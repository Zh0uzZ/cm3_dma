//------------------------------------------------------------------------------
// The confidential and proprietary information contained in this file may
// only be used by a person authorised under and to the extent permitted
// by a subsisting licensing agreement from ARM Limited.
//
//            (C) COPYRIGHT 2017 ARM Limited.
//                ALL RIGHTS RESERVED
//
// This entire notice must be reproduced on all copies of this file
// and copies of this file may only be made by a person if such person is
// permitted to do so under the terms of a subsisting license agreement
// from ARM Limited.
//
//      SVN Information
//
//      Checked In          : $$
//
//      Revision            : $$
//
//      Release Information : CM3DesignStart-r0p0-02rel0
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Cortex-M3 DesignStart processor logic level
//------------------------------------------------------------------------------

module cortexm3ds_logic
(ISOLATEn, RETAINn, nTRST, SWCLKTCK, SWDITMS, TDI,
PORESETn, SYSRESETn, RSTBYPASS, CGBYPASS, FCLK, HCLK, TRACECLKIN, STCLK,
STCALIB, AUXFAULT, BIGEND, INTISR, INTNMI, HREADYI, HRDATAI, HRESPI,
IFLUSH, HREADYD, HRDATAD, HRESPD, EXRESPD, SE, HREADYS, HRDATAS, HRESPS,
EXRESPS, EDBGRQ, DBGRESTART, RXEV, SLEEPHOLDREQn, WICENREQ,
FIXMASTERTYPE, TSVALUEB, MPUDISABLE, DBGEN, NIDEN, CDBGPWRUPACK,
DNOTITRANS, TDO, nTDOEN, SWDOEN, SWDO, SWV, JTAGNSW, TRACECLK, TRACEDATA
, HTRANSI, HSIZEI, HADDRI, HBURSTI, HPROTI, MEMATTRI, HTRANSD, HSIZED,
HADDRD, HBURSTD, HPROTD, MEMATTRD, HMASTERD, EXREQD, HWRITED, HWDATAD,
HTRANSS, HSIZES, HADDRS, HBURSTS, HPROTS, MEMATTRS, HMASTERS, EXREQS,
HWRITES, HWDATAS, HMASTLOCKS, BRCHSTAT, HALTED, LOCKUP, SLEEPING,
SLEEPDEEP, ETMINTNUM, ETMINTSTAT, SYSRESETREQ, TXEV, TRCENA, CURRPRI,
DBGRESTARTED, SLEEPHOLDACKn, GATEHCLK, HTMDHADDR, HTMDHTRANS, HTMDHSIZE,
HTMDHBURST, HTMDHPROT, HTMDHWDATA, HTMDHWRITE, HTMDHRDATA, HTMDHREADY,
HTMDHRESP, WICENACK, WAKEUP, CDBGPWRUPREQ, vis_r0_o, vis_r1_o, vis_r2_o,
vis_r3_o, vis_r4_o, vis_r5_o, vis_r6_o, vis_r7_o, vis_r8_o, vis_r9_o,
vis_r10_o, vis_r11_o, vis_r12_o, vis_msp_o, vis_psp_o, vis_pc_o);

input [25:0] STCALIB;
input [31:0] AUXFAULT;
input [239:0] INTISR;
input [31:0] HRDATAI;
input [1:0] HRESPI;
input [31:0] HRDATAD;
input [1:0] HRESPD;
input [31:0] HRDATAS;
input [1:0] HRESPS;
input [47:0] TSVALUEB;
output [3:0] TRACEDATA;
output [1:0] HTRANSI;
output [2:0] HSIZEI;
output [31:0] HADDRI;
output [2:0] HBURSTI;
output [3:0] HPROTI;
output [1:0] MEMATTRI;
output [1:0] HTRANSD;
output [2:0] HSIZED;
output [31:0] HADDRD;
output [2:0] HBURSTD;
output [3:0] HPROTD;
output [1:0] MEMATTRD;
output [1:0] HMASTERD;
output [31:0] HWDATAD;
output [1:0] HTRANSS;
output [2:0] HSIZES;
output [31:0] HADDRS;
output [2:0] HBURSTS;
output [3:0] HPROTS;
output [1:0] MEMATTRS;
output [1:0] HMASTERS;
output [31:0] HWDATAS;
output [3:0] BRCHSTAT;
output [8:0] ETMINTNUM;
output [2:0] ETMINTSTAT;
output [7:0] CURRPRI;
output [31:0] HTMDHADDR;
output [1:0] HTMDHTRANS;
output [2:0] HTMDHSIZE;
output [2:0] HTMDHBURST;
output [3:0] HTMDHPROT;
output [31:0] HTMDHWDATA;
output [31:0] HTMDHRDATA;
output [1:0] HTMDHRESP;
output [31:0] vis_r0_o;
output [31:0] vis_r1_o;
output [31:0] vis_r2_o;
output [31:0] vis_r3_o;
output [31:0] vis_r4_o;
output [31:0] vis_r5_o;
output [31:0] vis_r6_o;
output [31:0] vis_r7_o;
output [31:0] vis_r8_o;
output [31:0] vis_r9_o;
output [31:0] vis_r10_o;
output [31:0] vis_r11_o;
output [31:0] vis_r12_o;
output [31:2] vis_msp_o;
output [31:2] vis_psp_o;
output [31:1] vis_pc_o;
input ISOLATEn;
input RETAINn;
input nTRST;
input SWCLKTCK;
input SWDITMS;
input TDI;
input PORESETn;
input SYSRESETn;
input RSTBYPASS;
input CGBYPASS;
input FCLK;
input HCLK;
input TRACECLKIN;
input STCLK;
input BIGEND;
input INTNMI;
input HREADYI;
input IFLUSH;
input HREADYD;
input EXRESPD;
input SE;
input HREADYS;
input EXRESPS;
input EDBGRQ;
input DBGRESTART;
input RXEV;
input SLEEPHOLDREQn;
input WICENREQ;
input FIXMASTERTYPE;
input MPUDISABLE;
input DBGEN;
input NIDEN;
input CDBGPWRUPACK;
input DNOTITRANS;
output TDO;
output nTDOEN;
output SWDOEN;
output SWDO;
output SWV;
output JTAGNSW;
output TRACECLK;
output EXREQD;
output HWRITED;
output EXREQS;
output HWRITES;
output HMASTLOCKS;
output HALTED;
output LOCKUP;
output SLEEPING;
output SLEEPDEEP;
output SYSRESETREQ;
output TXEV;
output TRCENA;
output DBGRESTARTED;
output SLEEPHOLDACKn;
output GATEHCLK;
output HTMDHWRITE;
output HTMDHREADY;
output WICENACK;
output WAKEUP;
output CDBGPWRUPREQ;

wire Ox9dt6, Cy9dt6, Py9dt6, Ez9dt6, Sz9dt6, G0adt6, T0adt6, D1adt6, R1adt6, K2adt6;
wire W2adt6, H3adt6, S3adt6, D4adt6, M4adt6, Y4adt6, L5adt6, X5adt6, K6adt6, O7adt6;
wire P8adt6, O9adt6, Oaadt6, Pbadt6, Lcadt6, Kdadt6, Ieadt6, Ffadt6, Yfadt6, Zgadt6;
wire Aiadt6, Fjadt6, Kkadt6, Iladt6, Nmadt6, Inadt6, Doadt6, Dpadt6, Aqadt6, Dradt6;
wire Esadt6, Dtadt6, Fuadt6, Evadt6, Cwadt6, Xwadt6, Txadt6, Ryadt6, Ozadt6, R0bdt6;
wire L1bdt6, K2bdt6, L3bdt6, K4bdt6, M5bdt6, M6bdt6, G7bdt6, H8bdt6, A9bdt6, Aabdt6;
wire Cbbdt6, Bcbdt6, Ldbdt6, Uebdt6, Kgbdt6, Zhbdt6, Jjbdt6, Tkbdt6, Cmbdt6, Knbdt6;
wire Uobdt6, Bqbdt6, Mrbdt6, Usbdt6, Cubdt6, Ovbdt6, Axbdt6, Lybdt6, Ozbdt6, X0cdt6;
wire J2cdt6, T3cdt6, I5cdt6, S6cdt6, B8cdt6, L9cdt6, Pacdt6, Fccdt6, Qdcdt6, Efcdt6;
wire Sgcdt6, Uicdt6, Nlcdt6, Aocdt6, Crcdt6, Ztcdt6, Ywcdt6, Wzcdt6, A3ddt6, V5ddt6;
wire T8ddt6, Nbddt6, Geddt6, Zgddt6, Vjddt6, Mmddt6, Loddt6, Pqddt6, Xsddt6, Tuddt6;
wire Qwddt6, Qyddt6, M0edt6, I2edt6, F4edt6, B6edt6, Z7edt6, W9edt6, Acedt6, Zdedt6;
wire Ofedt6, Dhedt6, Siedt6, Hkedt6, Wledt6, Lnedt6, Apedt6, Pqedt6, Esedt6, Ttedt6;
wire Ivedt6, Xwedt6, Myedt6, B0fdt6, Q1fdt6, F3fdt6, U4fdt6, J6fdt6, Y7fdt6, N9fdt6;
wire Cbfdt6, Rcfdt6, Gefdt6, Vffdt6, Khfdt6, Zifdt6, Okfdt6, Dmfdt6, Snfdt6, Hpfdt6;
wire Wqfdt6, Lsfdt6, Iufdt6, Lwfdt6, Oyfdt6, N0gdt6, L2gdt6, O4gdt6, D6gdt6, S7gdt6;
wire H9gdt6, Wagdt6, Lcgdt6, Aegdt6, Pfgdt6, Ehgdt6, Djgdt6, Elgdt6, Cngdt6, Xpgdt6;
wire Bsgdt6, Fugdt6, Jwgdt6, Nygdt6, R0hdt6, V2hdt6, Z4hdt6, D7hdt6, Q9hdt6, Ubhdt6;
wire Oehdt6, Sghdt6, Wihdt6, Alhdt6, Enhdt6, Iphdt6, Vrhdt6, Zthdt6, Dwhdt6, Hyhdt6;
wire L0idt6, P2idt6, T4idt6, X6idt6, B9idt6, Fbidt6, Jdidt6, Nfidt6, Rhidt6, Vjidt6;
wire Zlidt6, Doidt6, Hqidt6, Xsidt6, Bvidt6, Fxidt6, Jzidt6, N1jdt6, R3jdt6, V5jdt6;
wire Z7jdt6, Dajdt6, Gcjdt6, Jejdt6, Mgjdt6, Pijdt6, Skjdt6, Vmjdt6, Yojdt6, Brjdt6;
wire Etjdt6, Hvjdt6, Kxjdt6, Nzjdt6, Q1kdt6, T3kdt6, W5kdt6, Z7kdt6, Cakdt6, Fckdt6;
wire Iekdt6, Lgkdt6, Oikdt6, Rkkdt6, Umkdt6, Xokdt6, Arkdt6, Mtkdt6, Pvkdt6, Sxkdt6;
wire Vzkdt6, Y1ldt6, B4ldt6, E6ldt6, H8ldt6, Kaldt6, Ncldt6, Qeldt6, Tgldt6, Wildt6;
wire Zkldt6, Cnldt6, Fpldt6, Irldt6, Ltldt6, Ovldt6, Rxldt6, Uzldt6, X1mdt6, A4mdt6;
wire D6mdt6, G8mdt6, Jamdt6, Mcmdt6, Pemdt6, Sgmdt6, Vimdt6, Ykmdt6, Bnmdt6, Epmdt6;
wire Dsmdt6, Cvmdt6, Bymdt6, A1ndt6, Z3ndt6, Y6ndt6, X9ndt6, Wcndt6, Vfndt6, Uindt6;
wire Tlndt6, Sondt6, Rrndt6, Qundt6, Pxndt6, O0odt6, N3odt6, M6odt6, L9odt6, Kcodt6;
wire Jfodt6, Iiodt6, Hlodt6, Goodt6, Frodt6, Euodt6, Dxodt6, C0pdt6, A3pdt6, Y5pdt6;
wire W8pdt6, Ubpdt6, Sepdt6, Qhpdt6, Okpdt6, Mnpdt6, Kqpdt6, Itpdt6, Gwpdt6, Ezpdt6;
wire C2qdt6, A5qdt6, Y7qdt6, Waqdt6, Udqdt6, Sgqdt6, Qjqdt6, Omqdt6, Mpqdt6, Ksqdt6;
wire Ivqdt6, Gyqdt6, E1rdt6, C4rdt6, A7rdt6, Y9rdt6, Wcrdt6, Ufrdt6, Sirdt6, Qlrdt6;
wire Oordt6, Mrrdt6, Kurdt6, Ixrdt6, G0sdt6, E3sdt6, C6sdt6, A9sdt6, Ybsdt6, Wesdt6;
wire Uhsdt6, Sksdt6, Qnsdt6, Oqsdt6, Mtsdt6, Kwsdt6, Izsdt6, G2tdt6, E5tdt6, C8tdt6;
wire Abtdt6, Ydtdt6, Wgtdt6, Ujtdt6, Smtdt6, Qptdt6, Ostdt6, Mvtdt6, Kytdt6, I1udt6;
wire G4udt6, E7udt6, Caudt6, Adudt6, Yfudt6, Wiudt6, Uludt6, Soudt6, Qrudt6, Ouudt6;
wire Mxudt6, K0vdt6, I3vdt6, G6vdt6, E9vdt6, Ccvdt6, Afvdt6, Yhvdt6, Wkvdt6, Unvdt6;
wire Sqvdt6, Qtvdt6, Owvdt6, Mzvdt6, K2wdt6, I5wdt6, G8wdt6, Ebwdt6, Bewdt6, Ygwdt6;
wire Vjwdt6, Smwdt6, Ppwdt6, Mswdt6, Jvwdt6, Gywdt6, D1xdt6, A4xdt6, S7xdt6, Q9xdt6;
wire Wbxdt6, Zdxdt6, Wfxdt6, Whxdt6, Mkxdt6, Smxdt6, Yoxdt6, Erxdt6, Ktxdt6, Qvxdt6;
wire Wxxdt6, C0ydt6, I2ydt6, O4ydt6, U6ydt6, A9ydt6, Gbydt6, Mdydt6, Sfydt6, Yhydt6;
wire Ekydt6, Kmydt6, Qoydt6, Wqydt6, Btydt6, Gvydt6, Lxydt6, Qzydt6, V1zdt6, A4zdt6;
wire F6zdt6, K8zdt6, Pazdt6, Uczdt6, Zezdt6, Ehzdt6, Jjzdt6, Olzdt6, Tnzdt6, Ypzdt6;
wire Dszdt6, Iuzdt6, Nwzdt6, Syzdt6, X00et6, C30et6, H50et6, M70et6, R90et6, Wb0et6;
wire Be0et6, Gg0et6, Li0et6, Qk0et6, Vm0et6, Ap0et6, Fr0et6, Kt0et6, Pv0et6, Ux0et6;
wire Zz0et6, E21et6, J41et6, O61et6, T81et6, Ya1et6, Dd1et6, If1et6, Nh1et6, Sj1et6;
wire Xl1et6, Co1et6, Hq1et6, Ms1et6, Ru1et6, Ww1et6, Bz1et6, G12et6, L32et6, Q52et6;
wire Z72et6, Ea2et6, Jc2et6, Oe2et6, Bh2et6, Nj2et6, Yl2et6, Po2et6, Gr2et6, Vt2et6;
wire Ow2et6, Ez2et6, W13et6, M43et6, K73et6, Ca3et6, Lc3et6, Ue3et6, Dh3et6, Mj3et6;
wire Vl3et6, Eo3et6, Nq3et6, Ws3et6, Fv3et6, Ox3et6, Xz3et6, G24et6, P44et6, Y64et6;
wire H94et6, Qb4et6, Zd4et6, Ig4et6, Ri4et6, Al4et6, Jn4et6, Sp4et6, Bs4et6, Ku4et6;
wire Tw4et6, Cz4et6, L15et6, U35et6, D65et6, M85et6, Va5et6, Ed5et6, Nf5et6, Wh5et6;
wire Fk5et6, Om5et6, Xo5et6, Gr5et6, Pt5et6, Yv5et6, Hy5et6, Q06et6, Z26et6, I56et6;
wire R76et6, Aa6et6, Jc6et6, Se6et6, Bh6et6, Kj6et6, Tl6et6, Co6et6, Lq6et6, Us6et6;
wire Dv6et6, Mx6et6, Vz6et6, E27et6, N47et6, W67et6, F97et6, Ob7et6, Xd7et6, Gg7et6;
wire Vi7et6, Pl7et6, No7et6, Ir7et6, Ku7et6, Ex7et6, Xz7et6, U28et6, P58et6, L88et6;
wire Ua8et6, Dd8et6, Mf8et6, Vh8et6, Ek8et6, Nm8et6, Wo8et6, Fr8et6, Ot8et6, Xv8et6;
wire Gy8et6, P09et6, Y29et6, H59et6, Q79et6, Z99et6, Ic9et6, Re9et6, Ah9et6, Jj9et6;
wire Sl9et6, Bo9et6, Kq9et6, Ts9et6, Cv9et6, Lx9et6, Uz9et6, D2aet6, M4aet6, V6aet6;
wire E9aet6, Nbaet6, Wdaet6, Fgaet6, Oiaet6, Xkaet6, Gnaet6, Ppaet6, Yraet6, Huaet6;
wire Qwaet6, Zyaet6, I1bet6, R3bet6, A6bet6, J8bet6, Sabet6, Bdbet6, Kfbet6, Thbet6;
wire Pkbet6, Qmbet6, Qobet6, Oqbet6, Zrbet6, Itbet6, Qubet6, Awbet6, Lxbet6, Nybet6;
wire Vzbet6, E1cet6, L2cet6, U3cet6, D5cet6, O6cet6, A8cet6, E9cet6, Macet6, Wbcet6;
wire Hdcet6, Oecet6, Zfcet6, Fhcet6, Micet6, Sjcet6, Ykcet6, Emcet6, Sncet6, Gpcet6;
wire Uqcet6, Iscet6, Wtcet6, Kvcet6, Ywcet6, Mycet6, A0det6, O1det6, C3det6, Q4det6;
wire E6det6, S7det6, G9det6, Uadet6, Icdet6, Wddet6, Kfdet6, Ygdet6, Midet6, Akdet6;
wire Oldet6, Cndet6, Zodet6, Brdet6, Zsdet6, Zudet6, Ywdet6, Yydet6, X0eet6, W2eet6;
wire X4eet6, X6eet6, X8eet6, Cbeet6, Ddeet6, Ffeet6, Dheet6, Ijeet6, Mleet6, Nneet6;
wire Opeet6, Oreet6, Qteet6, Vveet6, Ayeet6, A0fet6, D2fet6, Y3fet6, T5fet6, R7fet6;
wire T9fet6, Hbfet6, Vcfet6, Jefet6, Xffet6, Lhfet6, Zifet6, Nkfet6, Bmfet6, Pnfet6;
wire Gpfet6, Lrfet6, Qtfet6, Ovfet6, Oxfet6, Ozfet6, S1get6, X3get6, V5get6, X7get6;
wire P9get6, Hcget6, Weget6, Phget6, Hkget6, Rmget6, Apget6, Orget6, Euget6, Qwget6;
wire Dzget6, P1het6, C4het6, P7het6, Cbhet6, Pehet6, Cihet6, Plhet6, Cphet6, Pshet6;
wire Cwhet6, Pzhet6, C3iet6, P6iet6, Caiet6, Pdiet6, Chiet6, Pkiet6, Coiet6, Priet6;
wire Cviet6, Pyiet6, C2jet6, P5jet6, C9jet6, Pcjet6, Cgjet6, Pjjet6, Cnjet6, Pqjet6;
wire Cujet6, Pxjet6, C1ket6, P4ket6, C8ket6, Pbket6, Cfket6, Piket6, Cmket6, Ppket6;
wire Ctket6, Pwket6, C0let6, P3let6, C7let6, Palet6, Celet6, Phlet6, Cllet6, Polet6;
wire Cslet6, Pvlet6, Czlet6, P2met6, C6met6, P9met6, Cdmet6, Pgmet6, Ckmet6, Pnmet6;
wire Crmet6, Pumet6, Cymet6, P1net6, C5net6, P8net6, Ccnet6, Senet6, Ihnet6, Ujnet6;
wire Gmnet6, Xnnet6, Spnet6, Ssnet6, Pvnet6, Iynet6, X0oet6, L3oet6, I6oet6, U8oet6;
wire Qboet6, Meoet6, Khoet6, Ekoet6, Wmoet6, Opoet6, Proet6, Qtoet6, Rvoet6, Sxoet6;
wire Tzoet6, U1pet6, V3pet6, W5pet6, X7pet6, Y9pet6, Zbpet6, Aepet6, Bgpet6, Cipet6;
wire Dkpet6, Empet6, Fopet6, Gqpet6, Hspet6, Iupet6, Jwpet6, Kypet6, L0qet6, M2qet6;
wire N4qet6, O6qet6, P8qet6, Qaqet6, Rcqet6, Seqet6, Tgqet6, Uiqet6, Vkqet6, Wmqet6;
wire Xoqet6, Yqqet6, Zsqet6, Avqet6, Bxqet6, Czqet6, D1ret6, E3ret6, F5ret6, G7ret6;
wire H9ret6, Ibret6, Jdret6, Kfret6, Lhret6, Mjret6, Nlret6, Onret6, Ppret6, Qrret6;
wire Rtret6, Svret6, Txret6, Uzret6, V1set6, W3set6, X5set6, Y7set6, Z9set6, Acset6;
wire Beset6, Cgset6, Diset6, Ekset6, Fmset6, Goset6, Hqset6, Isset6, Juset6, Kwset6;
wire Lyset6, M0tet6, N2tet6, O4tet6, P6tet6, Q8tet6, Ratet6, Sctet6, Tetet6, Ugtet6;
wire Vitet6, Wktet6, Xmtet6, Yotet6, Zqtet6, Attet6, Bvtet6, Cxtet6, Dztet6, E1uet6;
wire O3uet6, K6uet6, Y8uet6, Zauet6, Aduet6, Bfuet6, Chuet6, Djuet6, Eluet6, Fnuet6;
wire Gpuet6, Hruet6, Ituet6, Jvuet6, Kxuet6, Lzuet6, M1vet6, N3vet6, O5vet6, P7vet6;
wire Q9vet6, Rbvet6, Sdvet6, Tfvet6, Uhvet6, Vjvet6, Wlvet6, Xnvet6, Ypvet6, Zrvet6;
wire Auvet6, Bwvet6, Cyvet6, D0wet6, E2wet6, F4wet6, G6wet6, H8wet6, Iawet6, Jcwet6;
wire Kewet6, Lgwet6, Miwet6, Nkwet6, Omwet6, Powet6, Qqwet6, Rswet6, Suwet6, Twwet6;
wire Uywet6, V0xet6, W2xet6, X4xet6, Y6xet6, Z8xet6, Abxet6, Bdxet6, Cfxet6, Dhxet6;
wire Ejxet6, Flxet6, Gnxet6, Hpxet6, Irxet6, Jtxet6, Kvxet6, Qxxet6, Wzxet6, I2yet6;
wire S4yet6, M7yet6, X9yet6, Icyet6, Teyet6, Dhyet6, Sjyet6, Dmyet6, Woyet6, Hryet6;
wire Styet6, Ewyet6, Ryyet6, S0zet6, T2zet6, U4zet6, N7zet6, Gazet6, Xczet6, Mezet6;
wire Hgzet6, Bizet6, Rjzet6, Blzet6, Qmzet6, Cozet6, Ppzet6, Frzet6, Tszet6, Fvzet6;
wire Pxzet6, Pzzet6, P10ft6, P30ft6, P50ft6, P70ft6, P90ft6, Pb0ft6, Pd0ft6, Pf0ft6;
wire Ph0ft6, Pj0ft6, Pl0ft6, Zn0ft6, Lq0ft6, Bt0ft6, Ov0ft6, Ay0ft6, K01ft6, T21ft6;
wire F51ft6, U71ft6, Ja1ft6, Zb1ft6, Xc1ft6, Vd1ft6, Te1ft6, Rf1ft6, Pg1ft6, Nh1ft6;
wire Li1ft6, Jj1ft6, Tk1ft6, Dm1ft6, Nn1ft6, Xo1ft6, Hq1ft6, Rr1ft6, Ws1ft6, Cu1ft6;
wire Iv1ft6, Nw1ft6, Tx1ft6, Zy1ft6, D02ft6, M12ft6, W22ft6, L42ft6, Y52ft6, B82ft6;
wire Ea2ft6, Hc2ft6, Ke2ft6, Gg2ft6, Ei2ft6, Fk2ft6, Dm2ft6, Eo2ft6, Cq2ft6, Gs2ft6;
wire Hu2ft6, Gw2ft6, Gy2ft6, I03ft6, T13ft6, E33ft6, P43ft6, A63ft6, L73ft6, W83ft6;
wire Ha3ft6, Sb3ft6, Dd3ft6, Oe3ft6, Zf3ft6, Kh3ft6, Vi3ft6, Gk3ft6, Rl3ft6, Cn3ft6;
wire No3ft6, Yp3ft6, Jr3ft6, Us3ft6, Fu3ft6, Qv3ft6, Bx3ft6, My3ft6, Xz3ft6, I14ft6;
wire T24ft6, E44ft6, P54ft6, A74ft6, L84ft6, W94ft6, Qb4ft6, Id4ft6, Af4ft6, Ah4ft6;
wire Aj4ft6, Sk4ft6, Um4ft6, Po4ft6, Mq4ft6, Fs4ft6, Bu4ft6, Dw4ft6, Fy4ft6, A05ft6;
wire X15ft6, Q35ft6, M55ft6, O75ft6, J95ft6, Gb5ft6, Zc5ft6, Ve5ft6, Kg5ft6, Mi5ft6;
wire Hk5ft6, Em5ft6, Xn5ft6, Tp5ft6, Vr5ft6, Cu5ft6, Nw5ft6, Xy5ft6, D16ft6, Y26ft6;
wire E46ft6, H56ft6, X66ft6, D86ft6, I96ft6, La6ft6, Qb6ft6, Id6ft6, We6ft6, Og6ft6;
wire Ci6ft6, Ak6ft6, Tl6ft6, Ln6ft6, Ig27v6, Ci27v6, Rj27v6, Fl27v6, Mm27v6, Tn27v6;
wire Ap27v6, Hq27v6, Or27v6, Vs27v6, Nu27v6, Iw27v6, Px27v6, Wy27v6, D037v6, K137v6;
wire R237v6, Y337v6, F537v6, M637v6, T737v6, A937v6, Ha37v6, Ob37v6, Vc37v6, Ce37v6;
wire Jf37v6, Qg37v6, Xh37v6, Ej37v6, Lk37v6, Sl37v6, Zm37v6, Yo37v6, Gq37v6, Ur37v6;
wire Jt37v6, Bv37v6, Tw37v6, Ly37v6, D047v6, V147v6, I347v6, X447v6, P647v6, D847v6;
wire V947v6, Fb47v6, Oc47v6, Jd47v6, Ee47v6, Ye47v6, Qf47v6, Mg47v6, Kh47v6, Ii47v6;
wire Gj47v6, Ek47v6, Wk47v6, Sl47v6, Qm47v6, On47v6, Io47v6, Cp47v6, Up47v6, Mq47v6;
wire Qr47v6, Us47v6, Yt47v6, Jv47v6, Vw47v6, Fy47v6, Uz47v6, E157v6, M257v6, V357v6;
wire H557v6, S657v6, D857v6, R957v6, Ab57v6, Lc57v6, Ud57v6, Hf57v6, Tg57v6, Ii57v6;
wire Uj57v6, Cl57v6, Pm57v6, Yn57v6, Kp57v6, Tq57v6, Ds57v6, Lt57v6, Uu57v6, Hw57v6;
wire Sx57v6, Ez57v6, S067v6, F267v6, S367v6, D567v6, O667v6, X767v6, G967v6, Oa67v6;
wire Ub67v6, Uc67v6, Ud67v6, Ue67v6, Uf67v6, Ug67v6, Uh67v6, Ui67v6, Uj67v6, Uk67v6;
wire Ul67v6, Um67v6, Un67v6, Mp67v6, Gr67v6, At67v6, Zt67v6, Xu67v6, Vv67v6, Xw67v6;
wire Ox67v6, Fy67v6, Wy67v6, Xz67v6, T077v6, W177v6, A377v6, C477v6, X477v6, W577v6;
wire S677v6, O777v6, L877v6, I977v6, Sa77v6, Qc77v6, Ie77v6, Gg77v6, Uh77v6, Bj77v6;
wire Ok77v6, Gm77v6, Tn77v6, Dp77v6, Br77v6, Us77v6, Ru77v6, Uw77v6, Ty77v6, Q087v6;
wire G287v6, W387v6, L587v6, F787v6, B987v6, Ka87v6, Jc87v6, De87v6, Tf87v6, Ih87v6;
wire Fj87v6, Yk87v6, Xm87v6, Ro87v6, Uq87v6, Ds87v6, Mt87v6, Vu87v6, Ew87v6, Nx87v6;
wire Wy87v6, F097v6, O197v6, X297v6, G497v6, P597v6, Y697v6, H897v6, Q997v6, Za97v6;
wire Ic97v6, Rd97v6, Af97v6, Jg97v6, Sh97v6, Bj97v6, Kk97v6, Tl97v6, Cn97v6, Lo97v6;
wire Up97v6, Dr97v6, Ms97v6, Vt97v6, Ev97v6, Nw97v6, Cy97v6, Zz97v6, W1a7v6, W3a7v6;
wire Y5a7v6, U7a7v6, K9a7v6, Bba7v6, Vca7v6, Qea7v6, Oga7v6, Uia7v6, Rka7v6, Pma7v6;
wire Soa7v6, Mqa7v6, Gsa7v6, Lua7v6, Rwa7v6, Mya7v6, P0b7v6, J2b7v6, D4b7v6, T5b7v6;
wire P7b7v6, I9b7v6, Hbb7v6, Cdb7v6, Ifb7v6, Bhb7v6, Uib7v6, Tkb7v6, Rmb7v6, Oob7v6;
wire Hqb7v6, Jsb7v6, Ztb7v6, Qvb7v6, Qxb7v6, Lzb7v6, I1c7v6, Z2c7v6, Q4c7v6, N6c7v6;
wire H8c7v6, W9c7v6, Mbc7v6, Gdc7v6, Cfc7v6, Wgc7v6, Qic7v6, Kkc7v6, Emc7v6, Ync7v6;
wire Spc7v6, Frc7v6, Wsc7v6, Cuc7v6, Ivc7v6, Owc7v6, Uxc7v6, Azc7v6, G0d7v6, M1d7v6;
wire S2d7v6, Y3d7v6, E5d7v6, K6d7v6, Q7d7v6, W8d7v6, Cad7v6, Ibd7v6, Ocd7v6, Fed7v6;
wire Xfd7v6, Phd7v6, Fjd7v6, Kkd7v6, Bmd7v6, Lnd7v6, Vod7v6, Fqd7v6, Prd7v6, Zsd7v6;
wire Jud7v6, Tvd7v6, Dxd7v6, Nyd7v6, Xzd7v6, G1e7v6, M2e7v6, W3e7v6, B5e7v6, I6e7v6;
wire M7e7v6, M8e7v6, L9e7v6, Hae7v6, Hbe7v6, Hce7v6, Eee7v6, Lge7v6, Gie7v6, Jke7v6;
wire Ame7v6, Boe7v6, Zpe7v6, Xre7v6, Rte7v6, Kve7v6, Dxe7v6, Wye7v6, R0f7v6, F2f7v6;
wire A4f7v6, T5f7v6, J7f7v6, D9f7v6, Naf7v6, Xbf7v6, Hdf7v6, Ref7v6, Bgf7v6, Lhf7v6;
wire Vif7v6, Fkf7v6, Plf7v6, Zmf7v6, Jof7v6, Tpf7v6, Drf7v6, Ctf7v6, Vuf7v6, Mwf7v6;
wire Iyf7v6, P0g7v6, Z2g7v6, L5g7v6, X7g7v6, Jag7v6, Vcg7v6, Hfg7v6, Thg7v6, Vjg7v6;
wire Cmg7v6, Nog7v6, Brg7v6, Qtg7v6, Fwg7v6, Uyg7v6, J1h7v6, Y3h7v6, N6h7v6, W8h7v6;
wire D9h7v6, K9h7v6, R9h7v6, Y9h7v6, Fah7v6, Mah7v6, Tah7v6, Abh7v6, Hbh7v6, Obh7v6;
wire Vbh7v6, Cch7v6, Jch7v6, Qch7v6, Xch7v6, Edh7v6, Ldh7v6, Sdh7v6, Zdh7v6, Geh7v6;
wire Neh7v6, Ueh7v6, Bfh7v6, Ifh7v6, Pfh7v6, Wfh7v6, Dgh7v6, Kgh7v6, Rgh7v6, Ygh7v6;
wire Fhh7v6, Mhh7v6, Thh7v6, Aih7v6, Hih7v6, Oih7v6, Vih7v6, Cjh7v6, Jjh7v6, Qjh7v6;
wire Xjh7v6, Ekh7v6, Lkh7v6, Skh7v6, Zkh7v6, Glh7v6, Nlh7v6, Ulh7v6, Bmh7v6, Imh7v6;
wire Pmh7v6, Wmh7v6, Dnh7v6, Knh7v6, Rnh7v6, Ynh7v6, Foh7v6, Moh7v6, Toh7v6, Aph7v6;
wire Hph7v6, Oph7v6, Vph7v6, Cqh7v6, Jqh7v6, Qqh7v6, Xqh7v6, Erh7v6, Lrh7v6, Srh7v6;
wire Zrh7v6, Gsh7v6, Nsh7v6, Ush7v6, Bth7v6, Ith7v6, Pth7v6, Wth7v6, Duh7v6, Kuh7v6;
wire Ruh7v6, Yuh7v6, Fvh7v6, Mvh7v6, Tvh7v6, Awh7v6, Hwh7v6, Owh7v6, Vwh7v6, Cxh7v6;
wire Jxh7v6, Qxh7v6, Xxh7v6, Eyh7v6, Lyh7v6, Syh7v6, Zyh7v6, Gzh7v6, Nzh7v6, Uzh7v6;
wire B0i7v6, I0i7v6, P0i7v6, W0i7v6, D1i7v6, K1i7v6, R1i7v6, Y1i7v6, F2i7v6, M2i7v6;
wire T2i7v6, A3i7v6, H3i7v6, O3i7v6, V3i7v6, C4i7v6, J4i7v6, Q4i7v6, X4i7v6, E5i7v6;
wire L5i7v6, S5i7v6, Z5i7v6, G6i7v6, N6i7v6, U6i7v6, B7i7v6, I7i7v6, P7i7v6, W7i7v6;
wire D8i7v6, K8i7v6, R8i7v6, Y8i7v6, F9i7v6, M9i7v6, T9i7v6, Aai7v6, Hai7v6, Oai7v6;
wire Vai7v6, Cbi7v6, Jbi7v6, Qbi7v6, Xbi7v6, Eci7v6, Lci7v6, Sci7v6, Zci7v6, Gdi7v6;
wire Ndi7v6, Udi7v6, Bei7v6, Iei7v6, Pei7v6, Wei7v6, Dfi7v6, Kfi7v6, Rfi7v6, Yfi7v6;
wire Fgi7v6, Mgi7v6, Tgi7v6, Ahi7v6, Hhi7v6, Ohi7v6, Vhi7v6, Cii7v6, Jii7v6, Qii7v6;
wire Xii7v6, Eji7v6, Lji7v6, Sji7v6, Zji7v6, Gki7v6, Nki7v6, Uki7v6, Bli7v6, Ili7v6;
wire Pli7v6, Wli7v6, Dmi7v6, Kmi7v6, Rmi7v6, Ymi7v6, Fni7v6, Mni7v6, Tni7v6, Aoi7v6;
wire Hoi7v6, Ooi7v6, Voi7v6, Cpi7v6, Jpi7v6, Qpi7v6, Xpi7v6, Eqi7v6, Lqi7v6, Sqi7v6;
wire Zqi7v6, Gri7v6, Nri7v6, Uri7v6, Bsi7v6, Isi7v6, Psi7v6, Wsi7v6, Dti7v6, Kti7v6;
wire Rti7v6, Yti7v6, Fui7v6, Mui7v6, Tui7v6, Avi7v6, Hvi7v6, Ovi7v6, Vvi7v6, Cwi7v6;
wire Jwi7v6, Qwi7v6, Xwi7v6, Exi7v6, Lxi7v6, Sxi7v6, Zxi7v6, Gyi7v6, Nyi7v6, Uyi7v6;
wire Bzi7v6, Izi7v6, Pzi7v6, Wzi7v6, D0j7v6, K0j7v6, R0j7v6, Y0j7v6, F1j7v6, M1j7v6;
wire T1j7v6, A2j7v6, H2j7v6, O2j7v6, V2j7v6, C3j7v6, J3j7v6, Q3j7v6, X3j7v6, E4j7v6;
wire L4j7v6, S4j7v6, Z4j7v6, G5j7v6, N5j7v6, U5j7v6, B6j7v6, I6j7v6, P6j7v6, W6j7v6;
wire D7j7v6, K7j7v6, R7j7v6, Y7j7v6, F8j7v6, M8j7v6, T8j7v6, A9j7v6, H9j7v6, O9j7v6;
wire V9j7v6, Caj7v6, Jaj7v6, Qaj7v6, Xaj7v6, Ebj7v6, Lbj7v6, Sbj7v6, Zbj7v6, Gcj7v6;
wire Ncj7v6, Ucj7v6, Bdj7v6, Idj7v6, Pdj7v6, Wdj7v6, Dej7v6, Kej7v6, Rej7v6, Yej7v6;
wire Ffj7v6, Mfj7v6, Tfj7v6, Agj7v6, Hgj7v6, Ogj7v6, Vgj7v6, Chj7v6, Jhj7v6, Qhj7v6;
wire Xhj7v6, Eij7v6, Lij7v6, Sij7v6, Zij7v6, Gjj7v6, Njj7v6, Ujj7v6, Bkj7v6, Ikj7v6;
wire Pkj7v6, Wkj7v6, Dlj7v6, Klj7v6, Rlj7v6, Ylj7v6, Fmj7v6, Mmj7v6, Tmj7v6, Anj7v6;
wire Hnj7v6, Onj7v6, Vnj7v6, Coj7v6, Joj7v6, Qoj7v6, Xoj7v6, Epj7v6, Lpj7v6, Spj7v6;
wire Zpj7v6, Gqj7v6, Nqj7v6, Uqj7v6, Brj7v6, Irj7v6, Prj7v6, Wrj7v6, Dsj7v6, Ksj7v6;
wire Rsj7v6, Ysj7v6, Ftj7v6, Mtj7v6, Ttj7v6, Auj7v6, Huj7v6, Ouj7v6, Vuj7v6, Cvj7v6;
wire Jvj7v6, Qvj7v6, Xvj7v6, Ewj7v6, Lwj7v6, Swj7v6, Zwj7v6, Gxj7v6, Nxj7v6, Uxj7v6;
wire Byj7v6, Iyj7v6, Pyj7v6, Wyj7v6, Dzj7v6, Kzj7v6, Rzj7v6, Yzj7v6, F0k7v6, M0k7v6;
wire T0k7v6, A1k7v6, H1k7v6, O1k7v6, V1k7v6, C2k7v6, J2k7v6, Q2k7v6, X2k7v6, E3k7v6;
wire L3k7v6, S3k7v6, Z3k7v6, G4k7v6, N4k7v6, U4k7v6, B5k7v6, I5k7v6, P5k7v6, W5k7v6;
wire D6k7v6, K6k7v6, R6k7v6, Y6k7v6, F7k7v6, M7k7v6, T7k7v6, A8k7v6, H8k7v6, O8k7v6;
wire V8k7v6, C9k7v6, J9k7v6, Q9k7v6, X9k7v6, Eak7v6, Lak7v6, Sak7v6, Zak7v6, Gbk7v6;
wire Nbk7v6, Ubk7v6, Bck7v6, Ick7v6, Pck7v6, Wck7v6, Ddk7v6, Kdk7v6, Rdk7v6, Ydk7v6;
wire Fek7v6, Mek7v6, Tek7v6, Afk7v6, Hfk7v6, Ofk7v6, Vfk7v6, Cgk7v6, Jgk7v6, Qgk7v6;
wire Xgk7v6, Ehk7v6, Lhk7v6, Shk7v6, Zhk7v6, Gik7v6, Nik7v6, Uik7v6, Bjk7v6, Ijk7v6;
wire Pjk7v6, Wjk7v6, Dkk7v6, Kkk7v6, Rkk7v6, Ykk7v6, Flk7v6, Mlk7v6, Tlk7v6, Amk7v6;
wire Hmk7v6, Omk7v6, Vmk7v6, Cnk7v6, Jnk7v6, Qnk7v6, Xnk7v6, Eok7v6, Lok7v6, Sok7v6;
wire Zok7v6, Gpk7v6, Npk7v6, Upk7v6, Bqk7v6, Iqk7v6, Pqk7v6, Wqk7v6, Drk7v6, Krk7v6;
wire Rrk7v6, Yrk7v6, Fsk7v6, Msk7v6, Tsk7v6, Atk7v6, Htk7v6, Otk7v6, Vtk7v6, Cuk7v6;
wire Juk7v6, Quk7v6, Xuk7v6, Evk7v6, Lvk7v6, Svk7v6, Zvk7v6, Gwk7v6, Nwk7v6, Uwk7v6;
wire Bxk7v6, Ixk7v6, Pxk7v6, Wxk7v6, Dyk7v6, Kyk7v6, Ryk7v6, Yyk7v6, Fzk7v6, Mzk7v6;
wire Tzk7v6, A0l7v6, H0l7v6, O0l7v6, V0l7v6, C1l7v6, J1l7v6, Q1l7v6, X1l7v6, E2l7v6;
wire L2l7v6, S2l7v6, Z2l7v6, G3l7v6, N3l7v6, U3l7v6, B4l7v6, I4l7v6, P4l7v6, W4l7v6;
wire D5l7v6, K5l7v6, R5l7v6, Y5l7v6, F6l7v6, M6l7v6, T6l7v6, A7l7v6, H7l7v6, O7l7v6;
wire V7l7v6, C8l7v6, J8l7v6, Q8l7v6, X8l7v6, E9l7v6, L9l7v6, S9l7v6, Z9l7v6, Gal7v6;
wire Nal7v6, Ual7v6, Bbl7v6, Ibl7v6, Pbl7v6, Wbl7v6, Dcl7v6, Kcl7v6, Rcl7v6, Ycl7v6;
wire Fdl7v6, Mdl7v6, Tdl7v6, Ael7v6, Hel7v6, Oel7v6, Vel7v6, Cfl7v6, Jfl7v6, Qfl7v6;
wire Xfl7v6, Egl7v6, Lgl7v6, Sgl7v6, Zgl7v6, Ghl7v6, Nhl7v6, Uhl7v6, Bil7v6, Iil7v6;
wire Pil7v6, Wil7v6, Djl7v6, Kjl7v6, Rjl7v6, Yjl7v6, Fkl7v6, Mkl7v6, Tkl7v6, All7v6;
wire Hll7v6, Oll7v6, Vll7v6, Cml7v6, Jml7v6, Qml7v6, Xml7v6, Enl7v6, Lnl7v6, Snl7v6;
wire Znl7v6, Gol7v6, Nol7v6, Uol7v6, Bpl7v6, Ipl7v6, Ppl7v6, Wpl7v6, Dql7v6, Kql7v6;
wire Rql7v6, Yql7v6, Frl7v6, Mrl7v6, Trl7v6, Asl7v6, Hsl7v6, Osl7v6, Vsl7v6, Ctl7v6;
wire Jtl7v6, Qtl7v6, Xtl7v6, Eul7v6, Lul7v6, Sul7v6, Zul7v6, Gvl7v6, Nvl7v6, Uvl7v6;
wire Bwl7v6, Iwl7v6, Pwl7v6, Wwl7v6, Dxl7v6, Kxl7v6, Rxl7v6, Yxl7v6, Fyl7v6, Myl7v6;
wire Tyl7v6, Azl7v6, Hzl7v6, Ozl7v6, Vzl7v6, C0m7v6, J0m7v6, Q0m7v6, X0m7v6, E1m7v6;
wire L1m7v6, S1m7v6, Z1m7v6, G2m7v6, N2m7v6, U2m7v6, B3m7v6, I3m7v6, P3m7v6, W3m7v6;
wire D4m7v6, K4m7v6, R4m7v6, Y4m7v6, F5m7v6, M5m7v6, T5m7v6, A6m7v6, H6m7v6, O6m7v6;
wire V6m7v6, C7m7v6, J7m7v6, Q7m7v6, X7m7v6, E8m7v6, L8m7v6, S8m7v6, Z8m7v6, G9m7v6;
wire N9m7v6, U9m7v6, Bam7v6, Iam7v6, Pam7v6, Wam7v6, Dbm7v6, Kbm7v6, Rbm7v6, Ybm7v6;
wire Fcm7v6, Mcm7v6, Tcm7v6, Adm7v6, Hdm7v6, Odm7v6, Vdm7v6, Cem7v6, Jem7v6, Qem7v6;
wire Xem7v6, Efm7v6, Lfm7v6, Sfm7v6, Zfm7v6, Ggm7v6, Ngm7v6, Ugm7v6, Bhm7v6, Ihm7v6;
wire Phm7v6, Whm7v6, Dim7v6, Kim7v6, Rim7v6, Yim7v6, Fjm7v6, Mjm7v6, Tjm7v6, Akm7v6;
wire Hkm7v6, Okm7v6, Vkm7v6, Clm7v6, Jlm7v6, Qlm7v6, Xlm7v6, Emm7v6, Lmm7v6, Smm7v6;
wire Zmm7v6, Gnm7v6, Nnm7v6, Unm7v6, Bom7v6, Iom7v6, Pom7v6, Wom7v6, Dpm7v6, Kpm7v6;
wire Rpm7v6, Ypm7v6, Fqm7v6, Mqm7v6, Tqm7v6, Arm7v6, Hrm7v6, Orm7v6, Vrm7v6, Csm7v6;
wire Jsm7v6, Qsm7v6, Xsm7v6, Etm7v6, Ltm7v6, Stm7v6, Ztm7v6, Gum7v6, Num7v6, Uum7v6;
wire Bvm7v6, Ivm7v6, Pvm7v6, Wvm7v6, Dwm7v6, Kwm7v6, Rwm7v6, Ywm7v6, Fxm7v6, Mxm7v6;
wire Txm7v6, Aym7v6, Hym7v6, Oym7v6, Vym7v6, Czm7v6, Jzm7v6, Qzm7v6, Xzm7v6, E0n7v6;
wire L0n7v6, S0n7v6, Z0n7v6, G1n7v6, N1n7v6, U1n7v6, B2n7v6, I2n7v6, P2n7v6, W2n7v6;
wire D3n7v6, K3n7v6, R3n7v6, Y3n7v6, F4n7v6, M4n7v6, T4n7v6, A5n7v6, H5n7v6, O5n7v6;
wire V5n7v6, C6n7v6, J6n7v6, Q6n7v6, X6n7v6, E7n7v6, L7n7v6, S7n7v6, Z7n7v6, G8n7v6;
wire N8n7v6, U8n7v6, B9n7v6, I9n7v6, P9n7v6, W9n7v6, Dan7v6, Kan7v6, Ran7v6, Yan7v6;
wire Fbn7v6, Mbn7v6, Tbn7v6, Acn7v6, Hcn7v6, Ocn7v6, Vcn7v6, Cdn7v6, Jdn7v6, Qdn7v6;
wire Xdn7v6, Een7v6, Len7v6, Sen7v6, Zen7v6, Gfn7v6, Nfn7v6, Ufn7v6, Bgn7v6, Ign7v6;
wire Pgn7v6, Wgn7v6, Dhn7v6, Khn7v6, Rhn7v6, Yhn7v6, Fin7v6, Min7v6, Tin7v6, Ajn7v6;
wire Hjn7v6, Ojn7v6, Vjn7v6, Ckn7v6, Jkn7v6, Qkn7v6, Xkn7v6, Eln7v6, Lln7v6, Sln7v6;
wire Zln7v6, Gmn7v6, Nmn7v6, Umn7v6, Bnn7v6, Inn7v6, Pnn7v6, Wnn7v6, Don7v6, Kon7v6;
wire Ron7v6, Yon7v6, Fpn7v6, Mpn7v6, Tpn7v6, Aqn7v6, Hqn7v6, Oqn7v6, Vqn7v6, Crn7v6;
wire Jrn7v6, Qrn7v6, Xrn7v6, Esn7v6, Lsn7v6, Ssn7v6, Zsn7v6, Gtn7v6, Ntn7v6, Utn7v6;
wire Bun7v6, Iun7v6, Pun7v6, Wun7v6, Dvn7v6, Kvn7v6, Rvn7v6, Yvn7v6, Fwn7v6, Mwn7v6;
wire Twn7v6, Axn7v6, Hxn7v6, Oxn7v6, Vxn7v6, Cyn7v6, Jyn7v6, Qyn7v6, Xyn7v6, Ezn7v6;
wire Lzn7v6, Szn7v6, Zzn7v6, G0o7v6, N0o7v6, U0o7v6, B1o7v6, I1o7v6, P1o7v6, W1o7v6;
wire D2o7v6, K2o7v6, R2o7v6, Y2o7v6, F3o7v6, M3o7v6, T3o7v6, A4o7v6, H4o7v6, O4o7v6;
wire V4o7v6, C5o7v6, J5o7v6, Q5o7v6, X5o7v6, E6o7v6, L6o7v6, S6o7v6, Z6o7v6, G7o7v6;
wire N7o7v6, U7o7v6, B8o7v6, I8o7v6, P8o7v6, W8o7v6, D9o7v6, K9o7v6, R9o7v6, Y9o7v6;
wire Fao7v6, Mao7v6, Tao7v6, Abo7v6, Hbo7v6, Obo7v6, Vbo7v6, Cco7v6, Jco7v6, Qco7v6;
wire Xco7v6, Edo7v6, Ldo7v6, Sdo7v6, Zdo7v6, Geo7v6, Neo7v6, Ueo7v6, Bfo7v6, Ifo7v6;
wire Pfo7v6, Wfo7v6, Dgo7v6, Kgo7v6, Rgo7v6, Ygo7v6, Fho7v6, Mho7v6, Tho7v6, Aio7v6;
wire Hio7v6, Oio7v6, Vio7v6, Cjo7v6, Jjo7v6, Qjo7v6, Xjo7v6, Eko7v6, Lko7v6, Sko7v6;
wire Zko7v6, Glo7v6, Nlo7v6, Ulo7v6, Bmo7v6, Imo7v6, Pmo7v6, Wmo7v6, Dno7v6, Kno7v6;
wire Rno7v6, Yno7v6, Foo7v6, Moo7v6, Too7v6, Apo7v6, Hpo7v6, Opo7v6, Vpo7v6, Cqo7v6;
wire Jqo7v6, Qqo7v6, Xqo7v6, Ero7v6, Lro7v6, Sro7v6, Zro7v6, Gso7v6, Nso7v6, Uso7v6;
wire Bto7v6, Ito7v6, Pto7v6, Wto7v6, Duo7v6, Kuo7v6, Ruo7v6, Yuo7v6, Fvo7v6, Mvo7v6;
wire Tvo7v6, Awo7v6, Hwo7v6, Owo7v6, Vwo7v6, Cxo7v6, Jxo7v6, Qxo7v6, Xxo7v6, Eyo7v6;
wire Lyo7v6, Syo7v6, Zyo7v6, Gzo7v6, Nzo7v6, Uzo7v6, B0p7v6, I0p7v6, P0p7v6, W0p7v6;
wire D1p7v6, K1p7v6, R1p7v6, Y1p7v6, F2p7v6, M2p7v6, T2p7v6, A3p7v6, H3p7v6, O3p7v6;
wire V3p7v6, C4p7v6, J4p7v6, Q4p7v6, X4p7v6, E5p7v6, L5p7v6, S5p7v6, Z5p7v6, G6p7v6;
wire N6p7v6, U6p7v6, B7p7v6, I7p7v6, P7p7v6, W7p7v6, D8p7v6, K8p7v6, R8p7v6, Y8p7v6;
wire F9p7v6, M9p7v6, T9p7v6, Aap7v6, Hap7v6, Oap7v6, Vap7v6, Cbp7v6, Jbp7v6, Qbp7v6;
wire Xbp7v6, Ecp7v6, Lcp7v6, Scp7v6, Zcp7v6, Gdp7v6, Ndp7v6, Udp7v6, Bep7v6, Iep7v6;
wire Pep7v6, Wep7v6, Dfp7v6, Kfp7v6, Rfp7v6, Yfp7v6, Fgp7v6, Mgp7v6, Tgp7v6, Ahp7v6;
wire Hhp7v6, Ohp7v6, Vhp7v6, Cip7v6, Jip7v6, Qip7v6, Xip7v6, Ejp7v6, Ljp7v6, Sjp7v6;
wire Zjp7v6, Gkp7v6, Nkp7v6, Ukp7v6, Blp7v6, Ilp7v6, Plp7v6, Wlp7v6, Dmp7v6, Kmp7v6;
wire Rmp7v6, Ymp7v6, Fnp7v6, Mnp7v6, Tnp7v6, Aop7v6, Hop7v6, Oop7v6, Vop7v6, Cpp7v6;
wire Jpp7v6, Qpp7v6, Xpp7v6, Eqp7v6, Lqp7v6, Sqp7v6, Zqp7v6, Grp7v6, Nrp7v6, Urp7v6;
wire Bsp7v6, Isp7v6, Psp7v6, Wsp7v6, Dtp7v6, Ktp7v6, Rtp7v6, Ytp7v6, Fup7v6, Mup7v6;
wire Tup7v6, Avp7v6, Hvp7v6, Ovp7v6, Vvp7v6, Cwp7v6, Jwp7v6, Qwp7v6, Xwp7v6, Exp7v6;
wire Lxp7v6, Sxp7v6, Zxp7v6, Gyp7v6, Nyp7v6, Uyp7v6, Bzp7v6, Izp7v6, Pzp7v6, Wzp7v6;
wire D0q7v6, K0q7v6, R0q7v6, Y0q7v6, F1q7v6, M1q7v6, T1q7v6, A2q7v6, H2q7v6, O2q7v6;
wire V2q7v6, C3q7v6, J3q7v6, Q3q7v6, X3q7v6, E4q7v6, L4q7v6, S4q7v6, Z4q7v6, G5q7v6;
wire N5q7v6, U5q7v6, B6q7v6, I6q7v6, P6q7v6, W6q7v6, D7q7v6, K7q7v6, R7q7v6, Y7q7v6;
wire F8q7v6, M8q7v6, T8q7v6, A9q7v6, H9q7v6, O9q7v6, V9q7v6, Caq7v6, Jaq7v6, Qaq7v6;
wire Xaq7v6, Ebq7v6, Lbq7v6, Sbq7v6, Zbq7v6, Gcq7v6, Ncq7v6, Ucq7v6, Bdq7v6, Idq7v6;
wire Pdq7v6, Wdq7v6, Deq7v6, Keq7v6, Req7v6, Yeq7v6, Ffq7v6, Mfq7v6, Tfq7v6, Agq7v6;
wire Hgq7v6, Ogq7v6, Vgq7v6, Chq7v6, Jhq7v6, Qhq7v6, Xhq7v6, Eiq7v6, Liq7v6, Siq7v6;
wire Ziq7v6, Gjq7v6, Njq7v6, Ujq7v6, Bkq7v6, Ikq7v6, Pkq7v6, Wkq7v6, Dlq7v6, Klq7v6;
wire Rlq7v6, Ylq7v6, Fmq7v6, Mmq7v6, Tmq7v6, Anq7v6, Hnq7v6, Onq7v6, Vnq7v6, Coq7v6;
wire Joq7v6, Qoq7v6, Xoq7v6, Epq7v6, Lpq7v6, Spq7v6, Zpq7v6, Gqq7v6, Nqq7v6, Uqq7v6;
wire Brq7v6, Irq7v6, Prq7v6, Wrq7v6, Dsq7v6, Ksq7v6, Rsq7v6, Ysq7v6, Ftq7v6, Mtq7v6;
wire Ttq7v6, Auq7v6, Huq7v6, Ouq7v6, Vuq7v6, Cvq7v6, Jvq7v6, Qvq7v6, Xvq7v6, Ewq7v6;
wire Lwq7v6, Swq7v6, Zwq7v6, Gxq7v6, Nxq7v6, Uxq7v6, Byq7v6, Iyq7v6, Pyq7v6, Wyq7v6;
wire Dzq7v6, Kzq7v6, Rzq7v6, Yzq7v6, F0r7v6, M0r7v6, T0r7v6, A1r7v6, H1r7v6, O1r7v6;
wire V1r7v6, C2r7v6, J2r7v6, Q2r7v6, X2r7v6, E3r7v6, L3r7v6, S3r7v6, Z3r7v6, G4r7v6;
wire N4r7v6, U4r7v6, B5r7v6, I5r7v6, P5r7v6, W5r7v6, D6r7v6, K6r7v6, R6r7v6, Y6r7v6;
wire F7r7v6, M7r7v6, T7r7v6, A8r7v6, H8r7v6, O8r7v6, V8r7v6, C9r7v6, J9r7v6, Q9r7v6;
wire X9r7v6, Ear7v6, Lar7v6, Sar7v6, Zar7v6, Gbr7v6, Nbr7v6, Ubr7v6, Bcr7v6, Icr7v6;
wire Pcr7v6, Wcr7v6, Ddr7v6, Kdr7v6, Rdr7v6, Ydr7v6, Fer7v6, Mer7v6, Ter7v6, Afr7v6;
wire Hfr7v6, Ofr7v6, Vfr7v6, Cgr7v6, Jgr7v6, Qgr7v6, Xgr7v6, Ehr7v6, Lhr7v6, Shr7v6;
wire Zhr7v6, Gir7v6, Nir7v6, Uir7v6, Bjr7v6, Ijr7v6, Pjr7v6, Wjr7v6, Dkr7v6, Kkr7v6;
wire Rkr7v6, Ykr7v6, Flr7v6, Mlr7v6, Tlr7v6, Amr7v6, Hmr7v6, Omr7v6, Vmr7v6, Cnr7v6;
wire Jnr7v6, Qnr7v6, Xnr7v6, Eor7v6, Lor7v6, Sor7v6, Zor7v6, Gpr7v6, Npr7v6, Upr7v6;
wire Bqr7v6, Iqr7v6, Pqr7v6, Wqr7v6, Drr7v6, Krr7v6, Rrr7v6, Yrr7v6, Fsr7v6, Msr7v6;
wire Tsr7v6, Atr7v6, Htr7v6, Otr7v6, Vtr7v6, Cur7v6, Jur7v6, Qur7v6, Xur7v6, Evr7v6;
wire Lvr7v6, Svr7v6, Zvr7v6, Gwr7v6, Nwr7v6, Uwr7v6, Bxr7v6, Ixr7v6, Pxr7v6, Wxr7v6;
wire Dyr7v6, Kyr7v6, Ryr7v6, Yyr7v6, Fzr7v6, Mzr7v6, Tzr7v6, A0s7v6, H0s7v6, O0s7v6;
wire V0s7v6, C1s7v6, J1s7v6, Q1s7v6, X1s7v6, E2s7v6, L2s7v6, S2s7v6, Z2s7v6, G3s7v6;
wire N3s7v6, U3s7v6, B4s7v6, I4s7v6, P4s7v6, W4s7v6, D5s7v6, K5s7v6, R5s7v6, Y5s7v6;
wire F6s7v6, M6s7v6, T6s7v6, A7s7v6, H7s7v6, O7s7v6, V7s7v6, C8s7v6, J8s7v6, Q8s7v6;
wire X8s7v6, E9s7v6, L9s7v6, S9s7v6, Z9s7v6, Gas7v6, Nas7v6, Uas7v6, Bbs7v6, Ibs7v6;
wire Pbs7v6, Wbs7v6, Dcs7v6, Kcs7v6, Rcs7v6, Ycs7v6, Fds7v6, Mds7v6, Tds7v6, Aes7v6;
wire Hes7v6, Oes7v6, Ves7v6, Cfs7v6, Jfs7v6, Qfs7v6, Xfs7v6, Egs7v6, Lgs7v6, Sgs7v6;
wire Zgs7v6, Ghs7v6, Nhs7v6, Uhs7v6, Bis7v6, Iis7v6, Pis7v6, Wis7v6, Djs7v6, Kjs7v6;
wire Rjs7v6, Yjs7v6, Fks7v6, Mks7v6, Tks7v6, Als7v6, Hls7v6, Ols7v6, Vls7v6, Cms7v6;
wire Jms7v6, Qms7v6, Xms7v6, Ens7v6, Lns7v6, Sns7v6, Zns7v6, Gos7v6, Nos7v6, Uos7v6;
wire Bps7v6, Ips7v6, Pps7v6, Wps7v6, Dqs7v6, Kqs7v6, Rqs7v6, Yqs7v6, Frs7v6, Mrs7v6;
wire Trs7v6, Ass7v6, Hss7v6, Oss7v6, Vss7v6, Cts7v6, Jts7v6, Qts7v6, Xts7v6, Eus7v6;
wire Lus7v6, Sus7v6, Zus7v6, Gvs7v6, Nvs7v6, Uvs7v6, Bws7v6, Iws7v6, Pws7v6, Wws7v6;
wire Dxs7v6, Kxs7v6, Rxs7v6, Yxs7v6, Fys7v6, Mys7v6, Tys7v6, Azs7v6, Hzs7v6, Ozs7v6;
wire Vzs7v6, C0t7v6, J0t7v6, Q0t7v6, X0t7v6, E1t7v6, L1t7v6, S1t7v6, Z1t7v6, G2t7v6;
wire N2t7v6, U2t7v6, B3t7v6, I3t7v6, P3t7v6, W3t7v6, D4t7v6, K4t7v6, R4t7v6, Y4t7v6;
wire F5t7v6, M5t7v6, T5t7v6, A6t7v6, H6t7v6, O6t7v6, V6t7v6, C7t7v6, J7t7v6, Q7t7v6;
wire X7t7v6, E8t7v6, L8t7v6, S8t7v6, Z8t7v6, G9t7v6, N9t7v6, U9t7v6, Bat7v6, Iat7v6;
wire Pat7v6, Wat7v6, Dbt7v6, Kbt7v6, Rbt7v6, Ybt7v6, Fct7v6, Mct7v6, Tct7v6, Adt7v6;
wire Hdt7v6, Odt7v6, Vdt7v6, Cet7v6, Jet7v6, Qet7v6, Xet7v6, Eft7v6, Lft7v6, Sft7v6;
wire Zft7v6, Ggt7v6, Ngt7v6, Ugt7v6, Bht7v6, Iht7v6, Pht7v6, Wht7v6, Dit7v6, Kit7v6;
wire Rit7v6, Yit7v6, Fjt7v6, Mjt7v6, Tjt7v6, Akt7v6, Hkt7v6, Okt7v6, Vkt7v6, Clt7v6;
wire Jlt7v6, Qlt7v6, Xlt7v6, Emt7v6, Lmt7v6, Smt7v6, Zmt7v6, Gnt7v6, Nnt7v6, Unt7v6;
wire Bot7v6, Iot7v6, Pot7v6, Wot7v6, Dpt7v6, Kpt7v6, Rpt7v6, Ypt7v6, Fqt7v6, Mqt7v6;
wire Tqt7v6, Art7v6, Hrt7v6, Ort7v6, Vrt7v6, Cst7v6, Jst7v6, Qst7v6, Xst7v6, Ett7v6;
wire Ltt7v6, Stt7v6, Ztt7v6, Gut7v6, Nut7v6, Uut7v6, Bvt7v6, Ivt7v6, Pvt7v6, Wvt7v6;
wire Dwt7v6, Kwt7v6, Rwt7v6, Ywt7v6, Fxt7v6, Mxt7v6, Txt7v6, Ayt7v6, Hyt7v6, Oyt7v6;
wire Vyt7v6, Czt7v6, Jzt7v6, Qzt7v6, Xzt7v6, E0u7v6, L0u7v6, S0u7v6, Z0u7v6, G1u7v6;
wire N1u7v6, U1u7v6, B2u7v6, I2u7v6, P2u7v6, W2u7v6, D3u7v6, K3u7v6, R3u7v6, Y3u7v6;
wire F4u7v6, M4u7v6, T4u7v6, A5u7v6, H5u7v6, O5u7v6, V5u7v6, C6u7v6, J6u7v6, Q6u7v6;
wire X6u7v6, E7u7v6, L7u7v6, S7u7v6, Z7u7v6, G8u7v6, N8u7v6, U8u7v6, B9u7v6, I9u7v6;
wire P9u7v6, W9u7v6, Dau7v6, Kau7v6, Rau7v6, Yau7v6, Fbu7v6, Mbu7v6, Tbu7v6, Acu7v6;
wire Hcu7v6, Ocu7v6, Vcu7v6, Cdu7v6, Jdu7v6, Qdu7v6, Xdu7v6, Eeu7v6, Leu7v6, Seu7v6;
wire Zeu7v6, Gfu7v6, Nfu7v6, Ufu7v6, Bgu7v6, Igu7v6, Pgu7v6, Wgu7v6, Dhu7v6, Khu7v6;
wire Rhu7v6, Yhu7v6, Fiu7v6, Miu7v6, Tiu7v6, Aju7v6, Hju7v6, Oju7v6, Vju7v6, Cku7v6;
wire Jku7v6, Qku7v6, Xku7v6, Elu7v6, Llu7v6, Slu7v6, Zlu7v6, Gmu7v6, Nmu7v6, Umu7v6;
wire Bnu7v6, Inu7v6, Pnu7v6, Wnu7v6, Dou7v6, Kou7v6, Rou7v6, You7v6, Fpu7v6, Mpu7v6;
wire Tpu7v6, Aqu7v6, Hqu7v6, Oqu7v6, Vqu7v6, Cru7v6, Jru7v6, Qru7v6, Xru7v6, Esu7v6;
wire Lsu7v6, Ssu7v6, Zsu7v6, Gtu7v6, Ntu7v6, Utu7v6, Buu7v6, Iuu7v6, Puu7v6, Wuu7v6;
wire Dvu7v6, Kvu7v6, Rvu7v6, Yvu7v6, Fwu7v6, Mwu7v6, Twu7v6, Axu7v6, Hxu7v6, Oxu7v6;
wire Vxu7v6, Cyu7v6, Jyu7v6, Qyu7v6, Xyu7v6, Ezu7v6, Lzu7v6, Szu7v6, Zzu7v6, G0v7v6;
wire N0v7v6, U0v7v6, B1v7v6, I1v7v6, P1v7v6, W1v7v6, D2v7v6, K2v7v6, R2v7v6, Y2v7v6;
wire F3v7v6, M3v7v6, T3v7v6, A4v7v6, H4v7v6, O4v7v6, V4v7v6, C5v7v6, J5v7v6, Q5v7v6;
wire X5v7v6, E6v7v6, L6v7v6, S6v7v6, Z6v7v6, G7v7v6, N7v7v6, U7v7v6, B8v7v6, I8v7v6;
wire P8v7v6, W8v7v6, D9v7v6, K9v7v6, R9v7v6, Y9v7v6, Fav7v6, Mav7v6, Tav7v6, Abv7v6;
wire Hbv7v6, Obv7v6, Vbv7v6, Ccv7v6, Jcv7v6, Qcv7v6, Xcv7v6, Edv7v6, Ldv7v6, Sdv7v6;
wire Zdv7v6, Gev7v6, Nev7v6, Uev7v6, Bfv7v6, Ifv7v6, Pfv7v6, Wfv7v6, Dgv7v6, Kgv7v6;
wire Rgv7v6, Ygv7v6, Fhv7v6, Mhv7v6, Thv7v6, Aiv7v6, Hiv7v6, Oiv7v6, Viv7v6, Cjv7v6;
wire Jjv7v6, Qjv7v6, Xjv7v6, Ekv7v6, Lkv7v6, Skv7v6, Zkv7v6, Glv7v6, Nlv7v6, Ulv7v6;
wire Bmv7v6, Imv7v6, Pmv7v6, Wmv7v6, Dnv7v6, Knv7v6, Rnv7v6, Ynv7v6, Fov7v6, Mov7v6;
wire Tov7v6, Apv7v6, Hpv7v6, Opv7v6, Vpv7v6, Cqv7v6, Jqv7v6, Qqv7v6, Xqv7v6, Erv7v6;
wire Lrv7v6, Srv7v6, Zrv7v6, Gsv7v6, Nsv7v6, Usv7v6, Btv7v6, Itv7v6, Ptv7v6, Wtv7v6;
wire Duv7v6, Kuv7v6, Ruv7v6, Yuv7v6, Fvv7v6, Mvv7v6, Tvv7v6, Awv7v6, Hwv7v6, Owv7v6;
wire Vwv7v6, Cxv7v6, Jxv7v6, Qxv7v6, Xxv7v6, Eyv7v6, Lyv7v6, Syv7v6, Zyv7v6, Gzv7v6;
wire Nzv7v6, Uzv7v6, B0w7v6, I0w7v6, P0w7v6, W0w7v6, D1w7v6, K1w7v6, R1w7v6, Y1w7v6;
wire F2w7v6, M2w7v6, T2w7v6, A3w7v6, H3w7v6, O3w7v6, V3w7v6, C4w7v6, J4w7v6, Q4w7v6;
wire X4w7v6, E5w7v6, L5w7v6, S5w7v6, Z5w7v6, G6w7v6, N6w7v6, U6w7v6, B7w7v6, I7w7v6;
wire P7w7v6, W7w7v6, D8w7v6, K8w7v6, R8w7v6, Y8w7v6, F9w7v6, M9w7v6, T9w7v6, Aaw7v6;
wire Haw7v6, Oaw7v6, Vaw7v6, Cbw7v6, Jbw7v6, Qbw7v6, Xbw7v6, Ecw7v6, Lcw7v6, Scw7v6;
wire Zcw7v6, Gdw7v6, Ndw7v6, Udw7v6, Bew7v6, Iew7v6, Pew7v6, Wew7v6, Dfw7v6, Kfw7v6;
wire Rfw7v6, Yfw7v6, Fgw7v6, Mgw7v6, Tgw7v6, Ahw7v6, Hhw7v6, Ohw7v6, Vhw7v6, Ciw7v6;
wire Jiw7v6, Qiw7v6, Xiw7v6, Ejw7v6, Ljw7v6, Sjw7v6, Zjw7v6, Gkw7v6, Nkw7v6, Ukw7v6;
wire Blw7v6, Ilw7v6, Plw7v6, Wlw7v6, Dmw7v6, Kmw7v6, Rmw7v6, Ymw7v6, Fnw7v6, Mnw7v6;
wire Tnw7v6, Aow7v6, How7v6, Oow7v6, Vow7v6, Cpw7v6, Jpw7v6, Qpw7v6, Xpw7v6, Eqw7v6;
wire Lqw7v6, Sqw7v6, Zqw7v6, Grw7v6, Nrw7v6, Urw7v6, Bsw7v6, Isw7v6, Psw7v6, Wsw7v6;
wire Dtw7v6, Ktw7v6, Rtw7v6, Ytw7v6, Fuw7v6, Muw7v6, Tuw7v6, Avw7v6, Hvw7v6, Ovw7v6;
wire Vvw7v6, Cww7v6, Jww7v6, Qww7v6, Xww7v6, Exw7v6, Lxw7v6, Sxw7v6, Zxw7v6, Gyw7v6;
wire Nyw7v6, Uyw7v6, Bzw7v6, Izw7v6, Pzw7v6, Wzw7v6, D0x7v6, K0x7v6, R0x7v6, Y0x7v6;
wire F1x7v6, M1x7v6, T1x7v6, A2x7v6, H2x7v6, O2x7v6, V2x7v6, C3x7v6, J3x7v6, Q3x7v6;
wire X3x7v6, E4x7v6, L4x7v6, S4x7v6, Z4x7v6, G5x7v6, N5x7v6, U5x7v6, B6x7v6, I6x7v6;
wire P6x7v6, W6x7v6, D7x7v6, K7x7v6, R7x7v6, Y7x7v6, F8x7v6, M8x7v6, T8x7v6, A9x7v6;
wire H9x7v6, O9x7v6, V9x7v6, Cax7v6, Jax7v6, Qax7v6, Xax7v6, Ebx7v6, Lbx7v6, Sbx7v6;
wire Zbx7v6, Gcx7v6, Ncx7v6, Ucx7v6, Bdx7v6, Idx7v6, Pdx7v6, Wdx7v6, Dex7v6, Kex7v6;
wire Rex7v6, Yex7v6, Ffx7v6, Mfx7v6, Tfx7v6, Agx7v6, Hgx7v6, Ogx7v6, Vgx7v6, Chx7v6;
wire Jhx7v6, Qhx7v6, Xhx7v6, Eix7v6, Lix7v6, Six7v6, Zix7v6, Gjx7v6, Njx7v6, Ujx7v6;
wire Bkx7v6, Ikx7v6, Pkx7v6, Wkx7v6, Dlx7v6, Klx7v6, Rlx7v6, Ylx7v6, Fmx7v6, Mmx7v6;
wire Tmx7v6, Anx7v6, Hnx7v6, Onx7v6, Vnx7v6, Cox7v6, Jox7v6, Qox7v6, Xox7v6, Epx7v6;
wire Lpx7v6, Spx7v6, Zpx7v6, Gqx7v6, Nqx7v6, Uqx7v6, Brx7v6, Irx7v6, Prx7v6, Wrx7v6;
wire Dsx7v6, Ksx7v6, Rsx7v6, Ysx7v6, Ftx7v6, Mtx7v6, Ttx7v6, Aux7v6, Hux7v6, Oux7v6;
wire Vux7v6, Cvx7v6, Jvx7v6, Qvx7v6, Xvx7v6, Ewx7v6, Lwx7v6, Swx7v6, Zwx7v6, Gxx7v6;
wire Nxx7v6, Uxx7v6, Byx7v6, Iyx7v6, Pyx7v6, Wyx7v6, Dzx7v6, Kzx7v6, Rzx7v6, Yzx7v6;
wire F0y7v6, M0y7v6, T0y7v6, A1y7v6, H1y7v6, O1y7v6, V1y7v6, C2y7v6, J2y7v6, Q2y7v6;
wire X2y7v6, E3y7v6, L3y7v6, S3y7v6, Z3y7v6, G4y7v6, N4y7v6, U4y7v6, B5y7v6, I5y7v6;
wire P5y7v6, W5y7v6, D6y7v6, K6y7v6, R6y7v6, Y6y7v6, F7y7v6, M7y7v6, T7y7v6, A8y7v6;
wire H8y7v6, O8y7v6, V8y7v6, C9y7v6, J9y7v6, Q9y7v6, X9y7v6, Eay7v6, Lay7v6, Say7v6;
wire Zay7v6, Gby7v6, Nby7v6, Uby7v6, Bcy7v6, Icy7v6, Pcy7v6, Wcy7v6, Ddy7v6, Kdy7v6;
wire Rdy7v6, Ydy7v6, Fey7v6, Mey7v6, Tey7v6, Afy7v6, Hfy7v6, Ofy7v6, Vfy7v6, Cgy7v6;
wire Jgy7v6, Qgy7v6, Xgy7v6, Ehy7v6, Lhy7v6, Shy7v6, Zhy7v6, Giy7v6, Niy7v6, Uiy7v6;
wire Bjy7v6, Ijy7v6, Pjy7v6, Wjy7v6, Dky7v6, Kky7v6, Rky7v6, Yky7v6, Fly7v6, Mly7v6;
wire Tly7v6, Amy7v6, Hmy7v6, Omy7v6, Vmy7v6, Cny7v6, Jny7v6, Qny7v6, Xny7v6, Eoy7v6;
wire Loy7v6, Soy7v6, Zoy7v6, Gpy7v6, Npy7v6, Upy7v6, Bqy7v6, Iqy7v6, Pqy7v6, Wqy7v6;
wire Dry7v6, Kry7v6, Rry7v6, Yry7v6, Fsy7v6, Msy7v6, Tsy7v6, Aty7v6, Hty7v6, Oty7v6;
wire Vty7v6, Cuy7v6, Juy7v6, Quy7v6, Xuy7v6, Evy7v6, Lvy7v6, Svy7v6, Zvy7v6, Gwy7v6;
wire Nwy7v6, Uwy7v6, Bxy7v6, Ixy7v6, Pxy7v6, Wxy7v6, Dyy7v6, Kyy7v6, Ryy7v6, Yyy7v6;
wire Fzy7v6, Mzy7v6, Tzy7v6, A0z7v6, H0z7v6, O0z7v6, V0z7v6, C1z7v6, J1z7v6, Q1z7v6;
wire X1z7v6, E2z7v6, L2z7v6, S2z7v6, Z2z7v6, G3z7v6, N3z7v6, U3z7v6, B4z7v6, I4z7v6;
wire P4z7v6, W4z7v6, D5z7v6, K5z7v6, R5z7v6, Y5z7v6, F6z7v6, M6z7v6, T6z7v6, A7z7v6;
wire H7z7v6, O7z7v6, V7z7v6, C8z7v6, J8z7v6, Q8z7v6, X8z7v6, E9z7v6, L9z7v6, S9z7v6;
wire Z9z7v6, Gaz7v6, Naz7v6, Uaz7v6, Bbz7v6, Ibz7v6, Pbz7v6, Wbz7v6, Dcz7v6, Kcz7v6;
wire Rcz7v6, Ycz7v6, Fdz7v6, Mdz7v6, Tdz7v6, Aez7v6, Hez7v6, Oez7v6, Vez7v6, Cfz7v6;
wire Jfz7v6, Qfz7v6, Xfz7v6, Egz7v6, Lgz7v6, Sgz7v6, Zgz7v6, Ghz7v6, Nhz7v6, Uhz7v6;
wire Biz7v6, Iiz7v6, Piz7v6, Wiz7v6, Djz7v6, Kjz7v6, Rjz7v6, Yjz7v6, Fkz7v6, Mkz7v6;
wire Tkz7v6, Alz7v6, Hlz7v6, Olz7v6, Vlz7v6, Cmz7v6, Jmz7v6, Qmz7v6, Xmz7v6, Enz7v6;
wire Lnz7v6, Snz7v6, Znz7v6, Goz7v6, Noz7v6, Uoz7v6, Bpz7v6, Ipz7v6, Ppz7v6, Wpz7v6;
wire Dqz7v6, Kqz7v6, Rqz7v6, Yqz7v6, Frz7v6, Mrz7v6, Trz7v6, Asz7v6, Hsz7v6, Osz7v6;
wire Vsz7v6, Ctz7v6, Jtz7v6, Qtz7v6, Xtz7v6, Euz7v6, Luz7v6, Suz7v6, Zuz7v6, Gvz7v6;
wire Nvz7v6, Uvz7v6, Bwz7v6, Iwz7v6, Pwz7v6, Wwz7v6, Dxz7v6, Kxz7v6, Rxz7v6, Yxz7v6;
wire Fyz7v6, Myz7v6, Tyz7v6, Azz7v6, Hzz7v6, Ozz7v6, Vzz7v6, C008v6, J008v6, Q008v6;
wire X008v6, E108v6, L108v6, S108v6, Z108v6, G208v6, N208v6, U208v6, B308v6, I308v6;
wire P308v6, W308v6, D408v6, K408v6, R408v6, Y408v6, F508v6, M508v6, T508v6, A608v6;
wire H608v6, O608v6, V608v6, C708v6, J708v6, Q708v6, X708v6, E808v6, L808v6, S808v6;
wire Z808v6, G908v6, N908v6, U908v6, Ba08v6, Ia08v6, Pa08v6, Wa08v6, Db08v6, Kb08v6;
wire Rb08v6, Yb08v6, Fc08v6, Mc08v6, Tc08v6, Ad08v6, Hd08v6, Od08v6, Vd08v6, Ce08v6;
wire Je08v6, Qe08v6, Xe08v6, Ef08v6, Lf08v6, Sf08v6, Zf08v6, Gg08v6, Ng08v6, Ug08v6;
wire Bh08v6, Ih08v6, Ph08v6, Wh08v6, Di08v6, Ki08v6, Ri08v6, Yi08v6, Fj08v6, Mj08v6;
wire Tj08v6, Ak08v6, Hk08v6, Ok08v6, Vk08v6, Cl08v6, Jl08v6, Ql08v6, Xl08v6, Em08v6;
wire Lm08v6, Sm08v6, Zm08v6, Gn08v6, Nn08v6, Un08v6, Bo08v6, Io08v6, Po08v6, Wo08v6;
wire Dp08v6, Kp08v6, Rp08v6, Yp08v6, Fq08v6, Mq08v6, Tq08v6, Ar08v6, Hr08v6, Or08v6;
wire Vr08v6, Cs08v6, Js08v6, Qs08v6, Xs08v6, Et08v6, Lt08v6, St08v6, Zt08v6, Gu08v6;
wire Nu08v6, Uu08v6, Bv08v6, Iv08v6, Pv08v6, Wv08v6, Dw08v6, Kw08v6, Rw08v6, Yw08v6;
wire Fx08v6, Mx08v6, Tx08v6, Ay08v6, Hy08v6, Oy08v6, Vy08v6, Cz08v6, Jz08v6, Qz08v6;
wire Xz08v6, E018v6, L018v6, S018v6, Z018v6, G118v6, N118v6, U118v6, B218v6, I218v6;
wire P218v6, W218v6, D318v6, K318v6, R318v6, Y318v6, F418v6, M418v6, T418v6, A518v6;
wire H518v6, O518v6, V518v6, C618v6, J618v6, Q618v6, X618v6, E718v6, L718v6, S718v6;
wire Z718v6, G818v6, N818v6, U818v6, B918v6, I918v6, P918v6, W918v6, Da18v6, Ka18v6;
wire Ra18v6, Ya18v6, Fb18v6, Mb18v6, Tb18v6, Ac18v6, Hc18v6, Oc18v6, Vc18v6, Cd18v6;
wire Jd18v6, Qd18v6, Xd18v6, Ee18v6, Le18v6, Se18v6, Ze18v6, Gf18v6, Nf18v6, Uf18v6;
wire Bg18v6, Ig18v6, Pg18v6, Wg18v6, Dh18v6, Kh18v6, Rh18v6, Yh18v6, Fi18v6, Mi18v6;
wire Ti18v6, Aj18v6, Hj18v6, Oj18v6, Vj18v6, Ck18v6, Jk18v6, Qk18v6, Xk18v6, El18v6;
wire Ll18v6, Sl18v6, Zl18v6, Gm18v6, Nm18v6, Um18v6, Bn18v6, In18v6, Pn18v6, Wn18v6;
wire Do18v6, Ko18v6, Ro18v6, Yo18v6, Fp18v6, Mp18v6, Tp18v6, Aq18v6, Hq18v6, Oq18v6;
wire Vq18v6, Cr18v6, Jr18v6, Qr18v6, Xr18v6, Es18v6, Ls18v6, Ss18v6, Zs18v6, Gt18v6;
wire Nt18v6, Ut18v6, Bu18v6, Iu18v6, Pu18v6, Wu18v6, Dv18v6, Kv18v6, Rv18v6, Yv18v6;
wire Fw18v6, Mw18v6, Tw18v6, Ax18v6, Hx18v6, Ox18v6, Vx18v6, Cy18v6, Jy18v6, Qy18v6;
wire Xy18v6, Ez18v6, Lz18v6, Sz18v6, Zz18v6, G028v6, N028v6, U028v6, B128v6, I128v6;
wire P128v6, W128v6, D228v6, K228v6, R228v6, Y228v6, F328v6, M328v6, T328v6, A428v6;
wire H428v6, O428v6, V428v6, C528v6, J528v6, Q528v6, X528v6, E628v6, L628v6, S628v6;
wire Z628v6, G728v6, N728v6, U728v6, B828v6, I828v6, P828v6, W828v6, D928v6, K928v6;
wire R928v6, Y928v6, Fa28v6, Ma28v6, Ta28v6, Ab28v6, Hb28v6, Ob28v6, Vb28v6, Cc28v6;
wire Jc28v6, Qc28v6, Xc28v6, Ed28v6, Ld28v6, Sd28v6, Zd28v6, Ge28v6, Ne28v6, Ue28v6;
wire Bf28v6, If28v6, Pf28v6, Wf28v6, Dg28v6, Kg28v6, Rg28v6, Yg28v6, Fh28v6, Mh28v6;
wire Th28v6, Ai28v6, Hi28v6, Oi28v6, Vi28v6, Cj28v6, Jj28v6, Qj28v6, Xj28v6, Ek28v6;
wire Lk28v6, Sk28v6, Zk28v6, Gl28v6, Nl28v6, Ul28v6, Bm28v6, Im28v6, Pm28v6, Wm28v6;
wire Dn28v6, Kn28v6, Rn28v6, Yn28v6, Fo28v6, Mo28v6, To28v6, Ap28v6, Hp28v6, Op28v6;
wire Vp28v6, Cq28v6, Jq28v6, Qq28v6, Xq28v6, Er28v6, Lr28v6, Sr28v6, Zr28v6, Gs28v6;
wire Ns28v6, Us28v6, Bt28v6, It28v6, Pt28v6, Wt28v6, Du28v6, Ku28v6, Ru28v6, Yu28v6;
wire Fv28v6, Mv28v6, Tv28v6, Aw28v6, Hw28v6, Ow28v6, Vw28v6, Cx28v6, Jx28v6, Qx28v6;
wire Xx28v6, Ey28v6, Ly28v6, Sy28v6, Zy28v6, Gz28v6, Nz28v6, Uz28v6, B038v6, I038v6;
wire P038v6, W038v6, D138v6, K138v6, R138v6, Y138v6, F238v6, M238v6, T238v6, A338v6;
wire H338v6, O338v6, V338v6, C438v6, J438v6, Q438v6, X438v6, E538v6, L538v6, S538v6;
wire Z538v6, G638v6, N638v6, U638v6, B738v6, I738v6, P738v6, W738v6, D838v6, K838v6;
wire R838v6, Y838v6, F938v6, M938v6, T938v6, Aa38v6, Ha38v6, Oa38v6, Va38v6, Cb38v6;
wire Jb38v6, Qb38v6, Xb38v6, Ec38v6, Lc38v6, Sc38v6, Zc38v6, Gd38v6, Nd38v6, Ud38v6;
wire Be38v6, Ie38v6, Pe38v6, We38v6, Df38v6, Kf38v6, Rf38v6, Yf38v6, Fg38v6, Mg38v6;
wire Tg38v6, Ah38v6, Hh38v6, Oh38v6, Vh38v6, Ci38v6, Ji38v6, Qi38v6, Xi38v6, Ej38v6;
wire Lj38v6, Sj38v6, Zj38v6, Gk38v6, Nk38v6, Uk38v6, Bl38v6, Il38v6, Pl38v6, Wl38v6;
wire Dm38v6, Km38v6, Rm38v6, Ym38v6, Fn38v6, Mn38v6, Tn38v6, Ao38v6, Ho38v6, Oo38v6;
wire Vo38v6, Cp38v6, Jp38v6, Qp38v6, Xp38v6, Eq38v6, Lq38v6, Sq38v6, Zq38v6, Gr38v6;
wire Nr38v6, Ur38v6, Bs38v6, Is38v6, Ps38v6, Ws38v6, Dt38v6, Kt38v6, Rt38v6, Yt38v6;
wire Fu38v6, Mu38v6, Tu38v6, Av38v6, Hv38v6, Ov38v6, Vv38v6, Cw38v6, Jw38v6, Qw38v6;
wire Xw38v6, Ex38v6, Lx38v6, Sx38v6, Zx38v6, Gy38v6, Ny38v6, Uy38v6, Bz38v6, Iz38v6;
wire Pz38v6, Wz38v6, D048v6, K048v6, R048v6, Y048v6, F148v6, M148v6, T148v6, A248v6;
wire H248v6, O248v6, V248v6, C348v6, J348v6, Q348v6, X348v6, E448v6, L448v6, S448v6;
wire Z448v6, G548v6, N548v6, U548v6, B648v6, I648v6, P648v6, W648v6, D748v6, K748v6;
wire R748v6, Y748v6, F848v6, M848v6, T848v6, A948v6, H948v6, O948v6, V948v6, Ca48v6;
wire Ja48v6, Qa48v6, Xa48v6, Eb48v6, Lb48v6, Sb48v6, Zb48v6, Gc48v6, Nc48v6, Uc48v6;
wire Bd48v6, Id48v6, Pd48v6, Wd48v6, De48v6, Ke48v6, Re48v6, Ye48v6, Ff48v6, Mf48v6;
wire Tf48v6, Ag48v6, Hg48v6, Og48v6, Vg48v6, Ch48v6, Jh48v6, Qh48v6, Xh48v6, Ei48v6;
wire Li48v6, Si48v6, Zi48v6, Gj48v6, Nj48v6, Uj48v6, Bk48v6, Ik48v6, Pk48v6, Wk48v6;
wire Dl48v6, Kl48v6, Rl48v6, Yl48v6, Fm48v6, Mm48v6, Tm48v6, An48v6, Hn48v6, On48v6;
wire Vn48v6, Co48v6, Jo48v6, Qo48v6, Xo48v6, Ep48v6, Lp48v6, Sp48v6, Zp48v6, Gq48v6;
wire Nq48v6, Uq48v6, Br48v6, Ir48v6, Pr48v6, Wr48v6, Ds48v6, Ks48v6, Rs48v6, Ys48v6;
wire Ft48v6, Mt48v6, Tt48v6, Au48v6, Hu48v6, Ou48v6, Vu48v6, Cv48v6, Jv48v6, Qv48v6;
wire Xv48v6, Ew48v6, Lw48v6, Sw48v6, Zw48v6, Gx48v6, Nx48v6, Ux48v6, By48v6, Iy48v6;
wire Py48v6, Wy48v6, Dz48v6, Kz48v6, Rz48v6, Yz48v6, F058v6, M058v6, T058v6, A158v6;
wire H158v6, O158v6, V158v6, C258v6, J258v6, Q258v6, X258v6, E358v6, L358v6, S358v6;
wire Z358v6, G458v6, N458v6, U458v6, B558v6, I558v6, P558v6, W558v6, D658v6, K658v6;
wire R658v6, Y658v6, F758v6, M758v6, T758v6, A858v6, H858v6, O858v6, V858v6, C958v6;
wire J958v6, Q958v6, X958v6, Ea58v6, La58v6, Sa58v6, Za58v6, Gb58v6, Nb58v6, Ub58v6;
wire Bc58v6, Ic58v6, Pc58v6, Wc58v6, Dd58v6, Kd58v6, Rd58v6, Yd58v6, Fe58v6, Me58v6;
wire Te58v6, Af58v6, Hf58v6, Of58v6, Vf58v6, Cg58v6, Jg58v6, Qg58v6, Xg58v6, Eh58v6;
wire Lh58v6, Sh58v6, Zh58v6, Gi58v6, Ni58v6, Ui58v6, Bj58v6, Ij58v6, Pj58v6, Wj58v6;
wire Dk58v6, Kk58v6, Rk58v6, Yk58v6, Fl58v6, Ml58v6, Tl58v6, Am58v6, Hm58v6, Om58v6;
wire Vm58v6, Cn58v6, Jn58v6, Qn58v6, Xn58v6, Eo58v6, Lo58v6, So58v6, Zo58v6, Gp58v6;
wire Np58v6, Up58v6, Bq58v6, Iq58v6, Pq58v6, Wq58v6, Dr58v6, Kr58v6, Rr58v6, Yr58v6;
wire Fs58v6, Ms58v6, Ts58v6, At58v6, Ht58v6, Ot58v6, Vt58v6, Cu58v6, Ju58v6, Qu58v6;
wire Xu58v6, Ev58v6, Lv58v6, Sv58v6, Zv58v6, Gw58v6, Nw58v6, Uw58v6, Bx58v6, Ix58v6;
wire Px58v6, Wx58v6, Dy58v6, Ky58v6, Ry58v6, Yy58v6, Fz58v6, Mz58v6, Tz58v6, A068v6;
wire H068v6, O068v6, V068v6, C168v6, J168v6, Q168v6, X168v6, E268v6, L268v6, S268v6;
wire Z268v6, G368v6, N368v6, U368v6, B468v6, I468v6, P468v6, W468v6, D568v6, K568v6;
wire R568v6, Y568v6, F668v6, M668v6, T668v6, A768v6, H768v6, O768v6, V768v6, C868v6;
wire J868v6, Q868v6, X868v6, E968v6, L968v6, S968v6, Z968v6, Ga68v6, Na68v6, Ua68v6;
wire Bb68v6, Ib68v6, Pb68v6, Wb68v6, Dc68v6, Kc68v6, Rc68v6, Yc68v6, Fd68v6, Md68v6;
wire Td68v6, Ae68v6, He68v6, Oe68v6, Ve68v6, Cf68v6, Jf68v6, Qf68v6, Xf68v6, Eg68v6;
wire Lg68v6, Sg68v6, Zg68v6, Gh68v6, Nh68v6, Uh68v6, Bi68v6, Ii68v6, Pi68v6, Wi68v6;
wire Dj68v6, Kj68v6, Rj68v6, Yj68v6, Fk68v6, Mk68v6, Tk68v6, Al68v6, Hl68v6, Ol68v6;
wire Vl68v6, Cm68v6, Jm68v6, Qm68v6, Xm68v6, En68v6, Ln68v6, Sn68v6, Zn68v6, Go68v6;
wire No68v6, Uo68v6, Bp68v6, Ip68v6, Pp68v6, Wp68v6, Dq68v6, Kq68v6, Rq68v6, Yq68v6;
wire Fr68v6, Mr68v6, Tr68v6, As68v6, Hs68v6, Os68v6, Vs68v6, Ct68v6, Jt68v6, Qt68v6;
wire Xt68v6, Eu68v6, Lu68v6, Su68v6, Zu68v6, Gv68v6, Nv68v6, Uv68v6, Bw68v6, Iw68v6;
wire Pw68v6, Ww68v6, Dx68v6, Kx68v6, Rx68v6, Yx68v6, Fy68v6, My68v6, Ty68v6, Az68v6;
wire Hz68v6, Oz68v6, Vz68v6, C078v6, J078v6, Q078v6, X078v6, E178v6, L178v6, S178v6;
wire Z178v6, G278v6, N278v6, U278v6, B378v6, I378v6, P378v6, W378v6, D478v6, K478v6;
wire R478v6, Y478v6, F578v6, M578v6, T578v6, A678v6, H678v6, O678v6, V678v6, C778v6;
wire J778v6, Q778v6, X778v6, E878v6, L878v6, S878v6, Z878v6, G978v6, N978v6, U978v6;
wire Ba78v6, Ia78v6, Pa78v6, Wa78v6, Db78v6, Kb78v6, Rb78v6, Yb78v6, Fc78v6, Mc78v6;
wire Tc78v6, Ad78v6, Hd78v6, Od78v6, Vd78v6, Ce78v6, Je78v6, Qe78v6, Xe78v6, Ef78v6;
wire Lf78v6, Sf78v6, Zf78v6, Gg78v6, Ng78v6, Ug78v6, Bh78v6, Ih78v6, Ph78v6, Wh78v6;
wire Di78v6, Ki78v6, Ri78v6, Yi78v6, Fj78v6, Mj78v6, Tj78v6, Ak78v6, Hk78v6, Ok78v6;
wire Vk78v6, Cl78v6, Jl78v6, Ql78v6, Xl78v6, Em78v6, Lm78v6, Sm78v6, Zm78v6, Gn78v6;
wire Nn78v6, Un78v6, Bo78v6, Io78v6, Po78v6, Wo78v6, Dp78v6, Kp78v6, Rp78v6, Yp78v6;
wire Fq78v6, Mq78v6, Tq78v6, Ar78v6, Hr78v6, Or78v6, Vr78v6, Cs78v6, Js78v6, Qs78v6;
wire Xs78v6, Et78v6, Lt78v6, St78v6, Zt78v6, Gu78v6, Nu78v6, Uu78v6, Bv78v6, Iv78v6;
wire Pv78v6, Wv78v6, Dw78v6, Kw78v6, Rw78v6, Yw78v6, Fx78v6, Mx78v6, Tx78v6, Ay78v6;
wire Hy78v6, Oy78v6, Vy78v6, Cz78v6, Jz78v6, Qz78v6, Xz78v6, E088v6, L088v6, S088v6;
wire Z088v6, G188v6, N188v6, U188v6, B288v6, I288v6, P288v6, W288v6, D388v6, K388v6;
wire R388v6, Y388v6, F488v6, M488v6, T488v6, A588v6, H588v6, O588v6, V588v6, C688v6;
wire J688v6, Q688v6, X688v6, E788v6, L788v6, S788v6, Z788v6, G888v6, N888v6, U888v6;
wire B988v6, I988v6, P988v6, W988v6, Da88v6, Ka88v6, Ra88v6, Ya88v6, Fb88v6, Mb88v6;
wire Tb88v6, Ac88v6, Hc88v6, Oc88v6, Vc88v6, Cd88v6, Jd88v6, Qd88v6, Xd88v6, Ee88v6;
wire Le88v6, Se88v6, Ze88v6, Gf88v6, Nf88v6, Uf88v6, Bg88v6, Ig88v6, Pg88v6, Wg88v6;
wire Dh88v6, Kh88v6, Rh88v6, Yh88v6, Fi88v6, Mi88v6, Ti88v6, Aj88v6, Hj88v6, Oj88v6;
wire Vj88v6, Ck88v6, Jk88v6, Qk88v6, Xk88v6, El88v6, Ll88v6, Sl88v6, Zl88v6, Gm88v6;
wire Nm88v6, Um88v6, Bn88v6, In88v6, Pn88v6, Wn88v6, Do88v6, Ko88v6, Ro88v6, Yo88v6;
wire Fp88v6, Mp88v6, Tp88v6, Aq88v6, Hq88v6, Oq88v6, Vq88v6, Cr88v6, Jr88v6, Qr88v6;
wire Xr88v6, Es88v6, Ls88v6, Ss88v6, Zs88v6, Gt88v6, Nt88v6, Ut88v6, Bu88v6, Iu88v6;
wire Pu88v6, Wu88v6, Dv88v6, Kv88v6, Rv88v6, Yv88v6, Fw88v6, Mw88v6, Tw88v6, Ax88v6;
wire Hx88v6, Ox88v6, Vx88v6, Cy88v6, Jy88v6, Qy88v6, Xy88v6, Ez88v6, Lz88v6, Sz88v6;
wire Zz88v6, G098v6, N098v6, U098v6, B198v6, I198v6, P198v6, W198v6, D298v6, K298v6;
wire R298v6, Y298v6, F398v6, M398v6, T398v6, A498v6, H498v6, O498v6, V498v6, C598v6;
wire J598v6, Q598v6, X598v6, E698v6, L698v6, S698v6, Z698v6, G798v6, N798v6, U798v6;
wire B898v6, I898v6, P898v6, W898v6, D998v6, K998v6, R998v6, Y998v6, Fa98v6, Ma98v6;
wire Ta98v6, Ab98v6, Hb98v6, Ob98v6, Vb98v6, Cc98v6, Jc98v6, Qc98v6, Xc98v6, Ed98v6;
wire Ld98v6, Sd98v6, Zd98v6, Ge98v6, Ne98v6, Ue98v6, Bf98v6, If98v6, Pf98v6, Wf98v6;
wire Dg98v6, Kg98v6, Rg98v6, Yg98v6, Fh98v6, Mh98v6, Th98v6, Ai98v6, Hi98v6, Oi98v6;
wire Vi98v6, Cj98v6, Jj98v6, Qj98v6, Xj98v6, Ek98v6, Lk98v6, Sk98v6, Zk98v6, Gl98v6;
wire Nl98v6, Ul98v6, Bm98v6, Im98v6, Pm98v6, Wm98v6, Dn98v6, Kn98v6, Rn98v6, Yn98v6;
wire Fo98v6, Mo98v6, To98v6, Ap98v6, Hp98v6, Op98v6, Vp98v6, Cq98v6, Jq98v6, Qq98v6;
wire Xq98v6, Er98v6, Lr98v6, Sr98v6, Zr98v6, Gs98v6, Ns98v6, Us98v6, Bt98v6, It98v6;
wire Pt98v6, Wt98v6, Du98v6, Ku98v6, Ru98v6, Yu98v6, Fv98v6, Mv98v6, Tv98v6, Aw98v6;
wire Hw98v6, Ow98v6, Vw98v6, Cx98v6, Jx98v6, Qx98v6, Xx98v6, Ey98v6, Ly98v6, Sy98v6;
wire Zy98v6, Gz98v6, Nz98v6, Uz98v6, B0a8v6, I0a8v6, P0a8v6, W0a8v6, D1a8v6, K1a8v6;
wire R1a8v6, Y1a8v6, F2a8v6, M2a8v6, T2a8v6, A3a8v6, H3a8v6, O3a8v6, V3a8v6, C4a8v6;
wire J4a8v6, Q4a8v6, X4a8v6, E5a8v6, L5a8v6, S5a8v6, Z5a8v6, G6a8v6, N6a8v6, U6a8v6;
wire B7a8v6, I7a8v6, P7a8v6, W7a8v6, D8a8v6, K8a8v6, R8a8v6, Y8a8v6, F9a8v6, M9a8v6;
wire T9a8v6, Aaa8v6, Haa8v6, Oaa8v6, Vaa8v6, Cba8v6, Jba8v6, Qba8v6, Xba8v6, Eca8v6;
wire Lca8v6, Sca8v6, Zca8v6, Gda8v6, Nda8v6, Uda8v6, Bea8v6, Iea8v6, Pea8v6, Wea8v6;
wire Dfa8v6, Kfa8v6, Rfa8v6, Yfa8v6, Fga8v6, Mga8v6, Tga8v6, Aha8v6, Hha8v6, Oha8v6;
wire Vha8v6, Cia8v6, Jia8v6, Qia8v6, Xia8v6, Eja8v6, Lja8v6, Sja8v6, Zja8v6, Gka8v6;
wire Nka8v6, Uka8v6, Bla8v6, Ila8v6, Pla8v6, Wla8v6, Dma8v6, Kma8v6, Rma8v6, Yma8v6;
wire Fna8v6, Mna8v6, Tna8v6, Aoa8v6, Hoa8v6, Ooa8v6, Voa8v6, Cpa8v6, Jpa8v6, Qpa8v6;
wire Xpa8v6, Eqa8v6, Lqa8v6, Sqa8v6, Zqa8v6, Gra8v6, Nra8v6, Ura8v6, Bsa8v6, Isa8v6;
wire Psa8v6, Wsa8v6, Dta8v6, Kta8v6, Rta8v6, Yta8v6, Fua8v6, Mua8v6, Tua8v6, Ava8v6;
wire Hva8v6, Ova8v6, Vva8v6, Cwa8v6, Jwa8v6, Qwa8v6, Xwa8v6, Exa8v6, Lxa8v6, Sxa8v6;
wire Zxa8v6, Gya8v6, Nya8v6, Uya8v6, Bza8v6, Iza8v6, Pza8v6, Wza8v6, D0b8v6, K0b8v6;
wire R0b8v6, Y0b8v6, F1b8v6, M1b8v6, T1b8v6, A2b8v6, H2b8v6, O2b8v6, V2b8v6, C3b8v6;
wire J3b8v6, Q3b8v6, X3b8v6, E4b8v6, L4b8v6, S4b8v6, Z4b8v6, G5b8v6, N5b8v6, U5b8v6;
wire B6b8v6, I6b8v6, P6b8v6, W6b8v6, D7b8v6, K7b8v6, R7b8v6, Y7b8v6, F8b8v6, M8b8v6;
wire T8b8v6, A9b8v6, H9b8v6, O9b8v6, V9b8v6, Cab8v6, Jab8v6, Qab8v6, Xab8v6, Ebb8v6;
wire Lbb8v6, Sbb8v6, Zbb8v6, Gcb8v6, Ncb8v6, Ucb8v6, Bdb8v6, Idb8v6, Pdb8v6, Wdb8v6;
wire Deb8v6, Keb8v6, Reb8v6, Yeb8v6, Ffb8v6, Mfb8v6, Tfb8v6, Agb8v6, Hgb8v6, Ogb8v6;
wire Vgb8v6, Chb8v6, Jhb8v6, Qhb8v6, Xhb8v6, Eib8v6, Lib8v6, Sib8v6, Zib8v6, Gjb8v6;
wire Njb8v6, Ujb8v6, Bkb8v6, Ikb8v6, Pkb8v6, Wkb8v6, Dlb8v6, Klb8v6, Rlb8v6, Ylb8v6;
wire Fmb8v6, Mmb8v6, Tmb8v6, Anb8v6, Hnb8v6, Onb8v6, Vnb8v6, Cob8v6, Job8v6, Qob8v6;
wire Xob8v6, Epb8v6, Lpb8v6, Spb8v6, Zpb8v6, Gqb8v6, Nqb8v6, Uqb8v6, Brb8v6, Irb8v6;
wire Prb8v6, Wrb8v6, Dsb8v6, Ksb8v6, Rsb8v6, Ysb8v6, Ftb8v6, Mtb8v6, Ttb8v6, Aub8v6;
wire Hub8v6, Oub8v6, Vub8v6, Cvb8v6, Jvb8v6, Qvb8v6, Xvb8v6, Ewb8v6, Lwb8v6, Swb8v6;
wire Zwb8v6, Gxb8v6, Nxb8v6, Uxb8v6, Byb8v6, Iyb8v6, Pyb8v6, Wyb8v6, Dzb8v6, Kzb8v6;
wire Rzb8v6, Yzb8v6, F0c8v6, M0c8v6, T0c8v6, A1c8v6, H1c8v6, O1c8v6, V1c8v6, C2c8v6;
wire J2c8v6, Q2c8v6, X2c8v6, E3c8v6, L3c8v6, S3c8v6, Z3c8v6, G4c8v6, N4c8v6, U4c8v6;
wire B5c8v6, I5c8v6, P5c8v6, W5c8v6, D6c8v6, K6c8v6, R6c8v6, Y6c8v6, F7c8v6, M7c8v6;
wire T7c8v6, A8c8v6, H8c8v6, O8c8v6, V8c8v6, C9c8v6, J9c8v6, Q9c8v6, X9c8v6, Eac8v6;
wire Lac8v6, Sac8v6, Zac8v6, Gbc8v6, Nbc8v6, Ubc8v6, Bcc8v6, Icc8v6, Pcc8v6, Wcc8v6;
wire Ddc8v6, Kdc8v6, Rdc8v6, Ydc8v6, Fec8v6, Mec8v6, Tec8v6, Afc8v6, Hfc8v6, Ofc8v6;
wire Vfc8v6, Cgc8v6, Jgc8v6, Qgc8v6, Xgc8v6, Ehc8v6, Lhc8v6, Shc8v6, Zhc8v6, Gic8v6;
wire Nic8v6, Uic8v6, Bjc8v6, Ijc8v6, Pjc8v6, Wjc8v6, Dkc8v6, Kkc8v6, Rkc8v6, Ykc8v6;
wire Flc8v6, Mlc8v6, Tlc8v6, Amc8v6, Hmc8v6, Omc8v6, Vmc8v6, Cnc8v6, Jnc8v6, Qnc8v6;
wire Xnc8v6, Eoc8v6, Loc8v6, Soc8v6, Zoc8v6, Gpc8v6, Npc8v6, Upc8v6, Bqc8v6, Iqc8v6;
wire Pqc8v6, Wqc8v6, Drc8v6, Krc8v6, Rrc8v6, Yrc8v6, Fsc8v6, Msc8v6, Tsc8v6, Atc8v6;
wire Htc8v6, Otc8v6, Vtc8v6, Cuc8v6, Juc8v6, Quc8v6, Xuc8v6, Evc8v6, Lvc8v6, Svc8v6;
wire Zvc8v6, Gwc8v6, Nwc8v6, Uwc8v6, Bxc8v6, Ixc8v6, Pxc8v6, Wxc8v6, Dyc8v6, Kyc8v6;
wire Ryc8v6, Yyc8v6, Fzc8v6, Mzc8v6, Tzc8v6, A0d8v6, H0d8v6, O0d8v6, V0d8v6, C1d8v6;
wire J1d8v6, Q1d8v6, X1d8v6, E2d8v6, L2d8v6, S2d8v6, Z2d8v6, G3d8v6, N3d8v6, U3d8v6;
wire B4d8v6, I4d8v6, P4d8v6, W4d8v6, D5d8v6, K5d8v6, R5d8v6, Y5d8v6, F6d8v6, M6d8v6;
wire T6d8v6, A7d8v6, H7d8v6, O7d8v6, V7d8v6, C8d8v6, J8d8v6, Q8d8v6, X8d8v6, E9d8v6;
wire L9d8v6, S9d8v6, Z9d8v6, Gad8v6, Nad8v6, Uad8v6, Bbd8v6, Ibd8v6, Pbd8v6, Wbd8v6;
wire Dcd8v6, Kcd8v6, Rcd8v6, Ycd8v6, Fdd8v6, Mdd8v6, Tdd8v6, Aed8v6, Hed8v6, Oed8v6;
wire Ved8v6, Cfd8v6, Jfd8v6, Qfd8v6, Xfd8v6, Egd8v6, Lgd8v6, Sgd8v6, Zgd8v6, Ghd8v6;
wire Nhd8v6, Uhd8v6, Bid8v6, Iid8v6, Pid8v6, Wid8v6, Djd8v6, Kjd8v6, Rjd8v6, Yjd8v6;
wire Fkd8v6, Mkd8v6, Tkd8v6, Ald8v6, Hld8v6, Old8v6, Vld8v6, Cmd8v6, Jmd8v6, Qmd8v6;
wire Xmd8v6, End8v6, Lnd8v6, Snd8v6, Znd8v6, God8v6, Nod8v6, Uod8v6, Bpd8v6, Ipd8v6;
wire Ppd8v6, Wpd8v6, Dqd8v6, Kqd8v6, Rqd8v6, Yqd8v6, Frd8v6, Mrd8v6, Trd8v6, Asd8v6;
wire Hsd8v6, Osd8v6, Vsd8v6, Ctd8v6, Jtd8v6, Qtd8v6, Xtd8v6, Eud8v6, Lud8v6, Sud8v6;
wire Zud8v6, Gvd8v6, Nvd8v6, Uvd8v6, Bwd8v6, Iwd8v6, Pwd8v6, Wwd8v6, Dxd8v6, Kxd8v6;
wire Rxd8v6, Yxd8v6, Fyd8v6, Myd8v6, Tyd8v6, Azd8v6, Hzd8v6, Ozd8v6, Vzd8v6, C0e8v6;
wire J0e8v6, Q0e8v6, X0e8v6, E1e8v6, L1e8v6, S1e8v6, Z1e8v6, G2e8v6, N2e8v6, U2e8v6;
wire B3e8v6, I3e8v6, P3e8v6, W3e8v6, D4e8v6, K4e8v6, R4e8v6, Y4e8v6, F5e8v6, M5e8v6;
wire T5e8v6, A6e8v6, H6e8v6, O6e8v6, V6e8v6, C7e8v6, J7e8v6, Q7e8v6, X7e8v6, E8e8v6;
wire L8e8v6, S8e8v6, Z8e8v6, G9e8v6, N9e8v6, U9e8v6, Bae8v6, Iae8v6, Pae8v6, Wae8v6;
wire Dbe8v6, Kbe8v6, Rbe8v6, Ybe8v6, Fce8v6, Mce8v6, Tce8v6, Ade8v6, Hde8v6, Ode8v6;
wire Vde8v6, Cee8v6, Jee8v6, Qee8v6, Xee8v6, Efe8v6, Lfe8v6, Sfe8v6, Zfe8v6, Gge8v6;
wire Nge8v6, Uge8v6, Bhe8v6, Ihe8v6, Phe8v6, Whe8v6, Die8v6, Kie8v6, Rie8v6, Yie8v6;
wire Fje8v6, Mje8v6, Tje8v6, Ake8v6, Hke8v6, Oke8v6, Vke8v6, Cle8v6, Jle8v6, Qle8v6;
wire Xle8v6, Eme8v6, Lme8v6, Sme8v6, Zme8v6, Gne8v6, Nne8v6, Une8v6, Boe8v6, Ioe8v6;
wire Poe8v6, Woe8v6, Dpe8v6, Kpe8v6, Rpe8v6, Ype8v6, Fqe8v6, Mqe8v6, Tqe8v6, Are8v6;
wire Hre8v6, Ore8v6, Vre8v6, Cse8v6, Jse8v6, Qse8v6, Xse8v6, Ete8v6, Lte8v6, Ste8v6;
wire Zte8v6, Gue8v6, Nue8v6, Uue8v6, Bve8v6, Ive8v6, Pve8v6, Wve8v6, Dwe8v6, Kwe8v6;
wire Rwe8v6, Ywe8v6, Fxe8v6, Mxe8v6, Txe8v6, Aye8v6, Hye8v6, Oye8v6, Vye8v6, Cze8v6;
wire Jze8v6, Qze8v6, Xze8v6, E0f8v6, L0f8v6, S0f8v6, Z0f8v6, G1f8v6, N1f8v6, U1f8v6;
wire B2f8v6, I2f8v6, P2f8v6, W2f8v6, D3f8v6, K3f8v6, R3f8v6, Y3f8v6, F4f8v6, M4f8v6;
wire T4f8v6, A5f8v6, H5f8v6, O5f8v6, V5f8v6, C6f8v6, J6f8v6, Q6f8v6, X6f8v6, E7f8v6;
wire L7f8v6, S7f8v6, Z7f8v6, G8f8v6, N8f8v6, U8f8v6, B9f8v6, I9f8v6, P9f8v6, W9f8v6;
wire Daf8v6, Kaf8v6, Raf8v6, Yaf8v6, Fbf8v6, Mbf8v6, Tbf8v6, Acf8v6, Hcf8v6, Ocf8v6;
wire Vcf8v6, Cdf8v6, Jdf8v6, Qdf8v6, Xdf8v6, Eef8v6, Lef8v6, Sef8v6, Zef8v6, Gff8v6;
wire Nff8v6, Uff8v6, Bgf8v6, Igf8v6, Pgf8v6, Wgf8v6, Dhf8v6, Khf8v6, Rhf8v6, Yhf8v6;
wire Fif8v6, Mif8v6, Tif8v6, Ajf8v6, Hjf8v6, Ojf8v6, Vjf8v6, Ckf8v6, Jkf8v6, Qkf8v6;
wire Xkf8v6, Elf8v6, Llf8v6, Slf8v6, Zlf8v6, Gmf8v6, Nmf8v6, Umf8v6, Bnf8v6, Inf8v6;
wire Pnf8v6, Wnf8v6, Dof8v6, Kof8v6, Rof8v6, Yof8v6, Fpf8v6, Mpf8v6, Tpf8v6, Aqf8v6;
wire Hqf8v6, Oqf8v6, Vqf8v6, Crf8v6, Jrf8v6, Qrf8v6, Xrf8v6, Esf8v6, Lsf8v6, Ssf8v6;
wire Zsf8v6, Gtf8v6, Ntf8v6, Utf8v6, Buf8v6, Iuf8v6, Puf8v6, Wuf8v6, Dvf8v6, Kvf8v6;
wire Rvf8v6, Yvf8v6, Fwf8v6, Mwf8v6, Twf8v6, Axf8v6, Hxf8v6, Oxf8v6, Vxf8v6, Cyf8v6;
wire Jyf8v6, Qyf8v6, Xyf8v6, Ezf8v6, Lzf8v6, Szf8v6, Zzf8v6, G0g8v6, N0g8v6, U0g8v6;
wire B1g8v6, I1g8v6, P1g8v6, W1g8v6, D2g8v6, K2g8v6, R2g8v6, Y2g8v6, F3g8v6, M3g8v6;
wire T3g8v6, A4g8v6, H4g8v6, O4g8v6, V4g8v6, C5g8v6, J5g8v6, Q5g8v6, X5g8v6, E6g8v6;
wire L6g8v6, S6g8v6, Z6g8v6, G7g8v6, N7g8v6, U7g8v6, B8g8v6, I8g8v6, P8g8v6, W8g8v6;
wire D9g8v6, K9g8v6, R9g8v6, Y9g8v6, Fag8v6, Mag8v6, Tag8v6, Abg8v6, Hbg8v6, Obg8v6;
wire Vbg8v6, Ccg8v6, Jcg8v6, Qcg8v6, Xcg8v6, Edg8v6, Ldg8v6, Sdg8v6, Zdg8v6, Geg8v6;
wire Neg8v6, Ueg8v6, Bfg8v6, Ifg8v6, Pfg8v6, Wfg8v6, Dgg8v6, Kgg8v6, Rgg8v6, Ygg8v6;
wire Fhg8v6, Mhg8v6, Thg8v6, Aig8v6, Hig8v6, Oig8v6, Vig8v6, Cjg8v6, Jjg8v6, Qjg8v6;
wire Xjg8v6, Ekg8v6, Lkg8v6, Skg8v6, Zkg8v6, Glg8v6, Nlg8v6, Ulg8v6, Bmg8v6, Img8v6;
wire Pmg8v6, Wmg8v6, Dng8v6, Kng8v6, Rng8v6, Yng8v6, Fog8v6, Mog8v6, Tog8v6, Apg8v6;
wire Hpg8v6, Opg8v6, Vpg8v6, Cqg8v6, Jqg8v6, Qqg8v6, Xqg8v6, Erg8v6, Lrg8v6, Srg8v6;
wire Zrg8v6, Gsg8v6, Nsg8v6, Usg8v6, Btg8v6, Itg8v6, Ptg8v6, Wtg8v6, Dug8v6, Kug8v6;
wire Rug8v6, Yug8v6, Fvg8v6, Mvg8v6, Tvg8v6, Awg8v6, Hwg8v6, Owg8v6, Vwg8v6, Cxg8v6;
wire Jxg8v6, Qxg8v6, Xxg8v6, Eyg8v6, Lyg8v6, Syg8v6, Zyg8v6, Gzg8v6, Nzg8v6, Uzg8v6;
wire B0h8v6, I0h8v6, P0h8v6, W0h8v6, D1h8v6, K1h8v6, R1h8v6, Y1h8v6, F2h8v6, M2h8v6;
wire T2h8v6, A3h8v6, H3h8v6, O3h8v6, V3h8v6, C4h8v6, J4h8v6, Q4h8v6, X4h8v6, E5h8v6;
wire L5h8v6, S5h8v6, Z5h8v6, G6h8v6, N6h8v6, U6h8v6, B7h8v6, I7h8v6, P7h8v6, W7h8v6;
wire D8h8v6, K8h8v6, R8h8v6, Y8h8v6, F9h8v6, M9h8v6, T9h8v6, Aah8v6, Hah8v6, Oah8v6;
wire Vah8v6, Cbh8v6, Jbh8v6, Qbh8v6, Xbh8v6, Ech8v6, Lch8v6, Sch8v6, Zch8v6, Gdh8v6;
wire Ndh8v6, Udh8v6, Beh8v6, Ieh8v6, Peh8v6, Weh8v6, Dfh8v6, Kfh8v6, Rfh8v6, Yfh8v6;
wire Fgh8v6, Mgh8v6, Tgh8v6, Ahh8v6, Hhh8v6, Ohh8v6, Vhh8v6, Cih8v6, Jih8v6, Qih8v6;
wire Xih8v6, Ejh8v6, Ljh8v6, Sjh8v6, Zjh8v6, Gkh8v6, Nkh8v6, Ukh8v6, Blh8v6, Ilh8v6;
wire Plh8v6, Wlh8v6, Dmh8v6, Kmh8v6, Rmh8v6, Ymh8v6, Fnh8v6, Mnh8v6, Tnh8v6, Aoh8v6;
wire Hoh8v6, Ooh8v6, Voh8v6, Cph8v6, Jph8v6, Qph8v6, Xph8v6, Eqh8v6, Lqh8v6, Sqh8v6;
wire Zqh8v6, Grh8v6, Nrh8v6, Urh8v6, Bsh8v6, Ish8v6, Psh8v6, Wsh8v6, Dth8v6, Kth8v6;
wire Rth8v6, Yth8v6, Fuh8v6, Muh8v6, Tuh8v6, Avh8v6, Hvh8v6, Ovh8v6, Vvh8v6, Cwh8v6;
wire Jwh8v6, Qwh8v6, Xwh8v6, Exh8v6, Lxh8v6, Sxh8v6, Zxh8v6, Gyh8v6, Nyh8v6, Uyh8v6;
wire Bzh8v6, Izh8v6, Pzh8v6, Wzh8v6, D0i8v6, K0i8v6, R0i8v6, Y0i8v6, F1i8v6, M1i8v6;
wire T1i8v6, A2i8v6, H2i8v6, O2i8v6, V2i8v6, C3i8v6, J3i8v6, Q3i8v6, X3i8v6, E4i8v6;
wire L4i8v6, S4i8v6, Z4i8v6, G5i8v6, N5i8v6, U5i8v6, B6i8v6, I6i8v6, P6i8v6, W6i8v6;
wire D7i8v6, K7i8v6, R7i8v6, Y7i8v6, F8i8v6, M8i8v6, T8i8v6, A9i8v6, H9i8v6, O9i8v6;
wire V9i8v6, Cai8v6, Jai8v6, Qai8v6, Xai8v6, Ebi8v6, Lbi8v6, Sbi8v6, Zbi8v6, Gci8v6;
wire Nci8v6, Uci8v6, Bdi8v6, Idi8v6, Pdi8v6, Wdi8v6, Dei8v6, Kei8v6, Rei8v6, Yei8v6;
wire Ffi8v6, Mfi8v6, Tfi8v6, Agi8v6, Hgi8v6, Ogi8v6, Vgi8v6, Chi8v6, Jhi8v6, Qhi8v6;
wire Xhi8v6, Eii8v6, Lii8v6, Sii8v6, Zii8v6, Gji8v6, Nji8v6, Uji8v6, Bki8v6, Iki8v6;
wire Pki8v6, Wki8v6, Dli8v6, Kli8v6, Rli8v6, Yli8v6, Fmi8v6, Mmi8v6, Tmi8v6, Ani8v6;
wire Hni8v6, Oni8v6, Vni8v6, Coi8v6, Joi8v6, Qoi8v6, Xoi8v6, Epi8v6, Lpi8v6, Spi8v6;
wire Zpi8v6, Gqi8v6, Nqi8v6, Uqi8v6, Bri8v6, Iri8v6, Pri8v6, Wri8v6, Dsi8v6, Ksi8v6;
wire Rsi8v6, Ysi8v6, Fti8v6, Mti8v6, Tti8v6, Aui8v6, Hui8v6, Oui8v6, Vui8v6, Cvi8v6;
wire Jvi8v6, Qvi8v6, Xvi8v6, Ewi8v6, Lwi8v6, Swi8v6, Zwi8v6, Gxi8v6, Nxi8v6, Uxi8v6;
wire Byi8v6, Iyi8v6, Pyi8v6, Wyi8v6, Dzi8v6, Kzi8v6, Rzi8v6, Yzi8v6, F0j8v6, M0j8v6;
wire T0j8v6, A1j8v6, H1j8v6, O1j8v6, V1j8v6, C2j8v6, J2j8v6, Q2j8v6, X2j8v6, E3j8v6;
wire L3j8v6, S3j8v6, Z3j8v6, G4j8v6, N4j8v6, U4j8v6, B5j8v6, I5j8v6, P5j8v6, W5j8v6;
wire D6j8v6, K6j8v6, R6j8v6, Y6j8v6, F7j8v6, M7j8v6, T7j8v6, A8j8v6, H8j8v6, O8j8v6;
wire V8j8v6, C9j8v6, J9j8v6, Q9j8v6, X9j8v6, Eaj8v6, Laj8v6, Saj8v6, Zaj8v6, Gbj8v6;
wire Nbj8v6, Ubj8v6, Bcj8v6, Icj8v6, Pcj8v6, Wcj8v6, Ddj8v6, Kdj8v6, Rdj8v6, Ydj8v6;
wire Fej8v6, Mej8v6, Tej8v6, Afj8v6, Hfj8v6, Ofj8v6, Vfj8v6, Cgj8v6, Jgj8v6, Qgj8v6;
wire Xgj8v6, Ehj8v6, Lhj8v6, Shj8v6, Zhj8v6, Gij8v6, Nij8v6, Uij8v6, Bjj8v6, Ijj8v6;
wire Pjj8v6, Wjj8v6, Dkj8v6, Kkj8v6, Rkj8v6, Ykj8v6, Flj8v6, Mlj8v6, Tlj8v6, Amj8v6;
wire Hmj8v6, Omj8v6, Vmj8v6, Cnj8v6, Jnj8v6, Qnj8v6, Xnj8v6, Eoj8v6, Loj8v6, Soj8v6;
wire Zoj8v6, Gpj8v6, Npj8v6, Upj8v6, Bqj8v6, Iqj8v6, Pqj8v6, Wqj8v6, Drj8v6, Krj8v6;
wire Rrj8v6, Yrj8v6, Fsj8v6, Msj8v6, Tsj8v6, Atj8v6, Htj8v6, Otj8v6, Vtj8v6, Cuj8v6;
wire Juj8v6, Quj8v6, Xuj8v6, Evj8v6, Lvj8v6, Svj8v6, Zvj8v6, Gwj8v6, Nwj8v6, Uwj8v6;
wire Bxj8v6, Ixj8v6, Pxj8v6, Wxj8v6, Dyj8v6, Kyj8v6, Ryj8v6, Yyj8v6, Fzj8v6, Mzj8v6;
wire Tzj8v6, A0k8v6, H0k8v6, O0k8v6, V0k8v6, C1k8v6, J1k8v6, Q1k8v6, X1k8v6, E2k8v6;
wire L2k8v6, S2k8v6, Z2k8v6, G3k8v6, N3k8v6, U3k8v6, B4k8v6, I4k8v6, P4k8v6, W4k8v6;
wire D5k8v6, K5k8v6, R5k8v6, Y5k8v6, F6k8v6, M6k8v6, T6k8v6, A7k8v6, H7k8v6, O7k8v6;
wire V7k8v6, C8k8v6, J8k8v6, Q8k8v6, X8k8v6, E9k8v6, L9k8v6, S9k8v6, Z9k8v6, Gak8v6;
wire Nak8v6, Uak8v6, Bbk8v6, Ibk8v6, Pbk8v6, Wbk8v6, Dck8v6, Kck8v6, Rck8v6, Yck8v6;
wire Fdk8v6, Mdk8v6, Tdk8v6, Aek8v6, Hek8v6, Oek8v6, Vek8v6, Cfk8v6, Jfk8v6, Qfk8v6;
wire Xfk8v6, Egk8v6, Lgk8v6, Sgk8v6, Zgk8v6, Ghk8v6, Nhk8v6, Uhk8v6, Bik8v6, Iik8v6;
wire Pik8v6, Wik8v6, Djk8v6, Kjk8v6, Rjk8v6, Yjk8v6, Fkk8v6, Mkk8v6, Tkk8v6, Alk8v6;
wire Hlk8v6, Olk8v6, Vlk8v6, Cmk8v6, Jmk8v6, Qmk8v6, Xmk8v6, Enk8v6, Lnk8v6, Snk8v6;
wire Znk8v6, Gok8v6, Nok8v6, Uok8v6, Bpk8v6, Ipk8v6, Ppk8v6, Wpk8v6, Dqk8v6, Kqk8v6;
wire Rqk8v6, Yqk8v6, Frk8v6, Mrk8v6, Trk8v6, Ask8v6, Hsk8v6, Osk8v6, Vsk8v6, Ctk8v6;
wire Jtk8v6, Qtk8v6, Xtk8v6, Euk8v6, Luk8v6, Suk8v6, Zuk8v6, Gvk8v6, Nvk8v6, Uvk8v6;
wire Bwk8v6, Iwk8v6, Pwk8v6, Wwk8v6, Dxk8v6, Kxk8v6, Rxk8v6, Yxk8v6, Fyk8v6, Myk8v6;
wire Tyk8v6, Azk8v6, Hzk8v6, Ozk8v6, Vzk8v6, C0l8v6, J0l8v6, Q0l8v6, X0l8v6, E1l8v6;
wire L1l8v6, S1l8v6, Z1l8v6, G2l8v6, N2l8v6, U2l8v6, B3l8v6, I3l8v6, P3l8v6, W3l8v6;
wire D4l8v6, K4l8v6, R4l8v6, Y4l8v6, F5l8v6, M5l8v6, T5l8v6, A6l8v6, H6l8v6, O6l8v6;
wire V6l8v6, C7l8v6, J7l8v6, Q7l8v6, X7l8v6, E8l8v6, L8l8v6, S8l8v6, Z8l8v6, G9l8v6;
wire N9l8v6, U9l8v6, Bal8v6, Ial8v6, Pal8v6, Wal8v6, Dbl8v6, Kbl8v6, Rbl8v6, Ybl8v6;
wire Fcl8v6, Mcl8v6, Tcl8v6, Adl8v6, Hdl8v6, Odl8v6, Vdl8v6, Cel8v6, Jel8v6, Qel8v6;
wire Xel8v6, Efl8v6, Lfl8v6, Sfl8v6, Zfl8v6, Ggl8v6, Ngl8v6, Ugl8v6, Bhl8v6, Ihl8v6;
wire Phl8v6, Whl8v6, Dil8v6, Kil8v6, Ril8v6, Yil8v6, Fjl8v6, Mjl8v6, Tjl8v6, Akl8v6;
wire Hkl8v6, Okl8v6, Vkl8v6, Cll8v6, Jll8v6, Qll8v6, Xll8v6, Eml8v6, Lml8v6, Sml8v6;
wire Zml8v6, Gnl8v6, Nnl8v6, Unl8v6, Bol8v6, Iol8v6, Pol8v6, Wol8v6, Dpl8v6, Kpl8v6;
wire Rpl8v6, Ypl8v6, Fql8v6, Mql8v6, Tql8v6, Arl8v6, Hrl8v6, Orl8v6, Vrl8v6, Csl8v6;
wire Jsl8v6, Qsl8v6, Xsl8v6, Etl8v6, Ltl8v6, Stl8v6, Ztl8v6, Gul8v6, Nul8v6, Uul8v6;
wire Bvl8v6, Ivl8v6, Pvl8v6, Wvl8v6, Dwl8v6, Kwl8v6, Rwl8v6, Zyl8v6, H1m8v6, P3m8v6;
wire X5m8v6, F8m8v6, Gbm8v6, Hem8v6, Ihm8v6, Jkm8v6, Knm8v6, Lqm8v6, Mtm8v6, Nwm8v6;
wire Pzm8v6, R2n8v6, T5n8v6, V8n8v6, Xbn8v6, Zen8v6, Bin8v6, Dln8v6, Fon8v6, Hrn8v6;
wire Jun8v6, Lxn8v6, N0o8v6, P3o8v6, R6o8v6, T9o8v6, Vco8v6, Xfo8v6, Zio8v6, Bmo8v6;
wire Dpo8v6, Fso8v6, Gvo8v6, Hyo8v6, I1p8v6, J4p8v6, K7p8v6, Lap8v6, Mdp8v6, Ngp8v6;
wire Ojp8v6, Pmp8v6, Rpp8v6, Tsp8v6, Vvp8v6, Xyp8v6, Z1q8v6, B5q8v6, D8q8v6, Fbq8v6;
wire Heq8v6, Jhq8v6, Lkq8v6, Nnq8v6, Pqq8v6, Rtq8v6, Twq8v6, Vzq8v6, X2r8v6, Z5r8v6;
wire B9r8v6, Dcr8v6, Ffr8v6, Hir8v6, Xkr8v6, Nnr8v6, Dqr8v6, Tsr8v6, Svr8v6, Ryr8v6;
wire Q1s8v6, P4s8v6, O7s8v6, Nas8v6, Mds8v6, Lgs8v6, Kjs8v6, Jms8v6, Ips8v6, Hss8v6;
wire Gvs8v6, Fys8v6, E1t8v6, D4t8v6, C7t8v6, Bat8v6, Tct8v6, Let8v6, Bgt8v6, Rht8v6;
wire Hjt8v6, Ojt8v6, Vjt8v6, Ckt8v6, Jkt8v6, Qkt8v6, Xkt8v6, Elt8v6, Llt8v6, Slt8v6;
wire Zlt8v6, Gmt8v6, Nmt8v6, Umt8v6, Bnt8v6, Int8v6, Pnt8v6, Wnt8v6, Dot8v6, Kot8v6;
wire Rot8v6, Yot8v6, Fpt8v6, Mpt8v6, Tpt8v6, Aqt8v6, Hqt8v6, Oqt8v6, Vqt8v6, Crt8v6;
wire Jrt8v6, Qrt8v6, Xrt8v6, Est8v6, Lst8v6, Sst8v6, Zst8v6, Gtt8v6, Ntt8v6, Utt8v6;
wire But8v6, Iut8v6, Put8v6, Wut8v6, Dvt8v6, Kvt8v6, Rvt8v6, Yvt8v6, Fwt8v6, Mwt8v6;
wire Twt8v6, Axt8v6, Hxt8v6, Oxt8v6, Vxt8v6, Cyt8v6, Jyt8v6, Qyt8v6, Xyt8v6, Ezt8v6;
wire Lzt8v6, Szt8v6, Zzt8v6, G0u8v6, N0u8v6, U0u8v6, B1u8v6, I1u8v6, P1u8v6, W1u8v6;
wire D2u8v6, K2u8v6, R2u8v6, Y2u8v6, F3u8v6, M3u8v6, T3u8v6, A4u8v6, H4u8v6, O4u8v6;
wire V4u8v6, C5u8v6, J5u8v6, Q5u8v6, X5u8v6, E6u8v6, L6u8v6, S6u8v6, Z6u8v6, G7u8v6;
wire N7u8v6, U7u8v6, B8u8v6, I8u8v6, P8u8v6, W8u8v6, D9u8v6, K9u8v6, R9u8v6, Y9u8v6;
wire Fau8v6, Mau8v6, Tau8v6, Abu8v6, Hbu8v6, Obu8v6, Vbu8v6, Ccu8v6, Jcu8v6, Qcu8v6;
wire Xcu8v6, Edu8v6, Ldu8v6, Sdu8v6, Zdu8v6, Geu8v6, Neu8v6, Ueu8v6, Bfu8v6, Ifu8v6;
wire Pfu8v6, Wfu8v6, Dgu8v6, Kgu8v6, Rgu8v6, Ygu8v6, Fhu8v6, Mhu8v6, Thu8v6, Aiu8v6;
wire Hiu8v6, Oiu8v6, Viu8v6, Cju8v6, Jju8v6, Qju8v6, Xju8v6, Eku8v6, Lku8v6, Sku8v6;
wire Zku8v6, Glu8v6, Nlu8v6, Ulu8v6, Bmu8v6, Imu8v6, Pmu8v6, Wmu8v6, Dnu8v6, Knu8v6;
wire Rnu8v6, Ynu8v6, Fou8v6, Mou8v6, Tou8v6, Apu8v6, Hpu8v6, Opu8v6, Vpu8v6, Cqu8v6;
wire Jqu8v6, Qqu8v6, Xqu8v6, Eru8v6, Lru8v6, Sru8v6, Zru8v6, Gsu8v6, Nsu8v6, Usu8v6;
wire Btu8v6, Itu8v6, Ptu8v6, Wtu8v6, Duu8v6, Kuu8v6, Ruu8v6, Yuu8v6, Fvu8v6, Mvu8v6;
wire Tvu8v6, Awu8v6, Hwu8v6, Owu8v6, Vwu8v6, Cxu8v6, Jxu8v6, Qxu8v6, Xxu8v6, Eyu8v6;
wire Lyu8v6, Syu8v6, Zyu8v6, Gzu8v6, Nzu8v6, Uzu8v6, B0v8v6, I0v8v6, P0v8v6, W0v8v6;
wire D1v8v6, K1v8v6, R1v8v6, Y1v8v6, F2v8v6, M2v8v6, T2v8v6, A3v8v6, H3v8v6, O3v8v6;
wire V3v8v6, C4v8v6, J4v8v6, Q4v8v6, X4v8v6, E5v8v6, L5v8v6, S5v8v6, Z5v8v6, G6v8v6;
wire N6v8v6, U6v8v6, B7v8v6, I7v8v6, P7v8v6, W7v8v6, D8v8v6, K8v8v6, R8v8v6, Y8v8v6;
wire F9v8v6, M9v8v6, T9v8v6, Aav8v6, Hav8v6, Oav8v6, Vav8v6, Cbv8v6, Jbv8v6, Qbv8v6;
wire Xbv8v6, Ecv8v6, Lcv8v6, Scv8v6, Zcv8v6, Gdv8v6, Ndv8v6, Udv8v6, Bev8v6, Iev8v6;
wire Pev8v6, Wev8v6, Dfv8v6, Kfv8v6, Rfv8v6, Yfv8v6, Fgv8v6, Mgv8v6, Tgv8v6, Ahv8v6;
wire Hhv8v6, Ohv8v6, Vhv8v6, Civ8v6, Jiv8v6, Qiv8v6, Xiv8v6, Ejv8v6, Ljv8v6, Sjv8v6;
wire Zjv8v6, Gkv8v6, Nkv8v6, Ukv8v6, Blv8v6, Ilv8v6, Plv8v6, Wlv8v6, Dmv8v6, Kmv8v6;
wire Rmv8v6, Ymv8v6, Fnv8v6, Mnv8v6, Tnv8v6, Aov8v6, Hov8v6, Oov8v6, Vov8v6, Cpv8v6;
wire Jpv8v6, Qpv8v6, Xpv8v6, Eqv8v6, Lqv8v6, Sqv8v6, Zqv8v6, Grv8v6, Nrv8v6, Urv8v6;
wire Bsv8v6, Isv8v6, Psv8v6, Wsv8v6, Dtv8v6, Ktv8v6, Rtv8v6, Ytv8v6, Fuv8v6, Muv8v6;
wire Tuv8v6, Avv8v6, Hvv8v6, Ovv8v6, Vvv8v6, Cwv8v6, Jwv8v6, Qwv8v6, Xwv8v6, Exv8v6;
wire Lxv8v6, Sxv8v6, Zxv8v6, Gyv8v6, Nyv8v6, Uyv8v6, Bzv8v6, Izv8v6, Pzv8v6, Wzv8v6;
wire D0w8v6, K0w8v6, R0w8v6, Y0w8v6, F1w8v6, M1w8v6, T1w8v6, A2w8v6, H2w8v6, O2w8v6;
wire V2w8v6, C3w8v6, J3w8v6, Q3w8v6, X3w8v6, E4w8v6, L4w8v6, S4w8v6, Z4w8v6, G5w8v6;
wire N5w8v6, U5w8v6, B6w8v6, I6w8v6, P6w8v6, W6w8v6, D7w8v6, K7w8v6, R7w8v6, Y7w8v6;
wire F8w8v6, M8w8v6, T8w8v6, A9w8v6, H9w8v6, O9w8v6, V9w8v6, Caw8v6, Jaw8v6, Qaw8v6;
wire Xaw8v6, Ebw8v6, Lbw8v6, Sbw8v6, Zbw8v6, Gcw8v6, Ncw8v6, Ucw8v6, Bdw8v6, Idw8v6;
wire Pdw8v6, Wdw8v6, Dew8v6, Kew8v6, Rew8v6, Yew8v6, Ffw8v6, Mfw8v6, Tfw8v6, Agw8v6;
wire Hgw8v6, Ogw8v6, Vgw8v6, Chw8v6, Jhw8v6, Qhw8v6, Xhw8v6, Eiw8v6, Liw8v6, Siw8v6;
wire Ziw8v6, Gjw8v6, Njw8v6, Ujw8v6, Bkw8v6, Ikw8v6, Pkw8v6, Wkw8v6, Dlw8v6, Klw8v6;
wire Rlw8v6, Ylw8v6, Fmw8v6, Mmw8v6, Tmw8v6, Anw8v6, Hnw8v6, Onw8v6, Vnw8v6, Cow8v6;
wire Jow8v6, Qow8v6, Xow8v6, Epw8v6, Lpw8v6, Spw8v6, Zpw8v6, Gqw8v6, Nqw8v6, Uqw8v6;
wire Brw8v6, Irw8v6, Prw8v6, Wrw8v6, Dsw8v6, Ksw8v6, Rsw8v6, Ysw8v6, Ftw8v6, Mtw8v6;
wire Ttw8v6, Auw8v6, Huw8v6, Ouw8v6, Vuw8v6, Cvw8v6, Jvw8v6, Qvw8v6, Xvw8v6, Eww8v6;
wire Lww8v6, Sww8v6, Zww8v6, Gxw8v6, Nxw8v6, Uxw8v6, Byw8v6, Iyw8v6, Pyw8v6, Wyw8v6;
wire Dzw8v6, Kzw8v6, Rzw8v6, Yzw8v6, F0x8v6, M0x8v6, T0x8v6, A1x8v6, H1x8v6, O1x8v6;
wire V1x8v6, C2x8v6, J2x8v6, Q2x8v6, X2x8v6, E3x8v6, L3x8v6, S3x8v6, Z3x8v6, G4x8v6;
wire N4x8v6, U4x8v6, B5x8v6, I5x8v6, P5x8v6, W5x8v6, D6x8v6, K6x8v6, R6x8v6, Y6x8v6;
wire F7x8v6, M7x8v6, T7x8v6, A8x8v6, H8x8v6, O8x8v6, V8x8v6, C9x8v6, J9x8v6, Q9x8v6;
wire X9x8v6, Eax8v6, Lax8v6, Sax8v6, Zax8v6, Gbx8v6, Nbx8v6, Ubx8v6, Bcx8v6, Icx8v6;
wire Pcx8v6, Wcx8v6, Ddx8v6, Kdx8v6, Rdx8v6, Ydx8v6, Fex8v6, Mex8v6, Tex8v6, Afx8v6;
wire Hfx8v6, Ofx8v6, Vfx8v6, Cgx8v6, Jgx8v6, Qgx8v6, Xgx8v6, Ehx8v6, Lhx8v6, Shx8v6;
wire Zhx8v6, Gix8v6, Nix8v6, Uix8v6, Bjx8v6, Ijx8v6, Pjx8v6, Wjx8v6, Dkx8v6, Kkx8v6;
wire Rkx8v6, Ykx8v6, Flx8v6, Mlx8v6, Tlx8v6, Amx8v6, Hmx8v6, Omx8v6, Vmx8v6, Cnx8v6;
wire Jnx8v6, Qnx8v6, Xnx8v6, Eox8v6, Lox8v6, Sox8v6, Zox8v6, Gpx8v6, Npx8v6, Upx8v6;
wire Bqx8v6, Iqx8v6, Pqx8v6, Wqx8v6, Drx8v6, Krx8v6, Rrx8v6, Yrx8v6, Fsx8v6, Msx8v6;
wire Tsx8v6, Atx8v6, Htx8v6, Otx8v6, Vtx8v6, Cux8v6, Jux8v6, Qux8v6, Xux8v6, Evx8v6;
wire Lvx8v6, Svx8v6, Zvx8v6, Gwx8v6, Nwx8v6, Uwx8v6, Bxx8v6, Ixx8v6, Pxx8v6, Wxx8v6;
wire Dyx8v6, Kyx8v6, Ryx8v6, Yyx8v6, Fzx8v6, Mzx8v6, Tzx8v6, A0y8v6, H0y8v6, O0y8v6;
wire V0y8v6, C1y8v6, J1y8v6, Q1y8v6, X1y8v6, E2y8v6, L2y8v6, S2y8v6, Z2y8v6, G3y8v6;
wire N3y8v6, U3y8v6, B4y8v6, I4y8v6, P4y8v6, W4y8v6, D5y8v6, K5y8v6, R5y8v6, Y5y8v6;
wire F6y8v6, M6y8v6, T6y8v6, A7y8v6, H7y8v6, O7y8v6, V7y8v6, C8y8v6, J8y8v6, Q8y8v6;
wire X8y8v6, E9y8v6, L9y8v6, S9y8v6, Z9y8v6, Gay8v6, Nay8v6, Uay8v6, Bby8v6, Iby8v6;
wire Pby8v6, Wby8v6, Dcy8v6, Kcy8v6, Rcy8v6, Ycy8v6, Fdy8v6, Mdy8v6, Tdy8v6, Aey8v6;
wire Hey8v6, Oey8v6, Vey8v6, Cfy8v6, Jfy8v6, Qfy8v6, Xfy8v6, Egy8v6, Lgy8v6, Sgy8v6;
wire Zgy8v6, Ghy8v6, Nhy8v6, Uhy8v6, Biy8v6, Iiy8v6, Piy8v6, Wiy8v6, Djy8v6, Kjy8v6;
wire Rjy8v6, Yjy8v6, Fky8v6, Mky8v6, Tky8v6, Aly8v6, Hly8v6, Oly8v6, Vly8v6, Cmy8v6;
wire Jmy8v6, Qmy8v6, Xmy8v6, Eny8v6, Lny8v6, Sny8v6, Zny8v6, Goy8v6, Noy8v6, Uoy8v6;
wire Bpy8v6, Ipy8v6, Ppy8v6, Wpy8v6, Dqy8v6, Kqy8v6, Rqy8v6, Yqy8v6, Fry8v6, Mry8v6;
wire Try8v6, Asy8v6, Hsy8v6, Osy8v6, Vsy8v6, Cty8v6, Jty8v6, Qty8v6, Xty8v6, Euy8v6;
wire Luy8v6, Suy8v6, Zuy8v6, Gvy8v6, Nvy8v6, Uvy8v6, Bwy8v6, Iwy8v6, Pwy8v6, Wwy8v6;
wire Dxy8v6, Kxy8v6, Rxy8v6, Yxy8v6, Fyy8v6, Myy8v6, Tyy8v6, Azy8v6, Hzy8v6, Ozy8v6;
wire Vzy8v6, C0z8v6, J0z8v6, Q0z8v6, X0z8v6, E1z8v6, L1z8v6, S1z8v6, Z1z8v6, G2z8v6;
wire N2z8v6, U2z8v6, B3z8v6, I3z8v6, P3z8v6, W3z8v6, D4z8v6, K4z8v6, R4z8v6, Y4z8v6;
wire F5z8v6, M5z8v6, T5z8v6, A6z8v6, H6z8v6, O6z8v6, V6z8v6, C7z8v6, J7z8v6, Q7z8v6;
wire X7z8v6, E8z8v6, L8z8v6, S8z8v6, Z8z8v6, G9z8v6, N9z8v6, U9z8v6, Baz8v6, Iaz8v6;
wire Paz8v6, Waz8v6, Dbz8v6, Kbz8v6, Rbz8v6, Ybz8v6, Fcz8v6, Mcz8v6, Tcz8v6, Adz8v6;
wire Hdz8v6, Odz8v6, Vdz8v6, Cez8v6, Jez8v6, Qez8v6, Xez8v6, Efz8v6, Lfz8v6, Sfz8v6;
wire Zfz8v6, Ggz8v6, Ngz8v6, Ugz8v6, Bhz8v6, Ihz8v6, Phz8v6, Whz8v6, Diz8v6, Kiz8v6;
wire Riz8v6, Yiz8v6, Fjz8v6, Mjz8v6, Tjz8v6, Akz8v6, Hkz8v6, Okz8v6, Vkz8v6, Clz8v6;
wire Jlz8v6, Qlz8v6, Xlz8v6, Emz8v6, Lmz8v6, Smz8v6, Zmz8v6, Gnz8v6, Nnz8v6, Unz8v6;
wire Boz8v6, Ioz8v6, Poz8v6, Woz8v6, Dpz8v6, Kpz8v6, Rpz8v6, Ypz8v6, Fqz8v6, Mqz8v6;
wire Tqz8v6, Arz8v6, Hrz8v6, Orz8v6, Vrz8v6, Csz8v6, Jsz8v6, Qsz8v6, Xsz8v6, Etz8v6;
wire Ltz8v6, Stz8v6, Ztz8v6, Guz8v6, Nuz8v6, Uuz8v6, Bvz8v6, Ivz8v6, Pvz8v6, Wvz8v6;
wire Dwz8v6, Kwz8v6, Rwz8v6, Ywz8v6, Fxz8v6, Mxz8v6, Txz8v6, Ayz8v6, Hyz8v6, Oyz8v6;
wire Vyz8v6, Czz8v6, Jzz8v6, Qzz8v6, Xzz8v6, E009v6, L009v6, S009v6, Z009v6, G109v6;
wire N109v6, U109v6, B209v6, I209v6, P209v6, W209v6, D309v6, K309v6, R309v6, Y309v6;
wire F409v6, M409v6, T409v6, A509v6, H509v6, O509v6, V509v6, C609v6, J609v6, Q609v6;
wire X609v6, E709v6, L709v6, S709v6, Z709v6, G809v6, N809v6, U809v6, B909v6, I909v6;
wire P909v6, W909v6, Da09v6, Ka09v6, Ra09v6, Ya09v6, Fb09v6, Mb09v6, Tb09v6, Ac09v6;
wire Hc09v6, Oc09v6, Vc09v6, Cd09v6, Jd09v6, Qd09v6, Xd09v6, Ee09v6, Le09v6, Se09v6;
wire Ze09v6, Gf09v6, Nf09v6, Uf09v6, Bg09v6, Ig09v6, Pg09v6, Cnvmv6, Jnvmv6, Qnvmv6;
wire Xnvmv6, Eovmv6, Lovmv6, Sovmv6, Zovmv6, Gpvmv6, Npvmv6, Upvmv6, Bqvmv6, Iqvmv6;
wire Pqvmv6, Wqvmv6, Drvmv6, Krvmv6, Rrvmv6, Yrvmv6, Fsvmv6, Msvmv6, Tsvmv6, Atvmv6;
wire Htvmv6, Otvmv6, Vtvmv6, Cuvmv6, Juvmv6, Quvmv6, Xuvmv6, Evvmv6, Lvvmv6, Svvmv6;
wire Zvvmv6, Gwvmv6, Nwvmv6, Uwvmv6, Bxvmv6, Ixvmv6, Pxvmv6, Wxvmv6, Dyvmv6, Kyvmv6;
wire Ryvmv6, Yyvmv6, Fzvmv6, Mzvmv6, Tzvmv6, A0wmv6, H0wmv6, O0wmv6, V0wmv6, C1wmv6;
wire J1wmv6, Q1wmv6, X1wmv6, E2wmv6, L2wmv6, S2wmv6, Z2wmv6, G3wmv6, N3wmv6, U3wmv6;
wire B4wmv6, I4wmv6, P4wmv6, W4wmv6, D5wmv6, K5wmv6, R5wmv6, Y5wmv6, F6wmv6, M6wmv6;
wire T6wmv6, A7wmv6, H7wmv6, O7wmv6, V7wmv6, C8wmv6, J8wmv6, Q8wmv6, X8wmv6, E9wmv6;
wire L9wmv6, S9wmv6, Z9wmv6, Gawmv6, Nawmv6, Uawmv6, Bbwmv6, Ibwmv6, Pbwmv6, Wbwmv6;
wire Dcwmv6, Kcwmv6, Rcwmv6, Ycwmv6, Fdwmv6, Mdwmv6, Tdwmv6, Aewmv6, Hewmv6, Oewmv6;
wire Vewmv6, Cfwmv6, Jfwmv6, Qfwmv6, Xfwmv6, Egwmv6, Lgwmv6, Sgwmv6, Zgwmv6, Ghwmv6;
wire Nhwmv6, Uhwmv6, Biwmv6, Iiwmv6, Piwmv6, Wiwmv6, Djwmv6, Kjwmv6, Rjwmv6, Yjwmv6;
wire Fkwmv6, Mkwmv6, Tkwmv6, Alwmv6, Hlwmv6, Olwmv6, Vlwmv6, Cmwmv6, Jmwmv6, Qmwmv6;
wire Xmwmv6, Enwmv6, Lnwmv6, Snwmv6, Znwmv6, Gowmv6, Nowmv6, Uowmv6, Bpwmv6, Ipwmv6;
wire Ppwmv6, Wpwmv6, Dqwmv6, Kqwmv6, Rqwmv6, Yqwmv6, Frwmv6, Mrwmv6, Trwmv6, Aswmv6;
wire Hswmv6, Oswmv6, Vswmv6, Ctwmv6, Jtwmv6, Qtwmv6, Xtwmv6, Euwmv6, Luwmv6, Suwmv6;
wire Zuwmv6, Gvwmv6, Nvwmv6, Uvwmv6, Bwwmv6, Iwwmv6, Pwwmv6, Wwwmv6, Dxwmv6, Kxwmv6;
wire Rxwmv6, Yxwmv6, Fywmv6, Mywmv6, Tywmv6, Azwmv6, Hzwmv6, Ozwmv6, Vzwmv6, C0xmv6;
wire J0xmv6, Q0xmv6, X0xmv6, E1xmv6, L1xmv6, S1xmv6, Z1xmv6, G2xmv6, N2xmv6, U2xmv6;
wire B3xmv6, I3xmv6, P3xmv6, W3xmv6, D4xmv6, K4xmv6, R4xmv6, Y4xmv6, F5xmv6, M5xmv6;
wire T5xmv6, A6xmv6, H6xmv6, O6xmv6, V6xmv6, C7xmv6, J7xmv6, Q7xmv6, X7xmv6, E8xmv6;
wire L8xmv6, S8xmv6, Z8xmv6, G9xmv6, N9xmv6, U9xmv6, Baxmv6, Iaxmv6, Paxmv6, Waxmv6;
wire Dbxmv6, Kbxmv6, Rbxmv6, Ybxmv6, Fcxmv6, Mcxmv6, Tcxmv6, Adxmv6, Hdxmv6, Odxmv6;
wire Vdxmv6, Cexmv6, Jexmv6, Qexmv6, Xexmv6, Efxmv6, Lfxmv6, Sfxmv6, Zfxmv6, Ggxmv6;
wire Ngxmv6, Ugxmv6, Bhxmv6, Ihxmv6, Phxmv6, Whxmv6, Dixmv6, Kixmv6, Rixmv6, Yixmv6;
wire Fjxmv6, Mjxmv6, Tjxmv6, Akxmv6, Hkxmv6, Okxmv6, Vkxmv6, Clxmv6, Jlxmv6, Qlxmv6;
wire Xlxmv6, Emxmv6, Lmxmv6, Smxmv6, Zmxmv6, Gnxmv6, Nnxmv6, Unxmv6, Boxmv6, Ioxmv6;
wire Poxmv6, Woxmv6, Dpxmv6, Kpxmv6, Rpxmv6, Ypxmv6, Fqxmv6, Mqxmv6, Tqxmv6, Arxmv6;
wire Hrxmv6, Orxmv6, Vrxmv6, Csxmv6, Jsxmv6, Qsxmv6, Xsxmv6, Etxmv6, Ltxmv6, Stxmv6;
wire Ztxmv6, Guxmv6, Nuxmv6, Uuxmv6, Bvxmv6, Ivxmv6, Pvxmv6, Wvxmv6, Dwxmv6, Kwxmv6;
wire Rwxmv6, Ywxmv6, Fxxmv6, Mxxmv6, Txxmv6, Ayxmv6, Hyxmv6, Oyxmv6, Vyxmv6, Czxmv6;
wire Jzxmv6, Qzxmv6, Xzxmv6, E0ymv6, L0ymv6, S0ymv6, Z0ymv6, G1ymv6, N1ymv6, U1ymv6;
wire B2ymv6, I2ymv6, P2ymv6, W2ymv6, D3ymv6, K3ymv6, R3ymv6, Y3ymv6, F4ymv6, M4ymv6;
wire T4ymv6, A5ymv6, H5ymv6, O5ymv6, V5ymv6, C6ymv6, J6ymv6, Q6ymv6, X6ymv6, E7ymv6;
wire L7ymv6, S7ymv6, Z7ymv6, G8ymv6, N8ymv6, U8ymv6, B9ymv6, I9ymv6, P9ymv6, W9ymv6;
wire Daymv6, Kaymv6, Raymv6, Yaymv6, Fbymv6, Mbymv6, Tbymv6, Acymv6, Hcymv6, Ocymv6;
wire Vcymv6, Cdymv6, Jdymv6, Qdymv6, Xdymv6, Eeymv6, Leymv6, Seymv6, Zeymv6, Gfymv6;
wire Nfymv6, Ufymv6, Bgymv6, Igymv6, Pgymv6, Wgymv6, Dhymv6, Khymv6, Rhymv6, Yhymv6;
wire Fiymv6, Miymv6, Tiymv6, Ajymv6, Hjymv6, Ojymv6, Vjymv6, Ckymv6, Jkymv6, Qkymv6;
wire Xkymv6, Elymv6, Llymv6, Slymv6, Zlymv6, Gmymv6, Nmymv6, Umymv6, Bnymv6, Inymv6;
wire Pnymv6, Wnymv6, Doymv6, Koymv6, Roymv6, Yoymv6, Fpymv6, Mpymv6, Tpymv6, Aqymv6;
wire Hqymv6, Oqymv6, Vqymv6, Crymv6, Jrymv6, Qrymv6, Xrymv6, Esymv6, Lsymv6, Ssymv6;
wire Zsymv6, Gtymv6, Ntymv6, Utymv6, Buymv6, Iuymv6, Puymv6, Wuymv6, Dvymv6, Kvymv6;
wire Rvymv6, Yvymv6, Fwymv6, Mwymv6, Twymv6, Axymv6, Hxymv6, Oxymv6, Vxymv6, Cyymv6;
wire Jyymv6, Qyymv6, Xyymv6, Ezymv6, Lzymv6, Szymv6, Zzymv6, G0zmv6, N0zmv6, U0zmv6;
wire B1zmv6, I1zmv6, P1zmv6, W1zmv6, D2zmv6, K2zmv6, R2zmv6, Y2zmv6, F3zmv6, M3zmv6;
wire T3zmv6, A4zmv6, H4zmv6, O4zmv6, V4zmv6, C5zmv6, J5zmv6, Q5zmv6, X5zmv6, E6zmv6;
wire L6zmv6, S6zmv6, Z6zmv6, G7zmv6, N7zmv6, U7zmv6, B8zmv6, I8zmv6, P8zmv6, W8zmv6;
wire D9zmv6, K9zmv6, R9zmv6, Y9zmv6, Fazmv6, Mazmv6, Tazmv6, Abzmv6, Hbzmv6, Obzmv6;
wire Vbzmv6, Cczmv6, Jczmv6, Qczmv6, Xczmv6, Edzmv6, Ldzmv6, Sdzmv6, Zdzmv6, Gezmv6;
wire Nezmv6, Uezmv6, Bfzmv6, Ifzmv6, Pfzmv6, Wfzmv6, Dgzmv6, Kgzmv6, Rgzmv6, Ygzmv6;
wire Fhzmv6, Mhzmv6, Thzmv6, Aizmv6, Hizmv6, Oizmv6, Vizmv6, Cjzmv6, Jjzmv6, Qjzmv6;
wire Xjzmv6, Ekzmv6, Lkzmv6, Skzmv6, Zkzmv6, Glzmv6, Nlzmv6, Ulzmv6, Bmzmv6, Imzmv6;
wire Pmzmv6, Wmzmv6, Dnzmv6, Knzmv6, Rnzmv6, Ynzmv6, Fozmv6, Mozmv6, Tozmv6, Apzmv6;
wire Hpzmv6, Opzmv6, Vpzmv6, Cqzmv6, Jqzmv6, Qqzmv6, Xqzmv6, Erzmv6, Lrzmv6, Srzmv6;
wire Zrzmv6, Gszmv6, Nszmv6, Uszmv6, Btzmv6, Itzmv6, Ptzmv6, Wtzmv6, Duzmv6, Kuzmv6;
wire Ruzmv6, Yuzmv6, Fvzmv6, Mvzmv6, Tvzmv6, Awzmv6, Hwzmv6, Owzmv6, Vwzmv6, Cxzmv6;
wire Jxzmv6, Qxzmv6, Xxzmv6, Eyzmv6, Lyzmv6, Syzmv6, Zyzmv6, Gzzmv6, Nzzmv6, Uzzmv6;
wire B00nv6, I00nv6, P00nv6, W00nv6, D10nv6, K10nv6, R10nv6, Y10nv6, F20nv6, M20nv6;
wire T20nv6, A30nv6, H30nv6, O30nv6, V30nv6, C40nv6, J40nv6, Q40nv6, X40nv6, E50nv6;
wire L50nv6, S50nv6, Z50nv6, G60nv6, N60nv6, U60nv6, B70nv6, I70nv6, P70nv6, W70nv6;
wire D80nv6, K80nv6, R80nv6, Y80nv6, F90nv6, M90nv6, T90nv6, Aa0nv6, Ha0nv6, Oa0nv6;
wire Va0nv6, Cb0nv6, Jb0nv6, Qb0nv6, Xb0nv6, Ec0nv6, Lc0nv6, Sc0nv6, Zc0nv6, Gd0nv6;
wire Nd0nv6, Ud0nv6, Be0nv6, Ie0nv6, Pe0nv6, We0nv6, Df0nv6, Kf0nv6, Rf0nv6, Yf0nv6;
wire Fg0nv6, Mg0nv6, Tg0nv6, Ah0nv6, Hh0nv6, Oh0nv6, Vh0nv6, Ci0nv6, Ji0nv6, Qi0nv6;
wire Xi0nv6, Ej0nv6, Lj0nv6, Sj0nv6, Zj0nv6, Gk0nv6, Nk0nv6, Uk0nv6, Bl0nv6, Il0nv6;
wire Pl0nv6, Wl0nv6, Dm0nv6, Km0nv6, Rm0nv6, Ym0nv6, Fn0nv6, Mn0nv6, Tn0nv6, Ao0nv6;
wire Ho0nv6, Oo0nv6, Vo0nv6, Cp0nv6, Jp0nv6, Qp0nv6, Xp0nv6, Eq0nv6, Lq0nv6, Sq0nv6;
wire Zq0nv6, Gr0nv6, Nr0nv6, Ur0nv6, Bs0nv6, Is0nv6, Ps0nv6, Ws0nv6, Dt0nv6, Kt0nv6;
wire Rt0nv6, Yt0nv6, Fu0nv6, Mu0nv6, Tu0nv6, Av0nv6, Hv0nv6, Ov0nv6, Vv0nv6, Cw0nv6;
wire Jw0nv6, Qw0nv6, Xw0nv6, Ex0nv6, Lx0nv6, Sx0nv6, Zx0nv6, Gy0nv6, Ny0nv6, Uy0nv6;
wire Bz0nv6, Iz0nv6, Pz0nv6, Wz0nv6, D01nv6, K01nv6, R01nv6, Y01nv6, F11nv6, M11nv6;
wire T11nv6, A21nv6, H21nv6, O21nv6, V21nv6, C31nv6, J31nv6, Q31nv6, X31nv6, E41nv6;
wire L41nv6, S41nv6, Z41nv6, G51nv6, N51nv6, U51nv6, B61nv6, I61nv6, P61nv6, W61nv6;
wire D71nv6, K71nv6, R71nv6, Y71nv6, F81nv6, M81nv6, T81nv6, A91nv6, H91nv6, O91nv6;
wire V91nv6, Ca1nv6, Ja1nv6, Qa1nv6, Xa1nv6, Eb1nv6, Lb1nv6, Sb1nv6, Zb1nv6, Gc1nv6;
wire Nc1nv6, Uc1nv6, Bd1nv6, Id1nv6, Pd1nv6, Wd1nv6, De1nv6, Ke1nv6, Re1nv6, Ye1nv6;
wire Ff1nv6, Mf1nv6, Tf1nv6, Ag1nv6, Hg1nv6, Og1nv6, Vg1nv6, Ch1nv6, Jh1nv6, Qh1nv6;
wire Xh1nv6, Ei1nv6, Li1nv6, Si1nv6, Zi1nv6, Gj1nv6, Nj1nv6, Uj1nv6, Bk1nv6, Ik1nv6;
wire Pk1nv6, Wk1nv6, Dl1nv6, Kl1nv6, Rl1nv6, Yl1nv6, Fm1nv6, Mm1nv6, Tm1nv6, An1nv6;
wire Hn1nv6, On1nv6, Vn1nv6, Co1nv6, Jo1nv6, Qo1nv6, Xo1nv6, Ep1nv6, Lp1nv6, Sp1nv6;
wire Zp1nv6, Gq1nv6, Nq1nv6, Uq1nv6, Br1nv6, Ir1nv6, Pr1nv6, Wr1nv6, Ds1nv6, Ks1nv6;
wire Rs1nv6, Ys1nv6, Ft1nv6, Mt1nv6, Tt1nv6, Au1nv6, Hu1nv6, Ou1nv6, Vu1nv6, Cv1nv6;
wire Jv1nv6, Qv1nv6, Xv1nv6, Ew1nv6, Lw1nv6, Sw1nv6, Zw1nv6, Gx1nv6, Nx1nv6, Ux1nv6;
wire By1nv6, Iy1nv6, Py1nv6, Wy1nv6, Dz1nv6, Kz1nv6, Rz1nv6, Yz1nv6, F02nv6, M02nv6;
wire T02nv6, A12nv6, H12nv6, O12nv6, V12nv6, C22nv6, J22nv6, Q22nv6, X22nv6, E32nv6;
wire L32nv6, S32nv6, Z32nv6, G42nv6, N42nv6, U42nv6, B52nv6, I52nv6, P52nv6, W52nv6;
wire D62nv6, K62nv6, R62nv6, Y62nv6, F72nv6, M72nv6, T72nv6, A82nv6, H82nv6, O82nv6;
wire V82nv6, C92nv6, J92nv6, Q92nv6, X92nv6, Ea2nv6, La2nv6, Sa2nv6, Za2nv6, Gb2nv6;
wire Nb2nv6, Ub2nv6, Bc2nv6, Ic2nv6, Pc2nv6, Wc2nv6, Dd2nv6, Kd2nv6, Rd2nv6, Yd2nv6;
wire Fe2nv6, Me2nv6, Te2nv6, Af2nv6, Hf2nv6, Of2nv6, Vf2nv6, Cg2nv6, Jg2nv6, Qg2nv6;
wire Xg2nv6, Eh2nv6, Lh2nv6, Sh2nv6, Zh2nv6, Gi2nv6, Ni2nv6, Ui2nv6, Bj2nv6, Ij2nv6;
wire Pj2nv6, Wj2nv6, Dk2nv6, Kk2nv6, Rk2nv6, Yk2nv6, Fl2nv6, Ml2nv6, Tl2nv6, Am2nv6;
wire Hm2nv6, Om2nv6, Vm2nv6, Cn2nv6, Jn2nv6, Qn2nv6, Xn2nv6, Eo2nv6, Lo2nv6, So2nv6;
wire Zo2nv6, Gp2nv6, Np2nv6, Up2nv6, Bq2nv6, Iq2nv6, Pq2nv6, Wq2nv6, Dr2nv6, Kr2nv6;
wire Rr2nv6, Yr2nv6, Fs2nv6, Ms2nv6, Ts2nv6, At2nv6, Ht2nv6, Ot2nv6, Vt2nv6, Cu2nv6;
wire Ju2nv6, Qu2nv6, Xu2nv6, Ev2nv6, Lv2nv6, Sv2nv6, Zv2nv6, Gw2nv6, Nw2nv6, Uw2nv6;
wire Bx2nv6, Ix2nv6, Px2nv6, Wx2nv6, Dy2nv6, Ky2nv6, Ry2nv6, Yy2nv6, Fz2nv6, Mz2nv6;
wire Tz2nv6, A03nv6, H03nv6, O03nv6, V03nv6, C13nv6, J13nv6, Q13nv6, X13nv6, E23nv6;
wire L23nv6, S23nv6, Z23nv6, G33nv6, N33nv6, U33nv6, B43nv6, I43nv6, P43nv6, W43nv6;
wire D53nv6, K53nv6, R53nv6, Y53nv6, F63nv6, M63nv6, T63nv6, A73nv6, H73nv6, O73nv6;
wire V73nv6, C83nv6, J83nv6, Q83nv6, X83nv6, E93nv6, L93nv6, S93nv6, Z93nv6, Ga3nv6;
wire Na3nv6, Ua3nv6, Bb3nv6, Ib3nv6, Pb3nv6, Wb3nv6, Dc3nv6, Kc3nv6, Rc3nv6, Yc3nv6;
wire Fd3nv6, Md3nv6, Td3nv6, Ae3nv6, He3nv6, Oe3nv6, Ve3nv6, Cf3nv6, Jf3nv6, Qf3nv6;
wire Xf3nv6, Eg3nv6, Lg3nv6, Sg3nv6, Zg3nv6, Gh3nv6, Nh3nv6, Uh3nv6, Bi3nv6, Ii3nv6;
wire Pi3nv6, Wi3nv6, Dj3nv6, Kj3nv6, Rj3nv6, Yj3nv6, Fk3nv6, Mk3nv6, Tk3nv6, Al3nv6;
wire Hl3nv6, Ol3nv6, Vl3nv6, Cm3nv6, Jm3nv6, Qm3nv6, Xm3nv6, En3nv6, Ln3nv6, Sn3nv6;
wire Zn3nv6, Go3nv6, No3nv6, Uo3nv6, Bp3nv6, Ip3nv6, Pp3nv6, Wp3nv6, Dq3nv6, Kq3nv6;
wire Rq3nv6, Yq3nv6, Fr3nv6, Mr3nv6, Tr3nv6, As3nv6, Hs3nv6, Os3nv6, Vs3nv6, Ct3nv6;
wire Jt3nv6, Qt3nv6, Xt3nv6, Eu3nv6, Lu3nv6, Su3nv6, Zu3nv6, Gv3nv6, Nv3nv6, Uv3nv6;
wire Bw3nv6, Iw3nv6, Pw3nv6, Ww3nv6, Dx3nv6, Kx3nv6, Rx3nv6, Yx3nv6, Fy3nv6, My3nv6;
wire Ty3nv6, Az3nv6, Hz3nv6, Oz3nv6, Vz3nv6, C04nv6, J04nv6, Q04nv6, X04nv6, E14nv6;
wire L14nv6, S14nv6, Z14nv6, G24nv6, N24nv6, U24nv6, B34nv6, I34nv6, P34nv6, W34nv6;
wire D44nv6, K44nv6, R44nv6, Y44nv6, F54nv6, M54nv6, T54nv6, A64nv6, H64nv6, O64nv6;
wire V64nv6, C74nv6, J74nv6, Q74nv6, X74nv6, E84nv6, L84nv6, S84nv6, Z84nv6, G94nv6;
wire N94nv6, U94nv6, Ba4nv6, Ia4nv6, Pa4nv6, Wa4nv6, Db4nv6, Kb4nv6, Rb4nv6, Yb4nv6;
wire Fc4nv6, Mc4nv6, Tc4nv6, Ad4nv6, Hd4nv6, Od4nv6, Vd4nv6, Ce4nv6, Je4nv6, Qe4nv6;
wire Xe4nv6, Ef4nv6, Lf4nv6, Sf4nv6, Zf4nv6, Gg4nv6, Ng4nv6, Ug4nv6, Bh4nv6, Ih4nv6;
wire Ph4nv6, Wh4nv6, Di4nv6, Ki4nv6, Ri4nv6, Yi4nv6, Fj4nv6, Mj4nv6, Tj4nv6, Ak4nv6;
wire Hk4nv6, Ok4nv6, Vk4nv6, Cl4nv6, Jl4nv6, Ql4nv6, Xl4nv6, Em4nv6, Lm4nv6, Sm4nv6;
wire Zm4nv6, Gn4nv6, Nn4nv6, Un4nv6, Bo4nv6, Io4nv6, Po4nv6, Wo4nv6, Dp4nv6, Kp4nv6;
wire Rp4nv6, Yp4nv6, Fq4nv6, Mq4nv6, Tq4nv6, Ar4nv6, Hr4nv6, Or4nv6, Vr4nv6, Cs4nv6;
wire Js4nv6, Qs4nv6, Xs4nv6, Et4nv6, Lt4nv6, St4nv6, Zt4nv6, Gu4nv6, Nu4nv6, Uu4nv6;
wire Bv4nv6, Iv4nv6, Pv4nv6, Wv4nv6, Dw4nv6, Kw4nv6, Rw4nv6, Yw4nv6, Fx4nv6, Mx4nv6;
wire Tx4nv6, Ay4nv6, Hy4nv6, Oy4nv6, Vy4nv6, Cz4nv6, Jz4nv6, Qz4nv6, Xz4nv6, E05nv6;
wire L05nv6, S05nv6, Z05nv6, G15nv6, N15nv6, U15nv6, B25nv6, I25nv6, P25nv6, W25nv6;
wire D35nv6, K35nv6, R35nv6, Y35nv6, F45nv6, M45nv6, T45nv6, A55nv6, H55nv6, O55nv6;
wire V55nv6, C65nv6, J65nv6, Q65nv6, X65nv6, E75nv6, L75nv6, S75nv6, Z75nv6, G85nv6;
wire N85nv6, U85nv6, B95nv6, I95nv6, P95nv6, W95nv6, Da5nv6, Ka5nv6, Ra5nv6, Ya5nv6;
wire Fb5nv6, Mb5nv6, Tb5nv6, Ac5nv6, Hc5nv6, Oc5nv6, Vc5nv6, Cd5nv6, Jd5nv6, Qd5nv6;
wire Xd5nv6, Ee5nv6, Le5nv6, Se5nv6, Ze5nv6, Gf5nv6, Nf5nv6, Uf5nv6, Bg5nv6, Ig5nv6;
wire Pg5nv6, Wg5nv6, Dh5nv6, Kh5nv6, Rh5nv6, Yh5nv6, Fi5nv6, Mi5nv6, Ti5nv6, Aj5nv6;
wire Hj5nv6, Oj5nv6, Vj5nv6, Ck5nv6, Jk5nv6, Qk5nv6, Xk5nv6, El5nv6, Ll5nv6, Sl5nv6;
wire Zl5nv6, Gm5nv6, Nm5nv6, Um5nv6, Bn5nv6, In5nv6, Pn5nv6, Wn5nv6, Do5nv6, Ko5nv6;
wire Ro5nv6, Yo5nv6, Fp5nv6, Mp5nv6, Tp5nv6, Aq5nv6, Hq5nv6, Oq5nv6, Vq5nv6, Cr5nv6;
wire Jr5nv6, Qr5nv6, Xr5nv6, Es5nv6, Ls5nv6, Ss5nv6, Zs5nv6, Gt5nv6, Nt5nv6, Ut5nv6;
wire Bu5nv6, Iu5nv6, Pu5nv6, Wu5nv6, Dv5nv6, Kv5nv6, Rv5nv6, Yv5nv6, Fw5nv6, Mw5nv6;
wire Tw5nv6, Ax5nv6, Hx5nv6, Ox5nv6, Vx5nv6, Cy5nv6, Jy5nv6, Qy5nv6, Xy5nv6, Ez5nv6;
wire Lz5nv6, Sz5nv6, Zz5nv6, G06nv6, N06nv6, U06nv6, B16nv6, I16nv6, P16nv6, W16nv6;
wire D26nv6, K26nv6, R26nv6, Y26nv6, F36nv6, M36nv6, T36nv6, A46nv6, H46nv6, O46nv6;
wire V46nv6, C56nv6, J56nv6, Q56nv6, X56nv6, E66nv6, L66nv6, S66nv6, Z66nv6, G76nv6;
wire N76nv6, U76nv6, B86nv6, I86nv6, P86nv6, W86nv6, D96nv6, K96nv6, R96nv6, Y96nv6;
wire Fa6nv6, Ma6nv6, Ta6nv6, Ab6nv6, Hb6nv6, Ob6nv6, Vb6nv6, Cc6nv6, Jc6nv6, Qc6nv6;
wire Xc6nv6, Ed6nv6, Ld6nv6, Sd6nv6, Zd6nv6, Ge6nv6, Ne6nv6, Ue6nv6, Bf6nv6, If6nv6;
wire Pf6nv6, Wf6nv6, Dg6nv6, Kg6nv6, Rg6nv6, Yg6nv6, Fh6nv6, Mh6nv6, Th6nv6, Ai6nv6;
wire Hi6nv6, Oi6nv6, Vi6nv6, Cj6nv6, Jj6nv6, Qj6nv6, Xj6nv6, Ek6nv6, Lk6nv6, Sk6nv6;
wire Zk6nv6, Gl6nv6, Nl6nv6, Ul6nv6, Bm6nv6, Im6nv6, Pm6nv6, Wm6nv6, Dn6nv6, Kn6nv6;
wire Rn6nv6, Yn6nv6, Fo6nv6, Mo6nv6, To6nv6, Ap6nv6, Hp6nv6, Op6nv6, Vp6nv6, Cq6nv6;
wire Jq6nv6, Qq6nv6, Xq6nv6, Er6nv6, Lr6nv6, Sr6nv6, Zr6nv6, Gs6nv6, Ns6nv6, Us6nv6;
wire Bt6nv6, It6nv6, Pt6nv6, Wt6nv6, Du6nv6, Ku6nv6, Ru6nv6, Yu6nv6, Fv6nv6, Mv6nv6;
wire Tv6nv6, Aw6nv6, Hw6nv6, Ow6nv6, Vw6nv6, Cx6nv6, Jx6nv6, Qx6nv6, Xx6nv6, Ey6nv6;
wire Ly6nv6, Sy6nv6, Zy6nv6, Gz6nv6, Nz6nv6, Uz6nv6, B07nv6, I07nv6, P07nv6, W07nv6;
wire D17nv6, K17nv6, R17nv6, Y17nv6, F27nv6, M27nv6, T27nv6, A37nv6, H37nv6, O37nv6;
wire V37nv6, C47nv6, J47nv6, Q47nv6, X47nv6, E57nv6, L57nv6, S57nv6, Z57nv6, G67nv6;
wire N67nv6, U67nv6, B77nv6, I77nv6, P77nv6, W77nv6, D87nv6, K87nv6, R87nv6, Y87nv6;
wire F97nv6, M97nv6, T97nv6, Aa7nv6, Ha7nv6, Oa7nv6, Va7nv6, Cb7nv6, Jb7nv6, Qb7nv6;
wire Xb7nv6, Ec7nv6, Lc7nv6, Sc7nv6, Zc7nv6, Gd7nv6, Nd7nv6, Ud7nv6, Be7nv6, Ie7nv6;
wire Pe7nv6, We7nv6, Df7nv6, Kf7nv6, Rf7nv6, Yf7nv6, Fg7nv6, Mg7nv6, Tg7nv6, Ah7nv6;
wire Hh7nv6, Oh7nv6, Vh7nv6, Ci7nv6, Ji7nv6, Qi7nv6, Xi7nv6, Ej7nv6, Lj7nv6, Sj7nv6;
wire Zj7nv6, Gk7nv6, Nk7nv6, Uk7nv6, Bl7nv6, Il7nv6, Pl7nv6, Wl7nv6, Dm7nv6, Km7nv6;
wire Rm7nv6, Ym7nv6, Fn7nv6, Mn7nv6, Tn7nv6, Ao7nv6, Ho7nv6, Oo7nv6, Vo7nv6, Cp7nv6;
wire Jp7nv6, Qp7nv6, Xp7nv6, Eq7nv6, Lq7nv6, Sq7nv6, Zq7nv6, Gr7nv6, Nr7nv6, Ur7nv6;
wire Bs7nv6, Is7nv6, Ps7nv6, Ws7nv6, Dt7nv6, Kt7nv6, Rt7nv6, Yt7nv6, Fu7nv6, Mu7nv6;
wire Tu7nv6, Av7nv6, Hv7nv6, Ov7nv6, Vv7nv6, Cw7nv6, Jw7nv6, Qw7nv6, Xw7nv6, Ex7nv6;
wire Lx7nv6, Sx7nv6, Zx7nv6, Gy7nv6, Ny7nv6, Uy7nv6, Bz7nv6, Iz7nv6, Pz7nv6, Wz7nv6;
wire D08nv6, K08nv6, R08nv6, Y08nv6, F18nv6, M18nv6, T18nv6, A28nv6, H28nv6, O28nv6;
wire V28nv6, C38nv6, J38nv6, Q38nv6, X38nv6, E48nv6, L48nv6, S48nv6, Z48nv6, G58nv6;
wire N58nv6, U58nv6, B68nv6, I68nv6, P68nv6, W68nv6, D78nv6, K78nv6, R78nv6, Y78nv6;
wire F88nv6, M88nv6, T88nv6, A98nv6, H98nv6, O98nv6, V98nv6, Ca8nv6, Ja8nv6, Qa8nv6;
wire Xa8nv6, Eb8nv6, Lb8nv6, Sb8nv6, Zb8nv6, Gc8nv6, Nc8nv6, Uc8nv6, Bd8nv6, Id8nv6;
wire Pd8nv6, Wd8nv6, De8nv6, Ke8nv6, Re8nv6, Ye8nv6, Ff8nv6, Mf8nv6, Tf8nv6, Ag8nv6;
wire Hg8nv6, Og8nv6, Vg8nv6, Ch8nv6, Jh8nv6, Qh8nv6, Xh8nv6, Ei8nv6, Li8nv6, Si8nv6;
wire Zi8nv6, Gj8nv6, Nj8nv6, Uj8nv6, Bk8nv6, Ik8nv6, Pk8nv6, Wk8nv6, Dl8nv6, Kl8nv6;
wire Rl8nv6, Yl8nv6, Fm8nv6, Mm8nv6, Tm8nv6, An8nv6, Hn8nv6, On8nv6, Vn8nv6, Co8nv6;
wire Jo8nv6, Qo8nv6, Xo8nv6, Ep8nv6, Lp8nv6, Sp8nv6, Zp8nv6, Gq8nv6, Nq8nv6, Uq8nv6;
wire Br8nv6, Ir8nv6, Pr8nv6, Wr8nv6, Ds8nv6, Ks8nv6, Rs8nv6, Ys8nv6, Ft8nv6, Mt8nv6;
wire Tt8nv6, Au8nv6, Hu8nv6, Ou8nv6, Vu8nv6, Cv8nv6, Jv8nv6, Qv8nv6, Xv8nv6, Ew8nv6;
wire Lw8nv6, Sw8nv6, Zw8nv6, Gx8nv6, Nx8nv6, Ux8nv6, By8nv6, Iy8nv6, Py8nv6, Wy8nv6;
wire Dz8nv6, Kz8nv6, Rz8nv6, Yz8nv6, F09nv6, M09nv6, T09nv6, A19nv6, H19nv6, O19nv6;
wire V19nv6, C29nv6, J29nv6, Q29nv6, X29nv6, E39nv6, L39nv6, S39nv6, Z39nv6, G49nv6;
wire N49nv6, U49nv6, B59nv6, I59nv6, P59nv6, W59nv6, D69nv6, K69nv6, R69nv6, Y69nv6;
wire F79nv6, M79nv6, T79nv6, A89nv6, H89nv6, O89nv6, V89nv6, C99nv6, J99nv6, Q99nv6;
wire X99nv6, Ea9nv6, La9nv6, Sa9nv6, Za9nv6, Gb9nv6, Nb9nv6, Ub9nv6, Bc9nv6, Ic9nv6;
wire Pc9nv6, Wc9nv6, Dd9nv6, Kd9nv6, Rd9nv6, Yd9nv6, Fe9nv6, Me9nv6, Te9nv6, Af9nv6;
wire Hf9nv6, Of9nv6, Vf9nv6, Cg9nv6, Jg9nv6, Qg9nv6, Xg9nv6, Eh9nv6, Lh9nv6, Sh9nv6;
wire Zh9nv6, Gi9nv6, Ni9nv6, Ui9nv6, Bj9nv6, Ij9nv6, Pj9nv6, Wj9nv6, Dk9nv6, Kk9nv6;
wire Rk9nv6, Yk9nv6, Fl9nv6, Ml9nv6, Tl9nv6, Am9nv6, Hm9nv6, Om9nv6, Vm9nv6, Cn9nv6;
wire Jn9nv6, Qn9nv6, Xn9nv6, Eo9nv6, Lo9nv6, So9nv6, Zo9nv6, Gp9nv6, Np9nv6, Up9nv6;
wire Bq9nv6, Iq9nv6, Pq9nv6, Wq9nv6, Dr9nv6, Kr9nv6, Rr9nv6, Yr9nv6, Fs9nv6, Ms9nv6;
wire Ts9nv6, At9nv6, Ht9nv6, Ot9nv6, Vt9nv6, Cu9nv6, Ju9nv6, Qu9nv6, Xu9nv6, Ev9nv6;
wire Lv9nv6, Sv9nv6, Zv9nv6, Gw9nv6, Nw9nv6, Uw9nv6, Bx9nv6, Ix9nv6, Px9nv6, Wx9nv6;
wire Dy9nv6, Ky9nv6, Ry9nv6, Yy9nv6, Fz9nv6, Mz9nv6, Tz9nv6, A0anv6, H0anv6, O0anv6;
wire V0anv6, C1anv6, J1anv6, Q1anv6, X1anv6, E2anv6, L2anv6, S2anv6, Z2anv6, G3anv6;
wire N3anv6, U3anv6, B4anv6, I4anv6, P4anv6, W4anv6, D5anv6, K5anv6, R5anv6, Y5anv6;
wire F6anv6, M6anv6, T6anv6, A7anv6, H7anv6, O7anv6, V7anv6, C8anv6, J8anv6, Q8anv6;
wire X8anv6, E9anv6, L9anv6, S9anv6, Z9anv6, Gaanv6, Naanv6, Uaanv6, Bbanv6, Ibanv6;
wire Pbanv6, Wbanv6, Dcanv6, Kcanv6, Rcanv6, Ycanv6, Fdanv6, Mdanv6, Tdanv6, Aeanv6;
wire Heanv6, Oeanv6, Veanv6, Cfanv6, Jfanv6, Qfanv6, Xfanv6, Eganv6, Lganv6, Sganv6;
wire Zganv6, Ghanv6, Nhanv6, Uhanv6, Bianv6, Iianv6, Pianv6, Wianv6, Djanv6, Kjanv6;
wire Rjanv6, Yjanv6, Fkanv6, Mkanv6, Tkanv6, Alanv6, Hlanv6, Olanv6, Vlanv6, Cmanv6;
wire Jmanv6, Qmanv6, Xmanv6, Enanv6, Lnanv6, Snanv6, Znanv6, Goanv6, Noanv6, Uoanv6;
wire Bpanv6, Ipanv6, Ppanv6, Wpanv6, Dqanv6, Kqanv6, Rqanv6, Yqanv6, Franv6, Mranv6;
wire Tranv6, Asanv6, Hsanv6, Osanv6, Vsanv6, Ctanv6, Jtanv6, Qtanv6, Xtanv6, Euanv6;
wire Luanv6, Suanv6, Zuanv6, Gvanv6, Nvanv6, Uvanv6, Bwanv6, Iwanv6, Pwanv6, Wwanv6;
wire Dxanv6, Kxanv6, Rxanv6, Yxanv6, Fyanv6, Myanv6, Tyanv6, Azanv6, Hzanv6, Ozanv6;
wire Vzanv6, C0bnv6, J0bnv6, Q0bnv6, X0bnv6, E1bnv6, L1bnv6, S1bnv6, Z1bnv6, G2bnv6;
wire N2bnv6, U2bnv6, B3bnv6, I3bnv6, P3bnv6, W3bnv6, D4bnv6, K4bnv6, R4bnv6, Y4bnv6;
wire F5bnv6, M5bnv6, T5bnv6, A6bnv6, H6bnv6, O6bnv6, V6bnv6, C7bnv6, J7bnv6, Q7bnv6;
wire X7bnv6, E8bnv6, L8bnv6, S8bnv6, Z8bnv6, G9bnv6, N9bnv6, U9bnv6, Babnv6, Iabnv6;
wire Pabnv6, Wabnv6, Dbbnv6, Kbbnv6, Rbbnv6, Ybbnv6, Fcbnv6, Mcbnv6, Tcbnv6, Adbnv6;
wire Hdbnv6, Odbnv6, Vdbnv6, Cebnv6, Jebnv6, Qebnv6, Xebnv6, Efbnv6, Lfbnv6, Sfbnv6;
wire Zfbnv6, Ggbnv6, Ngbnv6, Ugbnv6, Bhbnv6, Ihbnv6, Phbnv6, Whbnv6, Dibnv6, Kibnv6;
wire Ribnv6, Yibnv6, Fjbnv6, Mjbnv6, Tjbnv6, Akbnv6, Hkbnv6, Okbnv6, Vkbnv6, Clbnv6;
wire Jlbnv6, Qlbnv6, Xlbnv6, Embnv6, Lmbnv6, Smbnv6, Zmbnv6, Gnbnv6, Nnbnv6, Unbnv6;
wire Bobnv6, Iobnv6, Pobnv6, Wobnv6, Dpbnv6, Kpbnv6, Rpbnv6, Ypbnv6, Fqbnv6, Mqbnv6;
wire Tqbnv6, Arbnv6, Hrbnv6, Orbnv6, Vrbnv6, Csbnv6, Jsbnv6, Qsbnv6, Xsbnv6, Etbnv6;
wire Ltbnv6, Stbnv6, Ztbnv6, Gubnv6, Nubnv6, Uubnv6, Bvbnv6, Ivbnv6, Pvbnv6, Wvbnv6;
wire Dwbnv6, Kwbnv6, Rwbnv6, Ywbnv6, Fxbnv6, Mxbnv6, Txbnv6, Aybnv6, Hybnv6, Oybnv6;
wire Vybnv6, Czbnv6, Jzbnv6, Qzbnv6, Xzbnv6, E0cnv6, L0cnv6, S0cnv6, Z0cnv6, G1cnv6;
wire N1cnv6, U1cnv6, B2cnv6, I2cnv6, P2cnv6, W2cnv6, D3cnv6, K3cnv6, R3cnv6, Y3cnv6;
wire F4cnv6, M4cnv6, T4cnv6, A5cnv6, H5cnv6, O5cnv6, V5cnv6, C6cnv6, J6cnv6, Q6cnv6;
wire X6cnv6, E7cnv6, L7cnv6, S7cnv6, Z7cnv6, G8cnv6, N8cnv6, U8cnv6, B9cnv6, I9cnv6;
wire P9cnv6, W9cnv6, Dacnv6, Kacnv6, Racnv6, Yacnv6, Fbcnv6, Mbcnv6, Tbcnv6, Accnv6;
wire Hccnv6, Occnv6, Vccnv6, Cdcnv6, Jdcnv6, Qdcnv6, Xdcnv6, Eecnv6, Lecnv6, Secnv6;
wire Zecnv6, Gfcnv6, Nfcnv6, Ufcnv6, Bgcnv6, Igcnv6, Pgcnv6, Wgcnv6, Dhcnv6, Khcnv6;
wire Rhcnv6, Yhcnv6, Ficnv6, Micnv6, Ticnv6, Ajcnv6, Hjcnv6, Ojcnv6, Vjcnv6, Ckcnv6;
wire Jkcnv6, Qkcnv6, Xkcnv6, Elcnv6, Llcnv6, Slcnv6, Zlcnv6, Gmcnv6, Nmcnv6, Umcnv6;
wire Bncnv6, Incnv6, Pncnv6, Wncnv6, Docnv6, Kocnv6, Rocnv6, Yocnv6, Fpcnv6, Mpcnv6;
wire Tpcnv6, Aqcnv6, Hqcnv6, Oqcnv6, Vqcnv6, Crcnv6, Jrcnv6, Qrcnv6, Xrcnv6, Escnv6;
wire Lscnv6, Sscnv6, Zscnv6, Gtcnv6, Ntcnv6, Utcnv6, Bucnv6, Iucnv6, Pucnv6, Wucnv6;
wire Dvcnv6, Kvcnv6, Rvcnv6, Yvcnv6, Fwcnv6, Mwcnv6, Twcnv6, Axcnv6, Hxcnv6, Oxcnv6;
wire Vxcnv6, Cycnv6, Jycnv6, Qycnv6, Xycnv6, Ezcnv6, Lzcnv6, Szcnv6, Zzcnv6, G0dnv6;
wire N0dnv6, U0dnv6, B1dnv6, I1dnv6, P1dnv6, W1dnv6, D2dnv6, K2dnv6, R2dnv6, Y2dnv6;
wire F3dnv6, M3dnv6, T3dnv6, A4dnv6, H4dnv6, O4dnv6, V4dnv6, C5dnv6, J5dnv6, Q5dnv6;
wire X5dnv6, E6dnv6, L6dnv6, S6dnv6, Z6dnv6, G7dnv6, N7dnv6, U7dnv6, B8dnv6, I8dnv6;
wire P8dnv6, W8dnv6, D9dnv6, K9dnv6, R9dnv6, Y9dnv6, Fadnv6, Madnv6, Tadnv6, Abdnv6;
wire Hbdnv6, Obdnv6, Vbdnv6, Ccdnv6, Jcdnv6, Qcdnv6, Xcdnv6, Eddnv6, Lddnv6, Sddnv6;
wire Zddnv6, Gednv6, Nednv6, Uednv6, Bfdnv6, Ifdnv6, Pfdnv6, Wfdnv6, Dgdnv6, Kgdnv6;
wire Rgdnv6, Ygdnv6, Fhdnv6, Mhdnv6, Thdnv6, Aidnv6, Hidnv6, Oidnv6, Vidnv6, Cjdnv6;
wire Jjdnv6, Qjdnv6, Xjdnv6, Ekdnv6, Lkdnv6, Skdnv6, Zkdnv6, Gldnv6, Nldnv6, Uldnv6;
wire Bmdnv6, Imdnv6, Pmdnv6, Wmdnv6, Dndnv6, Kndnv6, Rndnv6, Yndnv6, Fodnv6, Modnv6;
wire Todnv6, Apdnv6, Hpdnv6, Opdnv6, Vpdnv6, Cqdnv6, Jqdnv6, Qqdnv6, Xqdnv6, Erdnv6;
wire Lrdnv6, Srdnv6, Zrdnv6, Gsdnv6, Nsdnv6, Usdnv6, Btdnv6, Itdnv6, Ptdnv6, Wtdnv6;
wire Dudnv6, Kudnv6, Rudnv6, Yudnv6, Fvdnv6, Mvdnv6, Tvdnv6, Awdnv6, Hwdnv6, Owdnv6;
wire Vwdnv6, Cxdnv6, Jxdnv6, Qxdnv6, Xxdnv6, Eydnv6, Lydnv6, Sydnv6, Zydnv6, Gzdnv6;
wire Nzdnv6, Uzdnv6, B0env6, I0env6, P0env6, W0env6, D1env6, K1env6, R1env6, Y1env6;
wire F2env6, M2env6, T2env6, A3env6, H3env6, O3env6, V3env6, C4env6, J4env6, Q4env6;
wire X4env6, E5env6, L5env6, S5env6, Z5env6, G6env6, N6env6, U6env6, B7env6, I7env6;
wire P7env6, W7env6, D8env6, K8env6, R8env6, Y8env6, F9env6, M9env6, T9env6, Aaenv6;
wire Haenv6, Oaenv6, Vaenv6, Cbenv6, Jbenv6, Qbenv6, Xbenv6, Ecenv6, Lcenv6, Scenv6;
wire Zcenv6, Gdenv6, Ndenv6, Udenv6, Beenv6, Ieenv6, Peenv6, Weenv6, Dfenv6, Kfenv6;
wire Rfenv6, Yfenv6, Fgenv6, Mgenv6, Tgenv6, Ahenv6, Hhenv6, Ohenv6, Vhenv6, Cienv6;
wire Jienv6, Qienv6, Xienv6, Ejenv6, Ljenv6, Sjenv6, Zjenv6, Gkenv6, Nkenv6, Ukenv6;
wire Blenv6, Ilenv6, Plenv6, Wlenv6, Dmenv6, Kmenv6, Rmenv6, Ymenv6, Fnenv6, Mnenv6;
wire Tnenv6, Aoenv6, Hoenv6, Ooenv6, Voenv6, Cpenv6, Jpenv6, Qpenv6, Xpenv6, Eqenv6;
wire Lqenv6, Sqenv6, Zqenv6, Grenv6, Nrenv6, Urenv6, Bsenv6, Isenv6, Psenv6, Wsenv6;
wire Dtenv6, Ktenv6, Rtenv6, Ytenv6, Fuenv6, Muenv6, Tuenv6, Avenv6, Hvenv6, Ovenv6;
wire Vvenv6, Cwenv6, Jwenv6, Qwenv6, Xwenv6, Exenv6, Lxenv6, Sxenv6, Zxenv6, Gyenv6;
wire Nyenv6, Uyenv6, Bzenv6, Izenv6, Pzenv6, Wzenv6, D0fnv6, K0fnv6, R0fnv6, Y0fnv6;
wire F1fnv6, M1fnv6, T1fnv6, A2fnv6, H2fnv6, O2fnv6, V2fnv6, C3fnv6, J3fnv6, Q3fnv6;
wire X3fnv6, E4fnv6, L4fnv6, S4fnv6, Z4fnv6, G5fnv6, N5fnv6, U5fnv6, B6fnv6, I6fnv6;
wire P6fnv6, W6fnv6, D7fnv6, K7fnv6, R7fnv6, Y7fnv6, F8fnv6, M8fnv6, T8fnv6, A9fnv6;
wire H9fnv6, O9fnv6, V9fnv6, Cafnv6, Jafnv6, Qafnv6, Xafnv6, Ebfnv6, Lbfnv6, Sbfnv6;
wire Zbfnv6, Gcfnv6, Ncfnv6, Ucfnv6, Bdfnv6, Idfnv6, Pdfnv6, Wdfnv6, Defnv6, Kefnv6;
wire Refnv6, Yefnv6, Fffnv6, Mffnv6, Tffnv6, Agfnv6, Hgfnv6, Ogfnv6, Vgfnv6, Chfnv6;
wire Jhfnv6, Qhfnv6, Xhfnv6, Eifnv6, Lifnv6, Sifnv6, Zifnv6, Gjfnv6, Njfnv6, Ujfnv6;
wire Bkfnv6, Ikfnv6, Pkfnv6, Wkfnv6, Dlfnv6, Klfnv6, Rlfnv6, Ylfnv6, Fmfnv6, Mmfnv6;
wire Tmfnv6, Anfnv6, Hnfnv6, Onfnv6, Vnfnv6, Cofnv6, Jofnv6, Qofnv6, Xofnv6, Epfnv6;
wire Lpfnv6, Spfnv6, Zpfnv6, Gqfnv6, Nqfnv6, Uqfnv6, Brfnv6, Irfnv6, Prfnv6, Wrfnv6;
wire Dsfnv6, Ksfnv6, Rsfnv6, Ysfnv6, Ftfnv6, Mtfnv6, Ttfnv6, Aufnv6, Hufnv6, Oufnv6;
wire Vufnv6, Cvfnv6, Jvfnv6, Qvfnv6, Xvfnv6, Ewfnv6, Lwfnv6, Swfnv6, Zwfnv6, Gxfnv6;
wire Nxfnv6, Uxfnv6, Byfnv6, Iyfnv6, Pyfnv6, Wyfnv6, Dzfnv6, Kzfnv6, Rzfnv6, Yzfnv6;
wire F0gnv6, M0gnv6, T0gnv6, A1gnv6, H1gnv6, O1gnv6, V1gnv6, C2gnv6, J2gnv6, Q2gnv6;
wire X2gnv6, E3gnv6, L3gnv6, S3gnv6, Z3gnv6, G4gnv6, N4gnv6, U4gnv6, B5gnv6, I5gnv6;
wire P5gnv6, W5gnv6, D6gnv6, K6gnv6, R6gnv6, Y6gnv6, F7gnv6, M7gnv6, T7gnv6, A8gnv6;
wire H8gnv6, O8gnv6, V8gnv6, C9gnv6, J9gnv6, Q9gnv6, X9gnv6, Eagnv6, Lagnv6, Sagnv6;
wire Zagnv6, Gbgnv6, Nbgnv6, Ubgnv6, Bcgnv6, Icgnv6, Pcgnv6, Wcgnv6, Ddgnv6, Kdgnv6;
wire Rdgnv6, Ydgnv6, Fegnv6, Megnv6, Tegnv6, Afgnv6, Hfgnv6, Ofgnv6, Vfgnv6, Cggnv6;
wire Jggnv6, Qggnv6, Xggnv6, Ehgnv6, Lhgnv6, Shgnv6, Zhgnv6, Gignv6, Nignv6, Uignv6;
wire Bjgnv6, Ijgnv6, Pjgnv6, Wjgnv6, Dkgnv6, Kkgnv6, Rkgnv6, Ykgnv6, Flgnv6, Mlgnv6;
wire Tlgnv6, Amgnv6, Hmgnv6, Omgnv6, Vmgnv6, Cngnv6, Jngnv6, Qngnv6, Xngnv6, Eognv6;
wire Lognv6, Sognv6, Zognv6, Gpgnv6, Npgnv6, Upgnv6, Bqgnv6, Iqgnv6, Pqgnv6, Wqgnv6;
wire Drgnv6, Krgnv6, Rrgnv6, Yrgnv6, Fsgnv6, Msgnv6, Tsgnv6, Atgnv6, Htgnv6, Otgnv6;
wire Vtgnv6, Cugnv6, Jugnv6, Qugnv6, Xugnv6, Evgnv6, Lvgnv6, Svgnv6, Zvgnv6, Gwgnv6;
wire Nwgnv6, Uwgnv6, Bxgnv6, Ixgnv6, Pxgnv6, Wxgnv6, Dygnv6, Kygnv6, Rygnv6, Yygnv6;
wire Fzgnv6, Mzgnv6, Tzgnv6, A0hnv6, H0hnv6, O0hnv6, V0hnv6, C1hnv6, J1hnv6, Q1hnv6;
wire X1hnv6, E2hnv6, L2hnv6, S2hnv6, Z2hnv6, G3hnv6, N3hnv6, U3hnv6, B4hnv6, I4hnv6;
wire P4hnv6, W4hnv6, D5hnv6, K5hnv6, R5hnv6, Y5hnv6, F6hnv6, M6hnv6, T6hnv6, A7hnv6;
wire H7hnv6, O7hnv6, V7hnv6, C8hnv6, J8hnv6, Q8hnv6, X8hnv6, E9hnv6, L9hnv6, S9hnv6;
wire Z9hnv6, Gahnv6, Nahnv6, Uahnv6, Bbhnv6, Ibhnv6, Pbhnv6, Wbhnv6, Dchnv6, Kchnv6;
wire Rchnv6, Ychnv6, Fdhnv6, Mdhnv6, Tdhnv6, Aehnv6, Hehnv6, Oehnv6, Vehnv6, Cfhnv6;
wire Jfhnv6, Qfhnv6, Xfhnv6, Eghnv6, Lghnv6, Sghnv6, Zghnv6, Ghhnv6, Nhhnv6, Uhhnv6;
wire Bihnv6, Iihnv6, Pihnv6, Wihnv6, Djhnv6, Kjhnv6, Rjhnv6, Yjhnv6, Fkhnv6, Mkhnv6;
wire Tkhnv6, Alhnv6, Hlhnv6, Olhnv6, Vlhnv6, Cmhnv6, Jmhnv6, Qmhnv6, Xmhnv6, Enhnv6;
wire Lnhnv6, Snhnv6, Znhnv6, Gohnv6, Nohnv6, Uohnv6, Bphnv6, Iphnv6, Pphnv6, Wphnv6;
wire Dqhnv6, Kqhnv6, Rqhnv6, Yqhnv6, Frhnv6, Mrhnv6, Trhnv6, Ashnv6, Hshnv6, Oshnv6;
wire Vshnv6, Cthnv6, Jthnv6, Qthnv6, Xthnv6, Euhnv6, Luhnv6, Suhnv6, Zuhnv6, Gvhnv6;
wire Nvhnv6, Uvhnv6, Bwhnv6, Iwhnv6, Pwhnv6, Wwhnv6, Dxhnv6, Kxhnv6, Rxhnv6, Yxhnv6;
wire Fyhnv6, Myhnv6, Tyhnv6, Azhnv6, Hzhnv6, Ozhnv6, Vzhnv6, C0inv6, J0inv6, Q0inv6;
wire X0inv6, E1inv6, L1inv6, S1inv6, Z1inv6, G2inv6, N2inv6, U2inv6, B3inv6, I3inv6;
wire P3inv6, W3inv6, D4inv6, K4inv6, R4inv6, Y4inv6, F5inv6, M5inv6, T5inv6, A6inv6;
wire H6inv6, O6inv6, V6inv6, C7inv6, J7inv6, Q7inv6, X7inv6, E8inv6, L8inv6, S8inv6;
wire Z8inv6, G9inv6, N9inv6, U9inv6, Bainv6, Iainv6, Painv6, Wainv6, Dbinv6, Kbinv6;
wire Rbinv6, Ybinv6, Fcinv6, Mcinv6, Tcinv6, Adinv6, Hdinv6, Odinv6, Vdinv6, Ceinv6;
wire Jeinv6, Qeinv6, Xeinv6, Efinv6, Lfinv6, Sfinv6, Zfinv6, Gginv6, Nginv6, Uginv6;
wire Bhinv6, Ihinv6, Phinv6, Whinv6, Diinv6, Kiinv6, Riinv6, Yiinv6, Fjinv6, Mjinv6;
wire Tjinv6, Akinv6, Hkinv6, Okinv6, Vkinv6, Clinv6, Jlinv6, Qlinv6, Xlinv6, Eminv6;
wire Lminv6, Sminv6, Zminv6, Gninv6, Nninv6, Uninv6, Boinv6, Ioinv6, Poinv6, Woinv6;
wire Dpinv6, Kpinv6, Rpinv6, Ypinv6, Fqinv6, Mqinv6, Tqinv6, Arinv6, Hrinv6, Orinv6;
wire Vrinv6, Csinv6, Jsinv6, Qsinv6, Xsinv6, Etinv6, Ltinv6, Stinv6, Ztinv6, Guinv6;
wire Nuinv6, Uuinv6, Bvinv6, Ivinv6, Pvinv6, Wvinv6, Dwinv6, Kwinv6, Rwinv6, Ywinv6;
wire Fxinv6, Mxinv6, Txinv6, Ayinv6, Hyinv6, Oyinv6, Vyinv6, Czinv6, Jzinv6, Qzinv6;
wire Xzinv6, E0jnv6, L0jnv6, S0jnv6, Z0jnv6, G1jnv6, N1jnv6, U1jnv6, B2jnv6, I2jnv6;
wire P2jnv6, W2jnv6, D3jnv6, K3jnv6, R3jnv6, Y3jnv6, F4jnv6, M4jnv6, T4jnv6, A5jnv6;
wire H5jnv6, O5jnv6, V5jnv6, C6jnv6, J6jnv6, Q6jnv6, X6jnv6, E7jnv6, L7jnv6, S7jnv6;
wire Z7jnv6, G8jnv6, N8jnv6, U8jnv6, B9jnv6, I9jnv6, P9jnv6, W9jnv6, Dajnv6, Kajnv6;
wire Rajnv6, Yajnv6, Fbjnv6, Mbjnv6, Tbjnv6, Acjnv6, Hcjnv6, Ocjnv6, Vcjnv6, Cdjnv6;
wire Jdjnv6, Qdjnv6, Xdjnv6, Eejnv6, Lejnv6, Sejnv6, Zejnv6, Gfjnv6, Nfjnv6, Ufjnv6;
wire Bgjnv6, Igjnv6, Pgjnv6, Wgjnv6, Dhjnv6, Khjnv6, Rhjnv6, Yhjnv6, Fijnv6, Mijnv6;
wire Tijnv6, Ajjnv6, Hjjnv6, Ojjnv6, Vjjnv6, Ckjnv6, Jkjnv6, Qkjnv6, Xkjnv6, Eljnv6;
wire Lljnv6, Sljnv6, Zljnv6, Gmjnv6, Nmjnv6, Umjnv6, Bnjnv6, Injnv6, Pnjnv6, Wnjnv6;
wire Dojnv6, Kojnv6, Rojnv6, Yojnv6, Fpjnv6, Mpjnv6, Tpjnv6, Aqjnv6, Hqjnv6, Oqjnv6;
wire Vqjnv6, Crjnv6, Jrjnv6, Qrjnv6, Xrjnv6, Esjnv6, Lsjnv6, Ssjnv6, Zsjnv6, Gtjnv6;
wire Ntjnv6, Utjnv6, Bujnv6, Iujnv6, Pujnv6, Wujnv6, Dvjnv6, Kvjnv6, Rvjnv6, Yvjnv6;
wire Fwjnv6, Mwjnv6, Twjnv6, Axjnv6, Hxjnv6, Oxjnv6, Vxjnv6, Cyjnv6, Jyjnv6, Qyjnv6;
wire Xyjnv6, Ezjnv6, Lzjnv6, Szjnv6, Zzjnv6, G0knv6, N0knv6, U0knv6, B1knv6, I1knv6;
wire P1knv6, W1knv6, D2knv6, K2knv6, R2knv6, Y2knv6, F3knv6, M3knv6, T3knv6, A4knv6;
wire H4knv6, O4knv6, V4knv6, C5knv6, J5knv6, Q5knv6, X5knv6, E6knv6, L6knv6, S6knv6;
wire Z6knv6, G7knv6, N7knv6, U7knv6, B8knv6, I8knv6, P8knv6, W8knv6, D9knv6, K9knv6;
wire R9knv6, Y9knv6, Faknv6, Maknv6, Taknv6, Abknv6, Hbknv6, Obknv6, Vbknv6, Ccknv6;
wire Jcknv6, Qcknv6, Xcknv6, Edknv6, Ldknv6, Sdknv6, Zdknv6, Geknv6, Neknv6, Ueknv6;
wire Bfknv6, Ifknv6, Pfknv6, Wfknv6, Dgknv6, Kgknv6, Rgknv6, Ygknv6, Fhknv6, Mhknv6;
wire Thknv6, Aiknv6, Hiknv6, Oiknv6, Viknv6, Cjknv6, Jjknv6, Qjknv6, Xjknv6, Ekknv6;
wire Lkknv6, Skknv6, Zkknv6, Glknv6, Nlknv6, Ulknv6, Bmknv6, Imknv6, Pmknv6, Wmknv6;
wire Dnknv6, Knknv6, Rnknv6, Ynknv6, Foknv6, Moknv6, Toknv6, Apknv6, Hpknv6, Opknv6;
wire Vpknv6, Cqknv6, Jqknv6, Qqknv6, Xqknv6, Erknv6, Lrknv6, Srknv6, Zrknv6, Gsknv6;
wire Nsknv6, Usknv6, Btknv6, Itknv6, Ptknv6, Wtknv6, Duknv6, Kuknv6, Ruknv6, Yuknv6;
wire Fvknv6, Mvknv6, Tvknv6, Awknv6, Hwknv6, Owknv6, Vwknv6, Cxknv6, Jxknv6, Qxknv6;
wire Xxknv6, Eyknv6, Lyknv6, Syknv6, Zyknv6, Gzknv6, Nzknv6, Uzknv6, B0lnv6, I0lnv6;
wire P0lnv6, W0lnv6, D1lnv6, K1lnv6, R1lnv6, Y1lnv6, F2lnv6, M2lnv6, T2lnv6, A3lnv6;
wire H3lnv6, O3lnv6, V3lnv6, C4lnv6, J4lnv6, Q4lnv6, X4lnv6, E5lnv6, L5lnv6, S5lnv6;
wire Z5lnv6, G6lnv6, N6lnv6, U6lnv6, B7lnv6, I7lnv6, P7lnv6, W7lnv6, D8lnv6, K8lnv6;
wire R8lnv6, Y8lnv6, F9lnv6, M9lnv6, T9lnv6, Aalnv6, Halnv6, Oalnv6, Valnv6, Cblnv6;
wire Jblnv6, Qblnv6, Xblnv6, Eclnv6, Lclnv6, Sclnv6, Zclnv6, Gdlnv6, Ndlnv6, Udlnv6;
wire Belnv6, Ielnv6, Pelnv6, Welnv6, Dflnv6, Kflnv6, Rflnv6, Yflnv6, Fglnv6, Mglnv6;
wire Tglnv6, Ahlnv6, Hhlnv6, Ohlnv6, Vhlnv6, Cilnv6, Jilnv6, Qilnv6, Xilnv6, Ejlnv6;
wire Ljlnv6, Sjlnv6, Zjlnv6, Gklnv6, Nklnv6, Uklnv6, Bllnv6, Illnv6, Pllnv6, Wllnv6;
wire Dmlnv6, Kmlnv6, Rmlnv6, Ymlnv6, Fnlnv6, Mnlnv6, Tnlnv6, Aolnv6, Holnv6, Oolnv6;
wire Volnv6, Cplnv6, Jplnv6, Qplnv6, Xplnv6, Eqlnv6, Lqlnv6, Sqlnv6, Zqlnv6, Grlnv6;
wire Nrlnv6, Urlnv6, Bslnv6, Islnv6, Pslnv6, Wslnv6, Dtlnv6, Ktlnv6, Rtlnv6, Ytlnv6;
wire Fulnv6, Mulnv6, Tulnv6, Avlnv6, Hvlnv6, Ovlnv6, Vvlnv6, Cwlnv6, Jwlnv6, Qwlnv6;
wire Xwlnv6, Exlnv6, Lxlnv6, Sxlnv6, Zxlnv6, Gylnv6, Nylnv6, Uylnv6, Bzlnv6, Izlnv6;
wire Pzlnv6, Wzlnv6, D0mnv6, K0mnv6, R0mnv6, Y0mnv6, F1mnv6, M1mnv6, T1mnv6, A2mnv6;
wire H2mnv6, O2mnv6, V2mnv6, C3mnv6, J3mnv6, Q3mnv6, X3mnv6, E4mnv6, L4mnv6, S4mnv6;
wire Z4mnv6, G5mnv6, N5mnv6, U5mnv6, B6mnv6, I6mnv6, P6mnv6, W6mnv6, D7mnv6, K7mnv6;
wire R7mnv6, Y7mnv6, F8mnv6, M8mnv6, T8mnv6, A9mnv6, H9mnv6, O9mnv6, V9mnv6, Camnv6;
wire Jamnv6, Qamnv6, Xamnv6, Ebmnv6, Lbmnv6, Sbmnv6, Zbmnv6, Gcmnv6, Ncmnv6, Ucmnv6;
wire Bdmnv6, Idmnv6, Pdmnv6, Wdmnv6, Demnv6, Kemnv6, Remnv6, Yemnv6, Ffmnv6, Mfmnv6;
wire Tfmnv6, Agmnv6, Hgmnv6, Ogmnv6, Vgmnv6, Chmnv6, Jhmnv6, Qhmnv6, Xhmnv6, Eimnv6;
wire Limnv6, Simnv6, Zimnv6, Gjmnv6, Njmnv6, Ujmnv6, Bkmnv6, Ikmnv6, Pkmnv6, Wkmnv6;
wire Dlmnv6, Klmnv6, Rlmnv6, Ylmnv6, Fmmnv6, Mmmnv6, Tmmnv6, Anmnv6, Hnmnv6, Onmnv6;
wire Vnmnv6, Comnv6, Jomnv6, Qomnv6, Xomnv6, Epmnv6, Lpmnv6, Spmnv6, Zpmnv6, Gqmnv6;
wire Nqmnv6, Uqmnv6, Brmnv6, Irmnv6, Prmnv6, Wrmnv6, Dsmnv6, Ksmnv6, Rsmnv6, Ysmnv6;
wire Ftmnv6, Mtmnv6, Ttmnv6, Aumnv6, Humnv6, Oumnv6, Vumnv6, Cvmnv6, Jvmnv6, Qvmnv6;
wire Xvmnv6, Ewmnv6, Lwmnv6, Swmnv6, Zwmnv6, Gxmnv6, Nxmnv6, Uxmnv6, Bymnv6, Iymnv6;
wire Pymnv6, Wymnv6, Dzmnv6, Kzmnv6, Rzmnv6, Yzmnv6, F0nnv6, M0nnv6, T0nnv6, A1nnv6;
wire H1nnv6, O1nnv6, V1nnv6, C2nnv6, J2nnv6, Q2nnv6, X2nnv6, E3nnv6, L3nnv6, S3nnv6;
wire Z3nnv6, G4nnv6, N4nnv6, U4nnv6, B5nnv6, I5nnv6, P5nnv6, W5nnv6, D6nnv6, K6nnv6;
wire R6nnv6, Y6nnv6, F7nnv6, M7nnv6, T7nnv6, A8nnv6, H8nnv6, O8nnv6, V8nnv6, C9nnv6;
wire J9nnv6, Q9nnv6, X9nnv6, Eannv6, Lannv6, Sannv6, Zannv6, Gbnnv6, Nbnnv6, Ubnnv6;
wire Bcnnv6, Icnnv6, Pcnnv6, Wcnnv6, Ddnnv6, Kdnnv6, Rdnnv6, Ydnnv6, Fennv6, Mennv6;
wire Tennv6, Afnnv6, Hfnnv6, Ofnnv6, Vfnnv6, Cgnnv6, Jgnnv6, Qgnnv6, Xgnnv6, Ehnnv6;
wire Lhnnv6, Shnnv6, Zhnnv6, Ginnv6, Ninnv6, Uinnv6, Bjnnv6, Ijnnv6, Pjnnv6, Wjnnv6;
wire Dknnv6, Kknnv6, Rknnv6, Yknnv6, Flnnv6, Mlnnv6, Tlnnv6, Amnnv6, Hmnnv6, Omnnv6;
wire Vmnnv6, Cnnnv6, Jnnnv6, Qnnnv6, Xnnnv6, Eonnv6, Lonnv6, Sonnv6, Zonnv6, Gpnnv6;
wire Npnnv6, Upnnv6, Bqnnv6, Iqnnv6, Pqnnv6, Wqnnv6, Drnnv6, Krnnv6, Rrnnv6, Yrnnv6;
wire Fsnnv6, Msnnv6, Tsnnv6, Atnnv6, Htnnv6, Otnnv6, Vtnnv6, Cunnv6, Junnv6, Qunnv6;
wire Xunnv6, Evnnv6, Lvnnv6, Svnnv6, Zvnnv6, Gwnnv6, Nwnnv6, Uwnnv6, Bxnnv6, Ixnnv6;
wire Pxnnv6, Wxnnv6, Dynnv6, Kynnv6, Rynnv6, Yynnv6, Fznnv6, Mznnv6, Tznnv6, A0onv6;
wire H0onv6, O0onv6, V0onv6, C1onv6, J1onv6, Q1onv6, X1onv6, E2onv6, L2onv6, S2onv6;
wire Z2onv6, G3onv6, N3onv6, U3onv6, B4onv6, I4onv6, P4onv6, W4onv6, D5onv6, K5onv6;
wire R5onv6, Y5onv6, F6onv6, M6onv6, T6onv6, A7onv6, H7onv6, O7onv6, V7onv6, C8onv6;
wire J8onv6, Q8onv6, X8onv6, E9onv6, L9onv6, S9onv6, Z9onv6, Gaonv6, Naonv6, Uaonv6;
wire Bbonv6, Ibonv6, Pbonv6, Wbonv6, Dconv6, Kconv6, Rconv6, Yconv6, Fdonv6, Mdonv6;
wire Tdonv6, Aeonv6, Heonv6, Oeonv6, Veonv6, Cfonv6, Jfonv6, Qfonv6, Xfonv6, Egonv6;
wire Lgonv6, Sgonv6, Zgonv6, Ghonv6, Nhonv6, Uhonv6, Bionv6, Iionv6, Pionv6, Wionv6;
wire Djonv6, Kjonv6, Rjonv6, Yjonv6, Fkonv6, Mkonv6, Tkonv6, Alonv6, Hlonv6, Olonv6;
wire Vlonv6, Cmonv6, Jmonv6, Qmonv6, Xmonv6, Enonv6, Lnonv6, Snonv6, Znonv6, Goonv6;
wire Noonv6, Uoonv6, Bponv6, Iponv6, Pponv6, Wponv6, Dqonv6, Kqonv6, Rqonv6, Yqonv6;
wire Fronv6, Mronv6, Tronv6, Asonv6, Hsonv6, Osonv6, Vsonv6, Ctonv6, Jtonv6, Qtonv6;
wire Xtonv6, Euonv6, Luonv6, Suonv6, Zuonv6, Gvonv6, Nvonv6, Uvonv6, Bwonv6, Iwonv6;
wire Pwonv6, Wwonv6, Dxonv6, Kxonv6, Rxonv6, Yxonv6, Fyonv6, Myonv6, Tyonv6, Azonv6;
wire Hzonv6, Ozonv6, Vzonv6, C0pnv6, J0pnv6, Q0pnv6, X0pnv6, E1pnv6, L1pnv6, S1pnv6;
wire Z1pnv6, G2pnv6, N2pnv6, U2pnv6, B3pnv6, I3pnv6, P3pnv6, W3pnv6, D4pnv6, K4pnv6;
wire R4pnv6, Y4pnv6, F5pnv6, M5pnv6, T5pnv6, A6pnv6, H6pnv6, O6pnv6, V6pnv6, C7pnv6;
wire J7pnv6, Q7pnv6, X7pnv6, E8pnv6, L8pnv6, S8pnv6, Z8pnv6, G9pnv6, N9pnv6, U9pnv6;
wire Bapnv6, Iapnv6, Papnv6, Wapnv6, Dbpnv6, Kbpnv6, Rbpnv6, Ybpnv6, Fcpnv6, Mcpnv6;
wire Tcpnv6, Adpnv6, Hdpnv6, Odpnv6, Vdpnv6, Cepnv6, Jepnv6, Qepnv6, Xepnv6, Efpnv6;
wire Lfpnv6, Sfpnv6, Zfpnv6, Ggpnv6, Ngpnv6, Ugpnv6, Bhpnv6, Ihpnv6, Phpnv6, Whpnv6;
wire Dipnv6, Kipnv6, Ripnv6, Yipnv6, Fjpnv6, Mjpnv6, Tjpnv6, Akpnv6, Hkpnv6, Okpnv6;
wire Vkpnv6, Clpnv6, Jlpnv6, Qlpnv6, Xlpnv6, Empnv6, Lmpnv6, Smpnv6, Zmpnv6, Gnpnv6;
wire Nnpnv6, Unpnv6, Bopnv6, Iopnv6, Popnv6, Wopnv6, Dppnv6, Kppnv6, Rppnv6, Yppnv6;
wire Fqpnv6, Mqpnv6, Tqpnv6, Arpnv6, Hrpnv6, Orpnv6, Vrpnv6, Cspnv6, Jspnv6, Qspnv6;
wire Xspnv6, Etpnv6, Ltpnv6, Stpnv6, Ztpnv6, Gupnv6, Nupnv6, Uupnv6, Bvpnv6, Ivpnv6;
wire Pvpnv6, Wvpnv6, Dwpnv6, Kwpnv6, Rwpnv6, Ywpnv6, Fxpnv6, Mxpnv6, Txpnv6, Aypnv6;
wire Hypnv6, Oypnv6, Vypnv6, Czpnv6, Jzpnv6, Qzpnv6, Xzpnv6, E0qnv6, L0qnv6, S0qnv6;
wire Z0qnv6, G1qnv6, N1qnv6, U1qnv6, B2qnv6, I2qnv6, P2qnv6, W2qnv6, D3qnv6, K3qnv6;
wire R3qnv6, Y3qnv6, F4qnv6, M4qnv6, T4qnv6, A5qnv6, H5qnv6, O5qnv6, V5qnv6, C6qnv6;
wire J6qnv6, Q6qnv6, X6qnv6, E7qnv6, L7qnv6, S7qnv6, Z7qnv6, G8qnv6, N8qnv6, U8qnv6;
wire B9qnv6, I9qnv6, P9qnv6, W9qnv6, Daqnv6, Kaqnv6, Raqnv6, Yaqnv6, Fbqnv6, Mbqnv6;
wire Tbqnv6, Acqnv6, Hcqnv6, Ocqnv6, Vcqnv6, Cdqnv6, Jdqnv6, Qdqnv6, Xdqnv6, Eeqnv6;
wire Leqnv6, Seqnv6, Zeqnv6, Gfqnv6, Nfqnv6, Ufqnv6, Bgqnv6, Igqnv6, Pgqnv6, Wgqnv6;
wire Dhqnv6, Khqnv6, Rhqnv6, Yhqnv6, Fiqnv6, Miqnv6, Tiqnv6, Ajqnv6, Hjqnv6, Ojqnv6;
wire Vjqnv6, Ckqnv6, Jkqnv6, Qkqnv6, Xkqnv6, Elqnv6, Llqnv6, Slqnv6, Zlqnv6, Gmqnv6;
wire Nmqnv6, Umqnv6, Bnqnv6, Inqnv6, Pnqnv6, Wnqnv6, Doqnv6, Koqnv6, Roqnv6, Yoqnv6;
wire Fpqnv6, Mpqnv6, Tpqnv6, Aqqnv6, Hqqnv6, Oqqnv6, Vqqnv6, Crqnv6, Jrqnv6, Qrqnv6;
wire Xrqnv6, Esqnv6, Lsqnv6, Ssqnv6, Zsqnv6, Gtqnv6, Ntqnv6, Utqnv6, Buqnv6, Iuqnv6;
wire Puqnv6, Wuqnv6, Dvqnv6, Kvqnv6, Rvqnv6, Yvqnv6, Fwqnv6, Mwqnv6, Twqnv6, Axqnv6;
wire Hxqnv6, Oxqnv6, Vxqnv6, Cyqnv6, Jyqnv6, Qyqnv6, Xyqnv6, Ezqnv6, Lzqnv6, Szqnv6;
wire Zzqnv6, G0rnv6, N0rnv6, U0rnv6, B1rnv6, I1rnv6, P1rnv6, W1rnv6, D2rnv6, K2rnv6;
wire R2rnv6, Y2rnv6, F3rnv6, M3rnv6, T3rnv6, A4rnv6, H4rnv6, O4rnv6, V4rnv6, C5rnv6;
wire J5rnv6, Q5rnv6, X5rnv6, E6rnv6, L6rnv6, S6rnv6, Z6rnv6, G7rnv6, N7rnv6, U7rnv6;
wire B8rnv6, I8rnv6, P8rnv6, W8rnv6, D9rnv6, K9rnv6, R9rnv6, Y9rnv6, Farnv6, Marnv6;
wire Tarnv6, Abrnv6, Hbrnv6, Obrnv6, Vbrnv6, Ccrnv6, Jcrnv6, Qcrnv6, Xcrnv6, Edrnv6;
wire Ldrnv6, Sdrnv6, Zdrnv6, Gernv6, Nernv6, Uernv6, Bfrnv6, Ifrnv6, Pfrnv6, Wfrnv6;
wire Dgrnv6, Kgrnv6, Rgrnv6, Ygrnv6, Fhrnv6, Mhrnv6, Thrnv6, Airnv6, Hirnv6, Oirnv6;
wire Virnv6, Cjrnv6, Jjrnv6, Qjrnv6, Xjrnv6, Ekrnv6, Lkrnv6, Skrnv6, Zkrnv6, Glrnv6;
wire Nlrnv6, Ulrnv6, Bmrnv6, Imrnv6, Pmrnv6, Wmrnv6, Dnrnv6, Knrnv6, Rnrnv6, Ynrnv6;
wire Fornv6, Mornv6, Tornv6, Aprnv6, Hprnv6, Oprnv6, Vprnv6, Cqrnv6, Jqrnv6, Qqrnv6;
wire Xqrnv6, Errnv6, Lrrnv6, Srrnv6, Zrrnv6, Gsrnv6, Nsrnv6, Usrnv6, Btrnv6, Itrnv6;
wire Ptrnv6, Wtrnv6, Durnv6, Kurnv6, Rurnv6, Yurnv6, Fvrnv6, Mvrnv6, Tvrnv6, Awrnv6;
wire Hwrnv6, Owrnv6, Vwrnv6, Cxrnv6, Jxrnv6, Qxrnv6, Xxrnv6, Eyrnv6, Lyrnv6, Syrnv6;
wire Zyrnv6, Gzrnv6, Nzrnv6, Uzrnv6, B0snv6, I0snv6, P0snv6, W0snv6, D1snv6, K1snv6;
wire R1snv6, Y1snv6, F2snv6, M2snv6, T2snv6, A3snv6, H3snv6, O3snv6, V3snv6, C4snv6;
wire J4snv6, Q4snv6, X4snv6, E5snv6, L5snv6, S5snv6, Z5snv6, G6snv6, N6snv6, U6snv6;
wire B7snv6, I7snv6, P7snv6, W7snv6, D8snv6, K8snv6, R8snv6, Y8snv6, F9snv6, M9snv6;
wire T9snv6, Aasnv6, Hasnv6, Oasnv6, Vasnv6, Cbsnv6, Jbsnv6, Qbsnv6, Xbsnv6, Ecsnv6;
wire Lcsnv6, Scsnv6, Zcsnv6, Gdsnv6, Ndsnv6, Udsnv6, Besnv6, Iesnv6, Pesnv6, Wesnv6;
wire Dfsnv6, Kfsnv6, Rfsnv6, Yfsnv6, Fgsnv6, Mgsnv6, Tgsnv6, Ahsnv6, Hhsnv6, Ohsnv6;
wire Vhsnv6, Cisnv6, Jisnv6, Qisnv6, Xisnv6, Ejsnv6, Ljsnv6, Sjsnv6, Zjsnv6, Gksnv6;
wire Nksnv6, Uksnv6, Blsnv6, Ilsnv6, Plsnv6, Wlsnv6, Dmsnv6, Kmsnv6, Rmsnv6, Ymsnv6;
wire Fnsnv6, Mnsnv6, Tnsnv6, Aosnv6, Hosnv6, Oosnv6, Vosnv6, Cpsnv6, Jpsnv6, Qpsnv6;
wire Xpsnv6, Eqsnv6, Lqsnv6, Sqsnv6, Zqsnv6, Grsnv6, Nrsnv6, Ursnv6, Bssnv6, Issnv6;
wire Pssnv6, Wssnv6, Dtsnv6, Ktsnv6, Rtsnv6, Ytsnv6, Fusnv6, Musnv6, Tusnv6, Avsnv6;
wire Hvsnv6, Ovsnv6, Vvsnv6, Cwsnv6, Jwsnv6, Qwsnv6, Xwsnv6, Exsnv6, Lxsnv6, Sxsnv6;
wire Zxsnv6, Gysnv6, Nysnv6, Uysnv6, Bzsnv6, Izsnv6, Pzsnv6, Wzsnv6, D0tnv6, K0tnv6;
wire R0tnv6, Y0tnv6, F1tnv6, M1tnv6, T1tnv6, A2tnv6, H2tnv6, O2tnv6, V2tnv6, C3tnv6;
wire J3tnv6, Q3tnv6, X3tnv6, E4tnv6, L4tnv6, S4tnv6, Z4tnv6, G5tnv6, N5tnv6, U5tnv6;
wire B6tnv6, I6tnv6, P6tnv6, W6tnv6, D7tnv6, K7tnv6, R7tnv6, Y7tnv6, F8tnv6, M8tnv6;
wire T8tnv6, A9tnv6, H9tnv6, O9tnv6, V9tnv6, Catnv6, Jatnv6, Qatnv6, Xatnv6, Ebtnv6;
wire Lbtnv6, Sbtnv6, Zbtnv6, Gctnv6, Nctnv6, Uctnv6, Bdtnv6, Idtnv6, Pdtnv6, Wdtnv6;
wire Detnv6, Ketnv6, Retnv6, Yetnv6, Fftnv6, Mftnv6, Tftnv6, Agtnv6, Hgtnv6, Ogtnv6;
wire Vgtnv6, Chtnv6, Jhtnv6, Qhtnv6, Xhtnv6, Eitnv6, Litnv6, Sitnv6, Zitnv6, Gjtnv6;
wire Njtnv6, Ujtnv6, Bktnv6, Iktnv6, Pktnv6, Wktnv6, Dltnv6, Kltnv6, Rltnv6, Yltnv6;
wire Fmtnv6, Mmtnv6, Tmtnv6, Antnv6, Hntnv6, Ontnv6, Vntnv6, Cotnv6, Jotnv6, Qotnv6;
wire Xotnv6, Eptnv6, Lptnv6, Sptnv6, Zptnv6, Gqtnv6, Nqtnv6, Uqtnv6, Brtnv6, Irtnv6;
wire Prtnv6, Wrtnv6, Dstnv6, Kstnv6, Rstnv6, Ystnv6, Fttnv6, Mttnv6, Tttnv6, Autnv6;
wire Hutnv6, Outnv6, Vutnv6, Cvtnv6, Jvtnv6, Qvtnv6, Xvtnv6, Ewtnv6, Lwtnv6, Swtnv6;
wire Zwtnv6, Gxtnv6, Nxtnv6, Uxtnv6, Bytnv6, Iytnv6, Pytnv6, Wytnv6, Dztnv6, Kztnv6;
wire Rztnv6, Yztnv6, F0unv6, M0unv6, T0unv6, A1unv6, H1unv6, O1unv6, V1unv6, C2unv6;
wire J2unv6, Q2unv6, X2unv6, E3unv6, L3unv6, S3unv6, Z3unv6, G4unv6, N4unv6, U4unv6;
wire B5unv6, I5unv6, P5unv6, W5unv6, D6unv6, K6unv6, R6unv6, Y6unv6, F7unv6, M7unv6;
wire T7unv6, A8unv6, H8unv6, O8unv6, V8unv6, C9unv6, J9unv6, Q9unv6, X9unv6, Eaunv6;
wire Launv6, Saunv6, Zaunv6, Gbunv6, Nbunv6, Ubunv6, Bcunv6, Icunv6, Pcunv6, Wcunv6;
wire Ddunv6, Kdunv6, Rdunv6, Ydunv6, Feunv6, Meunv6, Teunv6, Afunv6, Hfunv6, Ofunv6;
wire Vfunv6, Cgunv6, Jgunv6, Qgunv6, Xgunv6, Ehunv6, Lhunv6, Shunv6, Zhunv6, Giunv6;
wire Niunv6, Uiunv6, Bjunv6, Ijunv6, Pjunv6, Wjunv6, Dkunv6, Kkunv6, Rkunv6, Ykunv6;
wire Flunv6, Mlunv6, Tlunv6, Amunv6, Hmunv6, Omunv6, Vmunv6, Cnunv6, Jnunv6, Qnunv6;
wire Xnunv6, Eounv6, Lounv6, Sounv6, Zounv6, Gpunv6, Npunv6, Upunv6, Bqunv6, Iqunv6;
wire Pqunv6, Wqunv6, Drunv6, Krunv6, Rrunv6, Yrunv6, Fsunv6, Msunv6, Tsunv6, Atunv6;
wire Htunv6, Otunv6, Vtunv6, Cuunv6, Juunv6, Quunv6, Xuunv6, Evunv6, Lvunv6, Svunv6;
wire Zvunv6, Gwunv6, Nwunv6, Uwunv6, Bxunv6, Ixunv6, Pxunv6, Wxunv6, Dyunv6, Kyunv6;
wire Ryunv6, Yyunv6, Fzunv6, Mzunv6, Tzunv6, A0vnv6, H0vnv6, O0vnv6, V0vnv6, C1vnv6;
wire J1vnv6, Q1vnv6, X1vnv6, E2vnv6, L2vnv6, S2vnv6, Z2vnv6, G3vnv6, N3vnv6, U3vnv6;
wire B4vnv6, I4vnv6, P4vnv6, W4vnv6, D5vnv6, K5vnv6, R5vnv6, Y5vnv6, F6vnv6, M6vnv6;
wire T6vnv6, A7vnv6, H7vnv6, O7vnv6, V7vnv6, C8vnv6, J8vnv6, Q8vnv6, X8vnv6, E9vnv6;
wire L9vnv6, S9vnv6, Z9vnv6, Gavnv6, Navnv6, Uavnv6, Bbvnv6, Ibvnv6, Pbvnv6, Wbvnv6;
wire Dcvnv6, Kcvnv6, Rcvnv6, Ycvnv6, Fdvnv6, Mdvnv6, Tdvnv6, Aevnv6, Hevnv6, Oevnv6;
wire Vevnv6, Cfvnv6, Jfvnv6, Qfvnv6, Xfvnv6, Egvnv6, Lgvnv6, Sgvnv6, Zgvnv6, Ghvnv6;
wire Nhvnv6, Uhvnv6, Bivnv6, Iivnv6, Pivnv6, Wivnv6, Djvnv6, Kjvnv6, Rjvnv6, Yjvnv6;
wire Fkvnv6, Mkvnv6, Tkvnv6, Alvnv6, Hlvnv6, Olvnv6, Vlvnv6, Cmvnv6, Jmvnv6, Qmvnv6;
wire Xmvnv6, Envnv6, Lnvnv6, Snvnv6, Znvnv6, Govnv6, Novnv6, Uovnv6, Bpvnv6, Ipvnv6;
wire Ppvnv6, Wpvnv6, Dqvnv6, Kqvnv6, Rqvnv6, Yqvnv6, Frvnv6, Mrvnv6, Trvnv6, Asvnv6;
wire Hsvnv6, Osvnv6, Vsvnv6, Ctvnv6, Jtvnv6, Qtvnv6, Xtvnv6, Euvnv6, Luvnv6, Suvnv6;
wire Zuvnv6, Gvvnv6, Nvvnv6, Uvvnv6, Bwvnv6, Iwvnv6, Pwvnv6, Wwvnv6, Dxvnv6, Kxvnv6;
wire Rxvnv6, Yxvnv6, Fyvnv6, Myvnv6, Tyvnv6, Azvnv6, Hzvnv6, Ozvnv6, Vzvnv6, C0wnv6;
wire J0wnv6, Q0wnv6, X0wnv6, E1wnv6, L1wnv6, S1wnv6, Z1wnv6, G2wnv6, N2wnv6, U2wnv6;
wire B3wnv6, I3wnv6, P3wnv6, W3wnv6, D4wnv6, K4wnv6, R4wnv6, Y4wnv6, F5wnv6, M5wnv6;
wire T5wnv6, A6wnv6, H6wnv6, O6wnv6, V6wnv6, C7wnv6, J7wnv6, Q7wnv6, X7wnv6, E8wnv6;
wire L8wnv6, S8wnv6, Z8wnv6, G9wnv6, N9wnv6, U9wnv6, Bawnv6, Iawnv6, Pawnv6, Wawnv6;
wire Dbwnv6, Kbwnv6, Rbwnv6, Ybwnv6, Fcwnv6, Mcwnv6, Tcwnv6, Adwnv6, Hdwnv6, Odwnv6;
wire Vdwnv6, Cewnv6, Jewnv6, Qewnv6, Xewnv6, Efwnv6, Lfwnv6, Sfwnv6, Zfwnv6, Ggwnv6;
wire Ngwnv6, Ugwnv6, Bhwnv6, Ihwnv6, Phwnv6, Whwnv6, Diwnv6, Kiwnv6, Riwnv6, Yiwnv6;
wire Fjwnv6, Mjwnv6, Tjwnv6, Akwnv6, Hkwnv6, Okwnv6, Vkwnv6, Clwnv6, Jlwnv6, Qlwnv6;
wire Xlwnv6, Emwnv6, Lmwnv6, Smwnv6, Zmwnv6, Gnwnv6, Nnwnv6, Unwnv6, Bownv6, Iownv6;
wire Pownv6, Wownv6, Dpwnv6, Kpwnv6, Rpwnv6, Ypwnv6, Fqwnv6, Mqwnv6, Tqwnv6, Arwnv6;
wire Hrwnv6, Orwnv6, Vrwnv6, Cswnv6, Jswnv6, Qswnv6, Xswnv6, Etwnv6, Ltwnv6, Stwnv6;
wire Ztwnv6, Guwnv6, Nuwnv6, Uuwnv6, Bvwnv6, Ivwnv6, Pvwnv6, Wvwnv6, Dwwnv6, Kwwnv6;
wire Rwwnv6, Ywwnv6, Fxwnv6, Mxwnv6, Txwnv6, Aywnv6, Hywnv6, Oywnv6, Vywnv6, Czwnv6;
wire Jzwnv6, Qzwnv6, Xzwnv6, E0xnv6, L0xnv6, S0xnv6, Z0xnv6, G1xnv6, N1xnv6, U1xnv6;
wire B2xnv6, I2xnv6, P2xnv6, W2xnv6, D3xnv6, K3xnv6, R3xnv6, Y3xnv6, F4xnv6, M4xnv6;
wire T4xnv6, A5xnv6, H5xnv6, O5xnv6, V5xnv6, C6xnv6, J6xnv6, Q6xnv6, X6xnv6, E7xnv6;
wire L7xnv6, S7xnv6, Z7xnv6, G8xnv6, N8xnv6, U8xnv6, B9xnv6, I9xnv6, P9xnv6, W9xnv6;
wire Daxnv6, Kaxnv6, Raxnv6, Yaxnv6, Fbxnv6, Mbxnv6, Tbxnv6, Acxnv6, Hcxnv6, Ocxnv6;
wire Vcxnv6, Cdxnv6, Jdxnv6, Qdxnv6, Xdxnv6, Eexnv6, Lexnv6, Sexnv6, Zexnv6, Gfxnv6;
wire Nfxnv6, Ufxnv6, Bgxnv6, Igxnv6, Pgxnv6, Wgxnv6, Dhxnv6, Khxnv6, Rhxnv6, Yhxnv6;
wire Fixnv6, Mixnv6, Tixnv6, Ajxnv6, Hjxnv6, Ojxnv6, Vjxnv6, Ckxnv6, Jkxnv6, Qkxnv6;
wire Xkxnv6, Elxnv6, Llxnv6, Slxnv6, Zlxnv6, Gmxnv6, Nmxnv6, Umxnv6, Bnxnv6, Inxnv6;
wire Pnxnv6, Wnxnv6, Doxnv6, Koxnv6, Roxnv6, Yoxnv6, Fpxnv6, Mpxnv6, Tpxnv6, Aqxnv6;
wire Hqxnv6, Oqxnv6, Vqxnv6, Crxnv6, Jrxnv6, Qrxnv6, Xrxnv6, Esxnv6, Lsxnv6, Ssxnv6;
wire Zsxnv6, Gtxnv6, Ntxnv6, Utxnv6, Buxnv6, Iuxnv6, Puxnv6, Wuxnv6, Dvxnv6, Kvxnv6;
wire Rvxnv6, Yvxnv6, Fwxnv6, Mwxnv6, Twxnv6, Axxnv6, Hxxnv6, Oxxnv6, Vxxnv6, Cyxnv6;
wire Jyxnv6, Qyxnv6, Xyxnv6, Ezxnv6, Lzxnv6, Szxnv6, Zzxnv6, G0ynv6, N0ynv6, U0ynv6;
wire B1ynv6, I1ynv6, P1ynv6, W1ynv6, D2ynv6, K2ynv6, R2ynv6, Y2ynv6, F3ynv6, M3ynv6;
wire T3ynv6, A4ynv6, H4ynv6, O4ynv6, V4ynv6, C5ynv6, J5ynv6, Q5ynv6, X5ynv6, E6ynv6;
wire L6ynv6, S6ynv6, Z6ynv6, G7ynv6, N7ynv6, U7ynv6, B8ynv6, I8ynv6, P8ynv6, W8ynv6;
wire D9ynv6, K9ynv6, R9ynv6, Y9ynv6, Faynv6, Maynv6, Taynv6, Abynv6, Hbynv6, Obynv6;
wire Vbynv6, Ccynv6, Jcynv6, Qcynv6, Xcynv6, Edynv6, Ldynv6, Sdynv6, Zdynv6, Geynv6;
wire Neynv6, Ueynv6, Bfynv6, Ifynv6, Pfynv6, Wfynv6, Dgynv6, Kgynv6, Rgynv6, Ygynv6;
wire Fhynv6, Mhynv6, Thynv6, Aiynv6, Hiynv6, Oiynv6, Viynv6, Cjynv6, Jjynv6, Qjynv6;
wire Xjynv6, Ekynv6, Lkynv6, Skynv6, Zkynv6, Glynv6, Nlynv6, Ulynv6, Bmynv6, Imynv6;
wire Pmynv6, Wmynv6, Dnynv6, Knynv6, Rnynv6, Ynynv6, Foynv6, Moynv6, Toynv6, Apynv6;
wire Hpynv6, Opynv6, Vpynv6, Cqynv6, Jqynv6, Qqynv6, Xqynv6, Erynv6, Lrynv6, Srynv6;
wire Zrynv6, Gsynv6, Nsynv6, Usynv6, Btynv6, Itynv6, Ptynv6, Wtynv6, Duynv6, Kuynv6;
wire Ruynv6, Yuynv6, Fvynv6, Mvynv6, Tvynv6, Awynv6, Hwynv6, Owynv6, Vwynv6, Cxynv6;
wire Jxynv6, Qxynv6, Xxynv6, Eyynv6, Lyynv6, Syynv6, Zyynv6, Gzynv6, Nzynv6, Uzynv6;
wire B0znv6, I0znv6, P0znv6, W0znv6, D1znv6, K1znv6, R1znv6, Y1znv6, F2znv6, M2znv6;
wire T2znv6, A3znv6, H3znv6, O3znv6, V3znv6, C4znv6, J4znv6, Q4znv6, X4znv6, E5znv6;
wire L5znv6, S5znv6, Z5znv6, G6znv6, N6znv6, U6znv6, B7znv6, I7znv6, P7znv6, W7znv6;
wire D8znv6, K8znv6, R8znv6, Y8znv6, F9znv6, M9znv6, T9znv6, Aaznv6, Haznv6, Oaznv6;
wire Vaznv6, Cbznv6, Jbznv6, Qbznv6, Xbznv6, Ecznv6, Lcznv6, Scznv6, Zcznv6, Gdznv6;
wire Ndznv6, Udznv6, Beznv6, Ieznv6, Peznv6, Weznv6, Dfznv6, Kfznv6, Rfznv6, Yfznv6;
wire Fgznv6, Mgznv6, Tgznv6, Ahznv6, Hhznv6, Ohznv6, Vhznv6, Ciznv6, Jiznv6, Qiznv6;
wire Xiznv6, Ejznv6, Ljznv6, Sjznv6, Zjznv6, Gkznv6, Nkznv6, Ukznv6, Blznv6, Ilznv6;
wire Plznv6, Wlznv6, Dmznv6, Kmznv6, Rmznv6, Ymznv6, Fnznv6, Mnznv6, Tnznv6, Aoznv6;
wire Hoznv6, Ooznv6, Voznv6, Cpznv6, Jpznv6, Qpznv6, Xpznv6, Eqznv6, Lqznv6, Sqznv6;
wire Zqznv6, Grznv6, Nrznv6, Urznv6, Bsznv6, Isznv6, Psznv6, Wsznv6, Dtznv6, Ktznv6;
wire Rtznv6, Ytznv6, Fuznv6, Muznv6, Tuznv6, Avznv6, Hvznv6, Ovznv6, Vvznv6, Cwznv6;
wire Jwznv6, Qwznv6, Xwznv6, Exznv6, Lxznv6, Sxznv6, Zxznv6, Gyznv6, Nyznv6, Uyznv6;
wire Bzznv6, Izznv6, Pzznv6, Wzznv6, D00ov6, K00ov6, R00ov6, Y00ov6, F10ov6, M10ov6;
wire T10ov6, A20ov6, H20ov6, O20ov6, V20ov6, C30ov6, J30ov6, Q30ov6, X30ov6, E40ov6;
wire L40ov6, S40ov6, Z40ov6, G50ov6, N50ov6, U50ov6, B60ov6, I60ov6, P60ov6, W60ov6;
wire D70ov6, K70ov6, R70ov6, Y70ov6, F80ov6, M80ov6, T80ov6, A90ov6, H90ov6, O90ov6;
wire V90ov6, Ca0ov6, Ja0ov6, Qa0ov6, Xa0ov6, Eb0ov6, Lb0ov6, Sb0ov6, Zb0ov6, Gc0ov6;
wire Nc0ov6, Uc0ov6, Bd0ov6, Id0ov6, Pd0ov6, Wd0ov6, De0ov6, Ke0ov6, Re0ov6, Ye0ov6;
wire Ff0ov6, Mf0ov6, Tf0ov6, Ag0ov6, Hg0ov6, Og0ov6, Vg0ov6, Ch0ov6, Jh0ov6, Qh0ov6;
wire Xh0ov6, Ei0ov6, Li0ov6, Si0ov6, Zi0ov6, Gj0ov6, Nj0ov6, Uj0ov6, Bk0ov6, Ik0ov6;
wire Pk0ov6, Wk0ov6, Dl0ov6, Kl0ov6, Rl0ov6, Yl0ov6, Fm0ov6, Mm0ov6, Tm0ov6, An0ov6;
wire Hn0ov6, On0ov6, Vn0ov6, Co0ov6, Jo0ov6, Qo0ov6, Xo0ov6, Ep0ov6, Lp0ov6, Sp0ov6;
wire Zp0ov6, Gq0ov6, Nq0ov6, Uq0ov6, Br0ov6, Ir0ov6, Pr0ov6, Wr0ov6, Ds0ov6, Ks0ov6;
wire Rs0ov6, Ys0ov6, Ft0ov6, Mt0ov6, Tt0ov6, Au0ov6, Hu0ov6, Ou0ov6, Vu0ov6, Cv0ov6;
wire Jv0ov6, Qv0ov6, Xv0ov6, Ew0ov6, Lw0ov6, Sw0ov6, Zw0ov6, Gx0ov6, Nx0ov6, Ux0ov6;
wire By0ov6, Iy0ov6, Py0ov6, Wy0ov6, Dz0ov6, Kz0ov6, Rz0ov6, Yz0ov6, F01ov6, M01ov6;
wire T01ov6, A11ov6, H11ov6, O11ov6, V11ov6, C21ov6, J21ov6, Q21ov6, X21ov6, E31ov6;
wire L31ov6, S31ov6, Z31ov6, G41ov6, N41ov6, U41ov6, B51ov6, I51ov6, P51ov6, W51ov6;
wire D61ov6, K61ov6, R61ov6, Y61ov6, F71ov6, M71ov6, T71ov6, A81ov6, H81ov6, O81ov6;
wire V81ov6, C91ov6, J91ov6, Q91ov6, X91ov6, Ea1ov6, La1ov6, Sa1ov6, Za1ov6, Gb1ov6;
wire Nb1ov6, Ub1ov6, Bc1ov6, Ic1ov6, Pc1ov6, Wc1ov6, Dd1ov6, Kd1ov6, Rd1ov6, Yd1ov6;
wire Fe1ov6, Me1ov6, Te1ov6, Af1ov6, Hf1ov6, Of1ov6, Vf1ov6, Cg1ov6, Jg1ov6, Qg1ov6;
wire Xg1ov6, Eh1ov6, Lh1ov6, Sh1ov6, Zh1ov6, Gi1ov6, Ni1ov6, Ui1ov6, Bj1ov6, Ij1ov6;
wire Pj1ov6, Wj1ov6, Dk1ov6, Kk1ov6, Rk1ov6, Yk1ov6, Fl1ov6, Ml1ov6, Tl1ov6, Am1ov6;
wire Hm1ov6, Om1ov6, Vm1ov6, Cn1ov6, Jn1ov6, Qn1ov6, Xn1ov6, Eo1ov6, Lo1ov6, So1ov6;
wire Zo1ov6, Gp1ov6, Np1ov6, Up1ov6, Bq1ov6, Iq1ov6, Pq1ov6, Wq1ov6, Dr1ov6, Kr1ov6;
wire Rr1ov6, Yr1ov6, Fs1ov6, Ms1ov6, Ts1ov6, At1ov6, Ht1ov6, Ot1ov6, Vt1ov6, Cu1ov6;
wire Ju1ov6, Qu1ov6, Xu1ov6, Ev1ov6, Lv1ov6, Sv1ov6, Zv1ov6, Gw1ov6, Nw1ov6, Uw1ov6;
wire Bx1ov6, Ix1ov6, Px1ov6, Wx1ov6, Dy1ov6, Ky1ov6, Ry1ov6, Yy1ov6, Fz1ov6, Mz1ov6;
wire Tz1ov6, A02ov6, H02ov6, O02ov6, V02ov6, C12ov6, J12ov6, Q12ov6, X12ov6, E22ov6;
wire L22ov6, S22ov6, Z22ov6, G32ov6, N32ov6, U32ov6, B42ov6, I42ov6, P42ov6, W42ov6;
wire D52ov6, K52ov6, R52ov6, Y52ov6, F62ov6, M62ov6, T62ov6, A72ov6, H72ov6, O72ov6;
wire V72ov6, C82ov6, J82ov6, Q82ov6, X82ov6, E92ov6, L92ov6, S92ov6, Z92ov6, Ga2ov6;
wire Na2ov6, Ua2ov6, Bb2ov6, Ib2ov6, Pb2ov6, Wb2ov6, Dc2ov6, Kc2ov6, Rc2ov6, Yc2ov6;
wire Fd2ov6, Md2ov6, Td2ov6, Ae2ov6, He2ov6, Oe2ov6, Ve2ov6, Cf2ov6, Jf2ov6, Qf2ov6;
wire Xf2ov6, Eg2ov6, Lg2ov6, Sg2ov6, Zg2ov6, Gh2ov6, Nh2ov6, Uh2ov6, Bi2ov6, Ii2ov6;
wire Pi2ov6, Wi2ov6, Dj2ov6, Kj2ov6, Rj2ov6, Yj2ov6, Fk2ov6, Mk2ov6, Tk2ov6, Al2ov6;
wire Hl2ov6, Ol2ov6, Vl2ov6, Cm2ov6, Jm2ov6, Qm2ov6, Xm2ov6, En2ov6, Ln2ov6, Sn2ov6;
wire Zn2ov6, Go2ov6, No2ov6, Uo2ov6, Bp2ov6, Ip2ov6, Pp2ov6, Wp2ov6, Dq2ov6, Kq2ov6;
wire Rq2ov6, Yq2ov6, Fr2ov6, Mr2ov6, Tr2ov6, As2ov6, Hs2ov6, Os2ov6, Vs2ov6, Ct2ov6;
wire Jt2ov6, Qt2ov6, Xt2ov6, Eu2ov6, Lu2ov6, Su2ov6, Zu2ov6, Gv2ov6, Nv2ov6, Uv2ov6;
wire Bw2ov6, Iw2ov6, Pw2ov6, Ww2ov6, Dx2ov6, Kx2ov6, Rx2ov6, Yx2ov6, Fy2ov6, My2ov6;
wire Ty2ov6, Az2ov6, Hz2ov6, Oz2ov6, Vz2ov6, C03ov6, J03ov6, Q03ov6, X03ov6, E13ov6;
wire L13ov6, S13ov6, Z13ov6, G23ov6, N23ov6, U23ov6, B33ov6, I33ov6, P33ov6, W33ov6;
wire D43ov6, K43ov6, R43ov6, Y43ov6, F53ov6, M53ov6, T53ov6, A63ov6, H63ov6, O63ov6;
wire V63ov6, C73ov6, J73ov6, Q73ov6, X73ov6, E83ov6, L83ov6, S83ov6, Z83ov6, G93ov6;
wire N93ov6, U93ov6, Ba3ov6, Ia3ov6, Pa3ov6, Wa3ov6, Db3ov6, Kb3ov6, Rb3ov6, Yb3ov6;
wire Fc3ov6, Mc3ov6, Tc3ov6, Ad3ov6, Hd3ov6, Od3ov6, Vd3ov6, Ce3ov6, Je3ov6, Qe3ov6;
wire Xe3ov6, Ef3ov6, Lf3ov6, Sf3ov6, Zf3ov6, Gg3ov6, Ng3ov6, Ug3ov6, Bh3ov6, Ih3ov6;
wire Ph3ov6, Wh3ov6, Di3ov6, Ki3ov6, Ri3ov6, Yi3ov6, Fj3ov6, Mj3ov6, Tj3ov6, Ak3ov6;
wire Hk3ov6, Ok3ov6, Vk3ov6, Cl3ov6, Jl3ov6, Ql3ov6, Xl3ov6, Em3ov6, Lm3ov6, Sm3ov6;
wire Zm3ov6, Gn3ov6, Nn3ov6, Un3ov6, Bo3ov6, Io3ov6, Po3ov6, Wo3ov6, Dp3ov6, Kp3ov6;
wire Rp3ov6, Yp3ov6, Fq3ov6, Mq3ov6, Tq3ov6, Ar3ov6, Hr3ov6, Or3ov6, Vr3ov6, Cs3ov6;
wire Js3ov6, Qs3ov6, Xs3ov6, Et3ov6, Lt3ov6, St3ov6, Zt3ov6, Gu3ov6, Nu3ov6, Uu3ov6;
wire Bv3ov6, Iv3ov6, Pv3ov6, Wv3ov6, Dw3ov6, Kw3ov6, Rw3ov6, Yw3ov6, Fx3ov6, Mx3ov6;
wire Tx3ov6, Ay3ov6, Hy3ov6, Oy3ov6, Vy3ov6, Cz3ov6, Jz3ov6, Qz3ov6, Xz3ov6, E04ov6;
wire L04ov6, S04ov6, Z04ov6, G14ov6, N14ov6, U14ov6, B24ov6, I24ov6, P24ov6, W24ov6;
wire D34ov6, K34ov6, R34ov6, Y34ov6, F44ov6, M44ov6, T44ov6, A54ov6, H54ov6, O54ov6;
wire V54ov6, C64ov6, J64ov6, Q64ov6, X64ov6, E74ov6, L74ov6, S74ov6, Z74ov6, G84ov6;
wire N84ov6, U84ov6, B94ov6, I94ov6, P94ov6, W94ov6, Da4ov6, Ka4ov6, Ra4ov6, Ya4ov6;
wire Fb4ov6, Mb4ov6, Tb4ov6, Ac4ov6, Hc4ov6, Oc4ov6, Vc4ov6, Cd4ov6, Jd4ov6, Qd4ov6;
wire Xd4ov6, Ee4ov6, Le4ov6, Se4ov6, Ze4ov6, Gf4ov6, Nf4ov6, Uf4ov6, Bg4ov6, Ig4ov6;
wire Pg4ov6, Wg4ov6, Dh4ov6, Kh4ov6, Rh4ov6, Yh4ov6, Fi4ov6, Mi4ov6, Ti4ov6, Aj4ov6;
wire Hj4ov6, Oj4ov6, Vj4ov6, Ck4ov6, Jk4ov6, Qk4ov6, Xk4ov6, El4ov6, Ll4ov6, Sl4ov6;
wire Zl4ov6, Gm4ov6, Nm4ov6, Um4ov6, Bn4ov6, In4ov6, Pn4ov6, Wn4ov6, Do4ov6, Ko4ov6;
wire Ro4ov6, Yo4ov6, Fp4ov6, Mp4ov6, Tp4ov6, Aq4ov6, Hq4ov6, Oq4ov6, Vq4ov6, Cr4ov6;
wire Jr4ov6, Qr4ov6, Xr4ov6, Es4ov6, Ls4ov6, Ss4ov6, Zs4ov6, Gt4ov6, Nt4ov6, Ut4ov6;
wire Bu4ov6, Iu4ov6, Pu4ov6, Wu4ov6, Dv4ov6, Kv4ov6, Rv4ov6, Yv4ov6, Fw4ov6, Mw4ov6;
wire Tw4ov6, Ax4ov6, Hx4ov6, Ox4ov6, Vx4ov6, Cy4ov6, Jy4ov6, Qy4ov6, Xy4ov6, Ez4ov6;
wire Lz4ov6, Sz4ov6, Zz4ov6, G05ov6, N05ov6, U05ov6, B15ov6, I15ov6, P15ov6, W15ov6;
wire D25ov6, K25ov6, R25ov6, Y25ov6, F35ov6, M35ov6, T35ov6, A45ov6, H45ov6, O45ov6;
wire V45ov6, C55ov6, J55ov6, Q55ov6, X55ov6, E65ov6, L65ov6, S65ov6, Z65ov6, G75ov6;
wire N75ov6, U75ov6, B85ov6, I85ov6, P85ov6, W85ov6, D95ov6, K95ov6, R95ov6, Y95ov6;
wire Fa5ov6, Ma5ov6, Ta5ov6, Ab5ov6, Hb5ov6, Ob5ov6, Vb5ov6, Cc5ov6, Jc5ov6, Qc5ov6;
wire Xc5ov6, Ed5ov6, Ld5ov6, Sd5ov6, Zd5ov6, Ge5ov6, Ne5ov6, Ue5ov6, Bf5ov6, If5ov6;
wire Pf5ov6, Wf5ov6, Dg5ov6, Kg5ov6, Rg5ov6, Yg5ov6, Fh5ov6, Mh5ov6, Th5ov6, Ai5ov6;
wire Hi5ov6, Oi5ov6, Vi5ov6, Cj5ov6, Jj5ov6, Qj5ov6, Xj5ov6, Ek5ov6, Lk5ov6, Sk5ov6;
wire Zk5ov6, Gl5ov6, Nl5ov6, Ul5ov6, Bm5ov6, Im5ov6, Pm5ov6, Wm5ov6, Dn5ov6, Kn5ov6;
wire Rn5ov6, Yn5ov6, Fo5ov6, Mo5ov6, To5ov6, Ap5ov6, Hp5ov6, Op5ov6, Vp5ov6, Cq5ov6;
wire Jq5ov6, Qq5ov6, Xq5ov6, Er5ov6, Lr5ov6, Sr5ov6, Zr5ov6, Gs5ov6, Ns5ov6, Us5ov6;
wire Bt5ov6, It5ov6, Pt5ov6, Wt5ov6, Du5ov6, Ku5ov6, Ru5ov6, Yu5ov6, Fv5ov6, Mv5ov6;
wire Tv5ov6, Aw5ov6, Hw5ov6, Ow5ov6, Vw5ov6, Cx5ov6, Jx5ov6, Qx5ov6, Xx5ov6, Ey5ov6;
wire Ly5ov6, Sy5ov6, Zy5ov6, Gz5ov6, Nz5ov6, Uz5ov6, B06ov6, I06ov6, P06ov6, W06ov6;
wire D16ov6, K16ov6, R16ov6, Y16ov6, F26ov6, M26ov6, T26ov6, A36ov6, H36ov6, O36ov6;
wire V36ov6, C46ov6, J46ov6, Q46ov6, X46ov6, E56ov6, L56ov6, S56ov6, Z56ov6, G66ov6;
wire N66ov6, U66ov6, B76ov6, I76ov6, P76ov6, W76ov6, D86ov6, K86ov6, R86ov6, Y86ov6;
wire F96ov6, M96ov6, T96ov6, Aa6ov6, Ha6ov6, Oa6ov6, Va6ov6, Cb6ov6, Jb6ov6, Qb6ov6;
wire Xb6ov6, Ec6ov6, Lc6ov6, Sc6ov6, Zc6ov6, Gd6ov6, Nd6ov6, Ud6ov6, Be6ov6, Ie6ov6;
wire Pe6ov6, We6ov6, Df6ov6, Kf6ov6, Rf6ov6, Yf6ov6, Fg6ov6, Mg6ov6, Tg6ov6, Ah6ov6;
wire Hh6ov6, Oh6ov6, Vh6ov6, Ci6ov6, Ji6ov6, Qi6ov6, Xi6ov6, Ej6ov6, Lj6ov6, Sj6ov6;
wire Zj6ov6, Gk6ov6, Nk6ov6, Uk6ov6, Bl6ov6, Il6ov6, Pl6ov6, Wl6ov6, Dm6ov6, Km6ov6;
wire Rm6ov6, Ym6ov6, Fn6ov6, Mn6ov6, Tn6ov6, Ao6ov6, Ho6ov6, Oo6ov6, Vo6ov6, Cp6ov6;
wire Jp6ov6, Qp6ov6, Xp6ov6, Eq6ov6, Lq6ov6, Sq6ov6, Zq6ov6, Gr6ov6, Nr6ov6, Ur6ov6;
wire Bs6ov6, Is6ov6, Ps6ov6, Ws6ov6, Dt6ov6, Kt6ov6, Rt6ov6, Yt6ov6, Fu6ov6, Mu6ov6;
wire Tu6ov6, Av6ov6, Hv6ov6, Ov6ov6, Vv6ov6, Cw6ov6, Jw6ov6, Qw6ov6, Xw6ov6, Ex6ov6;
wire Lx6ov6, Sx6ov6, Zx6ov6, Gy6ov6, Ny6ov6, Uy6ov6, Bz6ov6, Iz6ov6, Pz6ov6, Wz6ov6;
wire D07ov6, K07ov6, R07ov6, Y07ov6, F17ov6, M17ov6, T17ov6, A27ov6, H27ov6, O27ov6;
wire V27ov6, C37ov6, J37ov6, Q37ov6, X37ov6, E47ov6, L47ov6, S47ov6, Z47ov6, G57ov6;
wire N57ov6, U57ov6, B67ov6, I67ov6, P67ov6, W67ov6, D77ov6, K77ov6, R77ov6, Y77ov6;
wire F87ov6, M87ov6, T87ov6, A97ov6, H97ov6, O97ov6, V97ov6, Ca7ov6, Ja7ov6, Qa7ov6;
wire Xa7ov6, Eb7ov6, Lb7ov6, Sb7ov6, Zb7ov6, Gc7ov6, Nc7ov6, Uc7ov6, Bd7ov6, Id7ov6;
wire Pd7ov6, Wd7ov6, De7ov6, Ke7ov6, Re7ov6, Ye7ov6, Ff7ov6, Mf7ov6, Tf7ov6, Ag7ov6;
wire Hg7ov6, Og7ov6, Vg7ov6, Ch7ov6, Jh7ov6, Qh7ov6, Xh7ov6, Ei7ov6, Li7ov6, Si7ov6;
wire Zi7ov6, Gj7ov6, Nj7ov6, Uj7ov6, Bk7ov6, Ik7ov6, Pk7ov6, Wk7ov6, Dl7ov6, Kl7ov6;
wire Rl7ov6, Yl7ov6, Fm7ov6, Mm7ov6, Tm7ov6, An7ov6, Hn7ov6, On7ov6, Vn7ov6, Co7ov6;
wire Jo7ov6, Qo7ov6, Xo7ov6, Ep7ov6, Lp7ov6, Sp7ov6, Zp7ov6, Gq7ov6, Nq7ov6, Uq7ov6;
wire Br7ov6, Ir7ov6, Pr7ov6, Wr7ov6, Ds7ov6, Ks7ov6, Rs7ov6, Ys7ov6, Ft7ov6, Mt7ov6;
wire Tt7ov6, Au7ov6, Hu7ov6, Ou7ov6, Vu7ov6, Cv7ov6, Jv7ov6, Qv7ov6, Xv7ov6, Ew7ov6;
wire Lw7ov6, Sw7ov6, Zw7ov6, Gx7ov6, Nx7ov6, Ux7ov6, By7ov6, Iy7ov6, Py7ov6, Wy7ov6;
wire Dz7ov6, Kz7ov6, Rz7ov6, Yz7ov6, F08ov6, M08ov6, T08ov6, A18ov6, H18ov6, O18ov6;
wire V18ov6, C28ov6, J28ov6, Q28ov6, X28ov6, E38ov6, L38ov6, S38ov6, Z38ov6, G48ov6;
wire N48ov6, U48ov6, B58ov6, I58ov6, P58ov6, W58ov6, D68ov6, K68ov6, R68ov6, Y68ov6;
wire F78ov6, M78ov6, T78ov6, A88ov6, H88ov6, O88ov6, V88ov6, C98ov6, J98ov6, Q98ov6;
wire X98ov6, Ea8ov6, La8ov6, Sa8ov6, Za8ov6, Gb8ov6, Nb8ov6, Ub8ov6, Bc8ov6, Ic8ov6;
wire Pc8ov6, Wc8ov6, Dd8ov6, Kd8ov6, Rd8ov6, Yd8ov6, Fe8ov6, Me8ov6, Te8ov6, Af8ov6;
wire Hf8ov6, Of8ov6, Vf8ov6, Cg8ov6, Jg8ov6, Qg8ov6, Xg8ov6, Eh8ov6, Lh8ov6, Sh8ov6;
wire Zh8ov6, Gi8ov6, Ni8ov6, Ui8ov6, Bj8ov6, Ij8ov6, Pj8ov6, Wj8ov6, Dk8ov6, Kk8ov6;
wire Rk8ov6, Yk8ov6, Fl8ov6, Ml8ov6, Tl8ov6, Am8ov6, Hm8ov6, Om8ov6, Vm8ov6, Cn8ov6;
wire Jn8ov6, Qn8ov6, Xn8ov6, Eo8ov6, Lo8ov6, So8ov6, Zo8ov6, Gp8ov6, Np8ov6, Up8ov6;
wire Bq8ov6, Iq8ov6, Pq8ov6, Wq8ov6, Dr8ov6, Kr8ov6, Rr8ov6, Yr8ov6, Fs8ov6, Ms8ov6;
wire Ts8ov6, At8ov6, Ht8ov6, Ot8ov6, Vt8ov6, Cu8ov6, Ju8ov6, Qu8ov6, Xu8ov6, Ev8ov6;
wire Lv8ov6, Sv8ov6, Zv8ov6, Gw8ov6, Nw8ov6, Uw8ov6, Bx8ov6, Ix8ov6, Px8ov6, Wx8ov6;
wire Dy8ov6, Ky8ov6, Ry8ov6, Yy8ov6, Fz8ov6, Mz8ov6, Tz8ov6, A09ov6, H09ov6, O09ov6;
wire V09ov6, C19ov6, J19ov6, Q19ov6, X19ov6, E29ov6, L29ov6, S29ov6, Z29ov6, G39ov6;
wire N39ov6, U39ov6, B49ov6, I49ov6, P49ov6, W49ov6, D59ov6, K59ov6, R59ov6, Y59ov6;
wire F69ov6, M69ov6, T69ov6, A79ov6, H79ov6, O79ov6, V79ov6, C89ov6, J89ov6, Q89ov6;
wire X89ov6, E99ov6, L99ov6, S99ov6, Z99ov6, Ga9ov6, Na9ov6, Ua9ov6, Bb9ov6, Ib9ov6;
wire Pb9ov6, Wb9ov6, Dc9ov6, Kc9ov6, Rc9ov6, Yc9ov6, Fd9ov6, Md9ov6, Td9ov6, Ae9ov6;
wire He9ov6, Oe9ov6, Ve9ov6, Cf9ov6, Jf9ov6, Qf9ov6, Xf9ov6, Eg9ov6, Lg9ov6, Sg9ov6;
wire Zg9ov6, Gh9ov6, Nh9ov6, Uh9ov6, Bi9ov6, Ii9ov6, Pi9ov6, Wi9ov6, Dj9ov6, Kj9ov6;
wire Rj9ov6, Yj9ov6, Fk9ov6, Mk9ov6, Tk9ov6, Al9ov6, Hl9ov6, Ol9ov6, Vl9ov6, Cm9ov6;
wire Jm9ov6, Qm9ov6, Xm9ov6, En9ov6, Ln9ov6, Sn9ov6, Zn9ov6, Go9ov6, No9ov6, Uo9ov6;
wire Bp9ov6, Ip9ov6, Pp9ov6, Wp9ov6, Dq9ov6, Kq9ov6, Rq9ov6, Yq9ov6, Fr9ov6, Mr9ov6;
wire Tr9ov6, As9ov6, Hs9ov6, Os9ov6, Vs9ov6, Ct9ov6, Jt9ov6, Qt9ov6, Xt9ov6, Eu9ov6;
wire Lu9ov6, Su9ov6, Zu9ov6, Gv9ov6, Nv9ov6, Uv9ov6, Bw9ov6, Iw9ov6, Pw9ov6, Ww9ov6;
wire Dx9ov6, Kx9ov6, Rx9ov6, Yx9ov6, Fy9ov6, My9ov6, Ty9ov6, Az9ov6, Hz9ov6, Oz9ov6;
wire Vz9ov6, C0aov6, J0aov6, Q0aov6, X0aov6, E1aov6, L1aov6, S1aov6, Z1aov6, G2aov6;
wire N2aov6, U2aov6, B3aov6, I3aov6, P3aov6, W3aov6, D4aov6, K4aov6, R4aov6, Y4aov6;
wire F5aov6, M5aov6, T5aov6, A6aov6, H6aov6, O6aov6, V6aov6, C7aov6, J7aov6, Q7aov6;
wire X7aov6, E8aov6, L8aov6, S8aov6, Z8aov6, G9aov6, N9aov6, U9aov6, Baaov6, Iaaov6;
wire Paaov6, Waaov6, Dbaov6, Kbaov6, Rbaov6, Ybaov6, Fcaov6, Mcaov6, Tcaov6, Adaov6;
wire Hdaov6, Odaov6, Vdaov6, Ceaov6, Jeaov6, Qeaov6, Xeaov6, Efaov6, Lfaov6, Sfaov6;
wire Zfaov6, Ggaov6, Ngaov6, Ugaov6, Bhaov6, Ihaov6, Phaov6, Whaov6, Diaov6, Kiaov6;
wire Riaov6, Yiaov6, Fjaov6, Mjaov6, Tjaov6, Akaov6, Hkaov6, Okaov6, Vkaov6, Claov6;
wire Jlaov6, Qlaov6, Xlaov6, Emaov6, Lmaov6, Smaov6, Zmaov6, Gnaov6, Nnaov6, Unaov6;
wire Boaov6, Ioaov6, Poaov6, Woaov6, Dpaov6, Kpaov6, Rpaov6, Ypaov6, Fqaov6, Mqaov6;
wire Tqaov6, Araov6, Hraov6, Oraov6, Vraov6, Csaov6, Jsaov6, Qsaov6, Xsaov6, Etaov6;
wire Ltaov6, Staov6, Ztaov6, Guaov6, Nuaov6, Uuaov6, Bvaov6, Ivaov6, Pvaov6, Wvaov6;
wire Dwaov6, Kwaov6, Rwaov6, Ywaov6, Fxaov6, Mxaov6, Txaov6, Ayaov6, Hyaov6, Oyaov6;
wire Vyaov6, Czaov6, Jzaov6, Qzaov6, Xzaov6, E0bov6, L0bov6, S0bov6, Z0bov6, G1bov6;
wire N1bov6, U1bov6, B2bov6, I2bov6, P2bov6, W2bov6, D3bov6, K3bov6, R3bov6, Y3bov6;
wire F4bov6, M4bov6, T4bov6, A5bov6, H5bov6, O5bov6, V5bov6, C6bov6, J6bov6, Q6bov6;
wire X6bov6, E7bov6, L7bov6, S7bov6, Z7bov6, G8bov6, N8bov6, U8bov6, B9bov6, I9bov6;
wire P9bov6, W9bov6, Dabov6, Kabov6, Rabov6, Yabov6, Fbbov6, Mbbov6, Tbbov6, Acbov6;
wire Hcbov6, Ocbov6, Vcbov6, Cdbov6, Jdbov6, Qdbov6, Xdbov6, Eebov6, Lebov6, Sebov6;
wire Zebov6, Gfbov6, Nfbov6, Ufbov6, Bgbov6, Igbov6, Pgbov6, Wgbov6, Dhbov6, Khbov6;
wire Rhbov6, Yhbov6, Fibov6, Mibov6, Tibov6, Ajbov6, Hjbov6, Ojbov6, Vjbov6, Ckbov6;
wire Jkbov6, Qkbov6, Xkbov6, Elbov6, Llbov6, Slbov6, Zlbov6, Gmbov6, Nmbov6, Umbov6;
wire Bnbov6, Inbov6, Pnbov6, Wnbov6, Dobov6, Kobov6, Robov6, Yobov6, Fpbov6, Mpbov6;
wire Tpbov6, Aqbov6, Hqbov6, Oqbov6, Vqbov6, Crbov6, Jrbov6, Qrbov6, Xrbov6, Esbov6;
wire Lsbov6, Ssbov6, Zsbov6, Gtbov6, Ntbov6, Utbov6, Bubov6, Iubov6, Pubov6, Wubov6;
wire Dvbov6, Kvbov6, Rvbov6, Yvbov6, Fwbov6, Mwbov6, Twbov6, Axbov6, Hxbov6, Oxbov6;
wire Vxbov6, Cybov6, Jybov6, Qybov6, Xybov6, Ezbov6, Lzbov6, Szbov6, Zzbov6, G0cov6;
wire N0cov6, U0cov6, B1cov6, I1cov6, P1cov6, W1cov6, D2cov6, K2cov6, R2cov6, Y2cov6;
wire F3cov6, M3cov6, T3cov6, A4cov6, H4cov6, O4cov6, V4cov6, C5cov6, J5cov6, Q5cov6;
wire X5cov6, E6cov6, L6cov6, S6cov6, Z6cov6, G7cov6, N7cov6, U7cov6, B8cov6, I8cov6;
wire P8cov6, W8cov6, D9cov6, K9cov6, R9cov6, Y9cov6, Facov6, Macov6, Tacov6, Abcov6;
wire Hbcov6, Obcov6, Vbcov6, Cccov6, Jccov6, Qccov6, Xccov6, Edcov6, Ldcov6, Sdcov6;
wire Zdcov6, Gecov6, Necov6, Uecov6, Bfcov6, Ifcov6, Pfcov6, Wfcov6, Dgcov6, Kgcov6;
wire Rgcov6, Ygcov6, Fhcov6, Mhcov6, Thcov6, Aicov6, Hicov6, Oicov6, Vicov6, Cjcov6;
wire Jjcov6, Qjcov6, Xjcov6, Ekcov6, Lkcov6, Skcov6, Zkcov6, Glcov6, Nlcov6, Ulcov6;
wire Bmcov6, Imcov6, Pmcov6, Wmcov6, Dncov6, Kncov6, Rncov6, Yncov6, Focov6, Mocov6;
wire Tocov6, Apcov6, Hpcov6, Opcov6, Vpcov6, Cqcov6, Jqcov6, Qqcov6, Xqcov6, Ercov6;
wire Lrcov6, Srcov6, Zrcov6, Gscov6, Nscov6, Uscov6, Btcov6, Itcov6, Ptcov6, Wtcov6;
wire Ducov6, Kucov6, Rucov6, Yucov6, Fvcov6, Mvcov6, Tvcov6, Awcov6, Hwcov6, Owcov6;
wire Vwcov6, Cxcov6, Jxcov6, Qxcov6, Xxcov6, Eycov6, Lycov6, Sycov6, Zycov6, Gzcov6;
wire Nzcov6, Uzcov6, B0dov6, I0dov6, P0dov6, W0dov6, D1dov6, K1dov6, R1dov6, Y1dov6;
wire F2dov6, M2dov6, T2dov6, A3dov6, H3dov6, O3dov6, V3dov6, C4dov6, J4dov6, Q4dov6;
wire X4dov6, E5dov6, L5dov6, S5dov6, Z5dov6, G6dov6, N6dov6, U6dov6, B7dov6, I7dov6;
wire P7dov6, W7dov6, D8dov6, K8dov6, R8dov6, Y8dov6, F9dov6, M9dov6, T9dov6, Aadov6;
wire Hadov6, Oadov6, Vadov6, Cbdov6, Jbdov6, Qbdov6, Xbdov6, Ecdov6, Lcdov6, Scdov6;
wire Zcdov6, Gddov6, Nddov6, Uddov6, Bedov6, Iedov6, Pedov6, Wedov6, Dfdov6, Kfdov6;
wire Rfdov6, Yfdov6, Fgdov6, Mgdov6, Tgdov6, Ahdov6, Hhdov6, Ohdov6, Vhdov6, Cidov6;
wire Jidov6, Qidov6, Xidov6, Ejdov6, Ljdov6, Sjdov6, Zjdov6, Gkdov6, Nkdov6, Ukdov6;
wire Bldov6, Ildov6, Pldov6, Wldov6, Dmdov6, Kmdov6, Rmdov6, Ymdov6, Fndov6, Mndov6;
wire Tndov6, Aodov6, Hodov6, Oodov6, Vodov6, Cpdov6, Jpdov6, Qpdov6, Xpdov6, Eqdov6;
wire Lqdov6, Sqdov6, Zqdov6, Grdov6, Nrdov6, Urdov6, Bsdov6, Isdov6, Psdov6, Wsdov6;
wire Dtdov6, Ktdov6, Rtdov6, Ytdov6, Fudov6, Mudov6, Tudov6, Avdov6, Hvdov6, Ovdov6;
wire Vvdov6, Cwdov6, Jwdov6, Qwdov6, Xwdov6, Exdov6, Lxdov6, Sxdov6, Zxdov6, Gydov6;
wire Nydov6, Uydov6, Bzdov6, Izdov6, Pzdov6, Wzdov6, D0eov6, K0eov6, R0eov6, Y0eov6;
wire F1eov6, M1eov6, T1eov6, A2eov6, H2eov6, O2eov6, V2eov6, C3eov6, J3eov6, Q3eov6;
wire X3eov6, E4eov6, L4eov6, S4eov6, Z4eov6, G5eov6, N5eov6, U5eov6, B6eov6, I6eov6;
wire P6eov6, W6eov6, D7eov6, K7eov6, R7eov6, Y7eov6, F8eov6, M8eov6, T8eov6, A9eov6;
wire H9eov6, O9eov6, V9eov6, Caeov6, Jaeov6, Qaeov6, Xaeov6, Ebeov6, Lbeov6, Sbeov6;
wire Zbeov6, Gceov6, Nceov6, Uceov6, Bdeov6, Ideov6, Pdeov6, Wdeov6, Deeov6, Keeov6;
wire Reeov6, Yeeov6, Ffeov6, Mfeov6, Tfeov6, Ageov6, Hgeov6, Ogeov6, Vgeov6, Cheov6;
wire Jheov6, Qheov6, Xheov6, Eieov6, Lieov6, Sieov6, Zieov6, Gjeov6, Njeov6, Ujeov6;
wire Bkeov6, Ikeov6, Pkeov6, Wkeov6, Dleov6, Kleov6, Rleov6, Yleov6, Fmeov6, Mmeov6;
wire Tmeov6, Aneov6, Hneov6, Oneov6, Vneov6, Coeov6, Joeov6, Qoeov6, Xoeov6, Epeov6;
wire Lpeov6, Speov6, Zpeov6, Gqeov6, Nqeov6, Uqeov6, Breov6, Ireov6, Preov6, Wreov6;
wire Dseov6, Kseov6, Rseov6, Yseov6, Fteov6, Mteov6, Tteov6, Aueov6, Hueov6, Oueov6;
wire Vueov6, Cveov6, Jveov6, Qveov6, Xveov6, Eweov6, Lweov6, Sweov6, Zweov6, Gxeov6;
wire Nxeov6, Uxeov6, Byeov6, Iyeov6, Pyeov6, Wyeov6, Dzeov6, Kzeov6, Rzeov6, Yzeov6;
wire F0fov6, M0fov6, T0fov6, A1fov6, H1fov6, O1fov6, V1fov6, C2fov6, J2fov6, Q2fov6;
wire X2fov6, E3fov6, L3fov6, S3fov6, Z3fov6, G4fov6, N4fov6, U4fov6, B5fov6, I5fov6;
wire P5fov6, W5fov6, D6fov6, K6fov6, R6fov6, Y6fov6, F7fov6, M7fov6, T7fov6, A8fov6;
wire H8fov6, O8fov6, V8fov6, C9fov6, J9fov6, Q9fov6, X9fov6, Eafov6, Lafov6, Safov6;
wire Zafov6, Gbfov6, Nbfov6, Ubfov6, Bcfov6, Icfov6, Pcfov6, Wcfov6, Ddfov6, Kdfov6;
wire Rdfov6, Ydfov6, Fefov6, Mefov6, Tefov6, Affov6, Hffov6, Offov6, Vffov6, Cgfov6;
wire Jgfov6, Qgfov6, Xgfov6, Ehfov6, Lhfov6, Shfov6, Zhfov6, Gifov6, Nifov6, Uifov6;
wire Bjfov6, Ijfov6, Pjfov6, Wjfov6, Dkfov6, Kkfov6, Rkfov6, Ykfov6, Flfov6, Mlfov6;
wire Tlfov6, Amfov6, Hmfov6, Omfov6, Vmfov6, Cnfov6, Jnfov6, Qnfov6, Xnfov6, Eofov6;
wire Lofov6, Sofov6, Zofov6, Gpfov6, Npfov6, Upfov6, Bqfov6, Iqfov6, Pqfov6, Wqfov6;
wire Drfov6, Krfov6, Rrfov6, Yrfov6, Fsfov6, Msfov6, Tsfov6, Atfov6, Htfov6, Otfov6;
wire Vtfov6, Cufov6, Jufov6, Qufov6, Xufov6, Evfov6, Lvfov6, Svfov6, Zvfov6, Gwfov6;
wire Nwfov6, Uwfov6, Bxfov6, Ixfov6, Pxfov6, Wxfov6, Dyfov6, Kyfov6, Ryfov6, Yyfov6;
wire Fzfov6, Mzfov6, Tzfov6, A0gov6, H0gov6, O0gov6, V0gov6, C1gov6, J1gov6, Q1gov6;
wire X1gov6, E2gov6, L2gov6, S2gov6, Z2gov6, G3gov6, N3gov6, U3gov6, B4gov6, I4gov6;
wire P4gov6, W4gov6, D5gov6, K5gov6, R5gov6, Y5gov6, F6gov6, M6gov6, T6gov6, A7gov6;
wire H7gov6, O7gov6, V7gov6, C8gov6, J8gov6, Q8gov6, X8gov6, E9gov6, L9gov6, S9gov6;
wire Z9gov6, Gagov6, Nagov6, Uagov6, Bbgov6, Ibgov6, Pbgov6, Wbgov6, Dcgov6, Kcgov6;
wire Rcgov6, Ycgov6, Fdgov6, Mdgov6, Tdgov6, Aegov6, Hegov6, Oegov6, Vegov6, Cfgov6;
wire Jfgov6, Qfgov6, Xfgov6, Eggov6, Lggov6, Sggov6, Zggov6, Ghgov6, Nhgov6, Uhgov6;
wire Bigov6, Iigov6, Pigov6, Wigov6, Djgov6, Kjgov6, Rjgov6, Yjgov6, Fkgov6, Mkgov6;
wire Tkgov6, Algov6, Hlgov6, Olgov6, Vlgov6, Cmgov6, Jmgov6, Qmgov6, Xmgov6, Engov6;
wire Lngov6, Sngov6, Zngov6, Gogov6, Nogov6, Uogov6, Bpgov6, Ipgov6, Ppgov6, Wpgov6;
wire Dqgov6, Kqgov6, Rqgov6, Yqgov6, Frgov6, Mrgov6, Trgov6, Asgov6, Hsgov6, Osgov6;
wire Vsgov6, Ctgov6, Jtgov6, Qtgov6, Xtgov6, Eugov6, Lugov6, Sugov6, Zugov6, Gvgov6;
wire Nvgov6, Uvgov6, Bwgov6, Iwgov6, Pwgov6, Wwgov6, Dxgov6, Kxgov6, Rxgov6, Yxgov6;
wire Fygov6, Mygov6, Tygov6, Azgov6, Hzgov6, Ozgov6, Vzgov6, C0hov6, J0hov6, Q0hov6;
wire X0hov6, E1hov6, L1hov6, S1hov6, Z1hov6, G2hov6, N2hov6, U2hov6, B3hov6, I3hov6;
wire P3hov6, W3hov6, D4hov6, K4hov6, R4hov6, Y4hov6, F5hov6, M5hov6, T5hov6, A6hov6;
wire H6hov6, O6hov6, V6hov6, C7hov6, J7hov6, Q7hov6, X7hov6, E8hov6, L8hov6, S8hov6;
wire Z8hov6, G9hov6, N9hov6, U9hov6, Bahov6, Iahov6, Pahov6, Wahov6, Dbhov6, Kbhov6;
wire Rbhov6, Ybhov6, Fchov6, Mchov6, Tchov6, Adhov6, Hdhov6, Odhov6, Vdhov6, Cehov6;
wire Jehov6, Qehov6, Xehov6, Efhov6, Lfhov6, Sfhov6, Zfhov6, Gghov6, Nghov6, Ughov6;
wire Bhhov6, Ihhov6, Phhov6, Whhov6, Dihov6, Kihov6, Rihov6, Yihov6, Fjhov6, Mjhov6;
wire Tjhov6, Akhov6, Hkhov6, Okhov6, Vkhov6, Clhov6, Jlhov6, Qlhov6, Xlhov6, Emhov6;
wire Lmhov6, Smhov6, Zmhov6, Gnhov6, Nnhov6, Unhov6, Bohov6, Iohov6, Pohov6, Wohov6;
wire Dphov6, Kphov6, Rphov6, Yphov6, Fqhov6, Mqhov6, Tqhov6, Arhov6, Hrhov6, Orhov6;
wire Vrhov6, Cshov6, Jshov6, Qshov6, Xshov6, Ethov6, Lthov6, Sthov6, Zthov6, Guhov6;
wire Nuhov6, Uuhov6, Bvhov6, Ivhov6, Pvhov6, Wvhov6, Dwhov6, Kwhov6, Rwhov6, Ywhov6;
wire Fxhov6, Mxhov6, Txhov6, Ayhov6, Hyhov6, Oyhov6, Vyhov6, Czhov6, Jzhov6, Qzhov6;
wire Xzhov6, E0iov6, L0iov6, S0iov6, Z0iov6, G1iov6, N1iov6, U1iov6, B2iov6, I2iov6;
wire P2iov6, W2iov6, D3iov6, K3iov6, R3iov6, Y3iov6, F4iov6, M4iov6, T4iov6, A5iov6;
wire H5iov6, O5iov6, V5iov6, C6iov6, J6iov6, Q6iov6, X6iov6, E7iov6, L7iov6, S7iov6;
wire Z7iov6, G8iov6, N8iov6, U8iov6, B9iov6, I9iov6, P9iov6, W9iov6, Daiov6, Kaiov6;
wire Raiov6, Yaiov6, Fbiov6, Mbiov6, Tbiov6, Aciov6, Hciov6, Ociov6, Vciov6, Cdiov6;
wire Jdiov6, Qdiov6, Xdiov6, Eeiov6, Leiov6, Seiov6, Zeiov6, Gfiov6, Nfiov6, Ufiov6;
wire Bgiov6, Igiov6, Pgiov6, Wgiov6, Dhiov6, Khiov6, Rhiov6, Yhiov6, Fiiov6, Miiov6;
wire Tiiov6, Ajiov6, Hjiov6, Ojiov6, Vjiov6, Ckiov6, Jkiov6, Qkiov6, Xkiov6, Eliov6;
wire Lliov6, Sliov6, Zliov6, Gmiov6, Nmiov6, Umiov6, Bniov6, Iniov6, Pniov6, Wniov6;
wire Doiov6, Koiov6, Roiov6, Yoiov6, Fpiov6, Mpiov6, Tpiov6, Aqiov6, Hqiov6, Oqiov6;
wire Vqiov6, Criov6, Jriov6, Qriov6, Xriov6, Esiov6, Lsiov6, Ssiov6, Zsiov6, Gtiov6;
wire Ntiov6, Utiov6, Buiov6, Iuiov6, Puiov6, Wuiov6, Dviov6, Kviov6, Rviov6, Yviov6;
wire Fwiov6, Mwiov6, Twiov6, Axiov6, Hxiov6, Oxiov6, Vxiov6, Cyiov6, Jyiov6, Qyiov6;
wire Xyiov6, Eziov6, Lziov6, Sziov6, Zziov6, G0jov6, N0jov6, U0jov6, B1jov6, I1jov6;
wire P1jov6, W1jov6, D2jov6, K2jov6, R2jov6, Y2jov6, F3jov6, M3jov6, T3jov6, A4jov6;
wire H4jov6, O4jov6, V4jov6, C5jov6, J5jov6, Q5jov6, X5jov6, E6jov6, L6jov6, S6jov6;
wire Z6jov6, G7jov6, N7jov6, U7jov6, B8jov6, I8jov6, P8jov6, W8jov6, D9jov6, K9jov6;
wire R9jov6, Y9jov6, Fajov6, Majov6, Tajov6, Abjov6, Hbjov6, Objov6, Vbjov6, Ccjov6;
wire Jcjov6, Qcjov6, Xcjov6, Edjov6, Ldjov6, Sdjov6, Zdjov6, Gejov6, Nejov6, Uejov6;
wire Bfjov6, Ifjov6, Pfjov6, Wfjov6, Dgjov6, Kgjov6, Rgjov6, Ygjov6, Fhjov6, Mhjov6;
wire Thjov6, Aijov6, Hijov6, Oijov6, Vijov6, Cjjov6, Jjjov6, Qjjov6, Xjjov6, Ekjov6;
wire Lkjov6, Skjov6, Zkjov6, Gljov6, Nljov6, Uljov6, Bmjov6, Imjov6, Pmjov6, Wmjov6;
wire Dnjov6, Knjov6, Rnjov6, Ynjov6, Fojov6, Mojov6, Tojov6, Apjov6, Hpjov6, Opjov6;
wire Vpjov6, Cqjov6, Jqjov6, Qqjov6, Xqjov6, Erjov6, Lrjov6, Srjov6, Zrjov6, Gsjov6;
wire Nsjov6, Usjov6, Btjov6, Itjov6, Ptjov6, Wtjov6, Dujov6, Kujov6, Rujov6, Yujov6;
wire Fvjov6, Mvjov6, Tvjov6, Awjov6, Hwjov6, Owjov6, Vwjov6, Cxjov6, Jxjov6, Qxjov6;
wire Xxjov6, Eyjov6, Lyjov6, Syjov6, Zyjov6, Gzjov6, Nzjov6, Uzjov6, B0kov6, I0kov6;
wire P0kov6, W0kov6, D1kov6, K1kov6, R1kov6, Y1kov6, F2kov6, M2kov6, T2kov6, A3kov6;
wire H3kov6, O3kov6, V3kov6, C4kov6, J4kov6, Q4kov6, X4kov6, E5kov6, L5kov6, S5kov6;
wire Z5kov6, G6kov6, N6kov6, U6kov6, B7kov6, I7kov6, P7kov6, W7kov6, D8kov6, K8kov6;
wire R8kov6, Y8kov6, F9kov6, M9kov6, T9kov6, Aakov6, Hakov6, Oakov6, Vakov6, Cbkov6;
wire Jbkov6, Qbkov6, Xbkov6, Eckov6, Lckov6, Sckov6, Zckov6, Gdkov6, Ndkov6, Udkov6;
wire Bekov6, Iekov6, Pekov6, Wekov6, Dfkov6, Kfkov6, Rfkov6, Yfkov6, Fgkov6, Mgkov6;
wire Tgkov6, Ahkov6, Hhkov6, Ohkov6, Vhkov6, Cikov6, Jikov6, Qikov6, Xikov6, Ejkov6;
wire Ljkov6, Sjkov6, Zjkov6, Gkkov6, Nkkov6, Ukkov6, Blkov6, Ilkov6, Plkov6, Wlkov6;
wire Dmkov6, Kmkov6, Rmkov6, Ymkov6, Fnkov6, Mnkov6, Tnkov6, Aokov6, Hokov6, Ookov6;
wire Vokov6, Cpkov6, Jpkov6, Qpkov6, Xpkov6, Eqkov6, Lqkov6, Sqkov6, Zqkov6, Grkov6;
wire Nrkov6, Urkov6, Bskov6, Iskov6, Pskov6, Wskov6, Dtkov6, Ktkov6, Rtkov6, Ytkov6;
wire Fukov6, Mukov6, Tukov6, Avkov6, Hvkov6, Ovkov6, Vvkov6, Cwkov6, Jwkov6, Qwkov6;
wire Xwkov6, Exkov6, Lxkov6, Sxkov6, Zxkov6, Gykov6, Nykov6, Uykov6, Bzkov6, Izkov6;
wire Pzkov6, Wzkov6, D0lov6, K0lov6, R0lov6, Y0lov6, F1lov6, M1lov6, T1lov6, A2lov6;
wire H2lov6, O2lov6, V2lov6, C3lov6, J3lov6, Q3lov6, X3lov6, E4lov6, L4lov6, S4lov6;
wire Z4lov6, G5lov6, N5lov6, U5lov6, B6lov6, I6lov6, P6lov6, W6lov6, D7lov6, K7lov6;
wire R7lov6, Y7lov6, F8lov6, M8lov6, T8lov6, A9lov6, H9lov6, O9lov6, V9lov6, Calov6;
wire Jalov6, Qalov6, Xalov6, Eblov6, Lblov6, Sblov6, Zblov6, Gclov6, Nclov6, Uclov6;
wire Bdlov6, Idlov6, Pdlov6, Wdlov6, Delov6, Kelov6, Relov6, Yelov6, Fflov6, Mflov6;
wire Tflov6, Aglov6, Hglov6, Oglov6, Vglov6, Chlov6, Jhlov6, Qhlov6, Xhlov6, Eilov6;
wire Lilov6, Silov6, Zilov6, Gjlov6, Njlov6, Ujlov6, Bklov6, Iklov6, Pklov6, Wklov6;
wire Dllov6, Kllov6, Rllov6, Yllov6, Fmlov6, Mmlov6, Tmlov6, Anlov6, Hnlov6, Onlov6;
wire Vnlov6, Colov6, Jolov6, Qolov6, Xolov6, Eplov6, Lplov6, Splov6, Zplov6, Gqlov6;
wire Nqlov6, Uqlov6, Brlov6, Irlov6, Prlov6, Wrlov6, Dslov6, Kslov6, Rslov6, Yslov6;
wire Ftlov6, Mtlov6, Ttlov6, Aulov6, Hulov6, Oulov6, Vulov6, Cvlov6, Jvlov6, Qvlov6;
wire Xvlov6, Ewlov6, Lwlov6, Swlov6, Zwlov6, Gxlov6, Nxlov6, Uxlov6, Bylov6, Iylov6;
wire Pylov6, Wylov6, Dzlov6, Kzlov6, Rzlov6, Yzlov6, F0mov6, M0mov6, T0mov6, A1mov6;
wire H1mov6, O1mov6, V1mov6, C2mov6, J2mov6, Q2mov6, X2mov6, E3mov6, L3mov6, S3mov6;
wire Z3mov6, G4mov6, N4mov6, U4mov6, B5mov6, I5mov6, P5mov6, W5mov6, D6mov6, K6mov6;
wire R6mov6, Y6mov6, F7mov6, M7mov6, T7mov6, A8mov6, H8mov6, O8mov6, V8mov6, C9mov6;
wire J9mov6, Q9mov6, X9mov6, Eamov6, Lamov6, Samov6, Zamov6, Gbmov6, Nbmov6, Ubmov6;
wire Bcmov6, Icmov6, Pcmov6, Wcmov6, Ddmov6, Kdmov6, Rdmov6, Ydmov6, Femov6, Memov6;
wire Temov6, Afmov6, Hfmov6, Ofmov6, Vfmov6, Cgmov6, Jgmov6, Qgmov6, Xgmov6, Ehmov6;
wire Lhmov6, Shmov6, Zhmov6, Gimov6, Nimov6, Uimov6, Bjmov6, Ijmov6, Pjmov6, Wjmov6;
wire Dkmov6, Kkmov6, Rkmov6, Ykmov6, Flmov6, Mlmov6, Tlmov6, Ammov6, Hmmov6, Ommov6;
wire Vmmov6, Cnmov6, Jnmov6, Qnmov6, Xnmov6, Eomov6, Lomov6, Somov6, Zomov6, Gpmov6;
wire Npmov6, Upmov6, Bqmov6, Iqmov6, Pqmov6, Wqmov6, Drmov6, Krmov6, Rrmov6, Yrmov6;
wire Fsmov6, Msmov6, Tsmov6, Atmov6, Htmov6, Otmov6, Vtmov6, Cumov6, Jumov6, Qumov6;
wire Xumov6, Evmov6, Lvmov6, Svmov6, Zvmov6, Gwmov6, Nwmov6, Uwmov6, Bxmov6, Ixmov6;
wire Pxmov6, Wxmov6, Dymov6, Kymov6, Rymov6, Yymov6, Fzmov6, Mzmov6, Tzmov6, A0nov6;
wire H0nov6, O0nov6, V0nov6, C1nov6, J1nov6, Q1nov6, X1nov6, E2nov6, L2nov6, S2nov6;
wire Z2nov6, G3nov6, N3nov6, U3nov6, B4nov6, I4nov6, P4nov6, W4nov6, D5nov6, K5nov6;
wire R5nov6, Y5nov6, F6nov6, M6nov6, T6nov6, A7nov6, H7nov6, O7nov6, V7nov6, C8nov6;
wire J8nov6, Q8nov6, X8nov6, E9nov6, L9nov6, S9nov6, Z9nov6, Ganov6, Nanov6, Uanov6;
wire Bbnov6, Ibnov6, Pbnov6, Wbnov6, Dcnov6, Kcnov6, Rcnov6, Ycnov6, Fdnov6, Mdnov6;
wire Tdnov6, Aenov6, Henov6, Oenov6, Venov6, Cfnov6, Jfnov6, Qfnov6, Xfnov6, Egnov6;
wire Lgnov6, Sgnov6, Zgnov6, Ghnov6, Nhnov6, Uhnov6, Binov6, Iinov6, Pinov6, Winov6;
wire Djnov6, Kjnov6, Rjnov6, Yjnov6, Fknov6, Mknov6, Tknov6, Alnov6, Hlnov6, Olnov6;
wire Vlnov6, Cmnov6, Jmnov6, Qmnov6, Xmnov6, Ennov6, Lnnov6, Snnov6, Znnov6, Gonov6;
wire Nonov6, Uonov6, Bpnov6, Ipnov6, Ppnov6, Wpnov6, Dqnov6, Kqnov6, Rqnov6, Yqnov6;
wire Frnov6, Mrnov6, Trnov6, Asnov6, Hsnov6, Osnov6, Vsnov6, Ctnov6, Jtnov6, Qtnov6;
wire Xtnov6, Eunov6, Lunov6, Sunov6, Zunov6, Gvnov6, Nvnov6, Uvnov6, Bwnov6, Iwnov6;
wire Pwnov6, Wwnov6, Dxnov6, Kxnov6, Rxnov6, Yxnov6, Fynov6, Mynov6, Tynov6, Aznov6;
wire Hznov6, Oznov6, Vznov6, C0oov6, J0oov6, Q0oov6, X0oov6, E1oov6, L1oov6, S1oov6;
wire Z1oov6, G2oov6, N2oov6, U2oov6, B3oov6, I3oov6, P3oov6, W3oov6, D4oov6, K4oov6;
wire R4oov6, Y4oov6, F5oov6, M5oov6, T5oov6, A6oov6, H6oov6, O6oov6, V6oov6, C7oov6;
wire J7oov6, Q7oov6, X7oov6, E8oov6, L8oov6, S8oov6, Z8oov6, G9oov6, N9oov6, U9oov6;
wire Baoov6, Iaoov6, Paoov6, Waoov6, Dboov6, Kboov6, Rboov6, Yboov6, Fcoov6, Mcoov6;
wire Tcoov6, Adoov6, Hdoov6, Odoov6, Vdoov6, Ceoov6, Jeoov6, Qeoov6, Xeoov6, Efoov6;
wire Lfoov6, Sfoov6, Zfoov6, Ggoov6, Ngoov6, Ugoov6, Bhoov6, Ihoov6, Phoov6, Whoov6;
wire Dioov6, Kioov6, Rioov6, Yioov6, Fjoov6, Mjoov6, Tjoov6, Akoov6, Hkoov6, Okoov6;
wire Vkoov6, Cloov6, Jloov6, Qloov6, Xloov6, Emoov6, Lmoov6, Smoov6, Zmoov6, Gnoov6;
wire Nnoov6, Unoov6, Booov6, Iooov6, Pooov6, Wooov6, Dpoov6, Kpoov6, Rpoov6, Ypoov6;
wire Fqoov6, Mqoov6, Tqoov6, Aroov6, Hroov6, Oroov6, Vroov6, Csoov6, Jsoov6, Qsoov6;
wire Xsoov6, Etoov6, Ltoov6, Stoov6, Ztoov6, Guoov6, Nuoov6, Uuoov6, Bvoov6, Ivoov6;
wire Pvoov6, Wvoov6, Dwoov6, Kwoov6, Rwoov6, Ywoov6, Fxoov6, Mxoov6, Txoov6, Ayoov6;
wire Hyoov6, Oyoov6, Vyoov6, Czoov6, Jzoov6, Qzoov6, Xzoov6, E0pov6, L0pov6, S0pov6;
wire Z0pov6, G1pov6, N1pov6, U1pov6, B2pov6, I2pov6, P2pov6, W2pov6, D3pov6, K3pov6;
wire R3pov6, Y3pov6, F4pov6, M4pov6, T4pov6, A5pov6, H5pov6, O5pov6, V5pov6, C6pov6;
wire J6pov6, Q6pov6, X6pov6, E7pov6, L7pov6, S7pov6, Z7pov6, G8pov6, N8pov6, U8pov6;
wire B9pov6, I9pov6, P9pov6, W9pov6, Dapov6, Kapov6, Rapov6, Yapov6, Fbpov6, Mbpov6;
wire Tbpov6, Acpov6, Hcpov6, Ocpov6, Vcpov6, Cdpov6, Jdpov6, Qdpov6, Xdpov6, Eepov6;
wire Lepov6, Sepov6, Zepov6, Gfpov6, Nfpov6, Ufpov6, Bgpov6, Igpov6, Pgpov6, Wgpov6;
wire Dhpov6, Khpov6, Rhpov6, Yhpov6, Fipov6, Mipov6, Tipov6, Ajpov6, Hjpov6, Ojpov6;
wire Vjpov6, Ckpov6, Jkpov6, Qkpov6, Xkpov6, Elpov6, Llpov6, Slpov6, Zlpov6, Gmpov6;
wire Nmpov6, Umpov6, Bnpov6, Inpov6, Pnpov6, Wnpov6, Dopov6, Kopov6, Ropov6, Yopov6;
wire Fppov6, Mppov6, Tppov6, Aqpov6, Hqpov6, Oqpov6, Vqpov6, Crpov6, Jrpov6, Qrpov6;
wire Xrpov6, Espov6, Lspov6, Sspov6, Zspov6, Gtpov6, Ntpov6, Utpov6, Bupov6, Iupov6;
wire Pupov6, Wupov6, Dvpov6, Kvpov6, Rvpov6, Yvpov6, Fwpov6, Mwpov6, Twpov6, Axpov6;
wire Hxpov6, Oxpov6, Vxpov6, Cypov6, Jypov6, Qypov6, Xypov6, Ezpov6, Lzpov6, Szpov6;
wire Zzpov6, G0qov6, N0qov6, U0qov6, B1qov6, I1qov6, P1qov6, W1qov6, D2qov6, K2qov6;
wire R2qov6, Y2qov6, F3qov6, M3qov6, T3qov6, A4qov6, H4qov6, O4qov6, V4qov6, C5qov6;
wire J5qov6, Q5qov6, X5qov6, E6qov6, L6qov6, S6qov6, Z6qov6, G7qov6, N7qov6, U7qov6;
wire B8qov6, I8qov6, P8qov6, W8qov6, D9qov6, K9qov6, R9qov6, Y9qov6, Faqov6, Maqov6;
wire Taqov6, Abqov6, Hbqov6, Obqov6, Vbqov6, Ccqov6, Jcqov6, Qcqov6, Xcqov6, Edqov6;
wire Ldqov6, Sdqov6, Zdqov6, Geqov6, Neqov6, Ueqov6, Bfqov6, Ifqov6, Pfqov6, Wfqov6;
wire Dgqov6, Kgqov6, Rgqov6, Ygqov6, Fhqov6, Mhqov6, Thqov6, Aiqov6, Hiqov6, Oiqov6;
wire Viqov6, Cjqov6, Jjqov6, Qjqov6, Xjqov6, Ekqov6, Lkqov6, Skqov6, Zkqov6, Glqov6;
wire Nlqov6, Ulqov6, Bmqov6, Imqov6, Pmqov6, Wmqov6, Dnqov6, Knqov6, Rnqov6, Ynqov6;
wire Foqov6, Moqov6, Toqov6, Apqov6, Hpqov6, Opqov6, Vpqov6, Cqqov6, Jqqov6, Qqqov6;
wire Xqqov6, Erqov6, Lrqov6, Srqov6, Zrqov6, Gsqov6, Nsqov6, Usqov6, Btqov6, Itqov6;
wire Ptqov6, Wtqov6, Duqov6, Kuqov6, Ruqov6, Yuqov6, Fvqov6, Mvqov6, Tvqov6, Awqov6;
wire Hwqov6, Owqov6, Vwqov6, Cxqov6, Jxqov6, Qxqov6, Xxqov6, Eyqov6, Lyqov6, Syqov6;
wire Zyqov6, Gzqov6, Nzqov6, Uzqov6, B0rov6, I0rov6, P0rov6, W0rov6, D1rov6, K1rov6;
wire R1rov6, Y1rov6, F2rov6, M2rov6, T2rov6, A3rov6, H3rov6, O3rov6, V3rov6, C4rov6;
wire J4rov6, Q4rov6, X4rov6, E5rov6, L5rov6, S5rov6, Z5rov6, G6rov6, N6rov6, U6rov6;
wire B7rov6, I7rov6, P7rov6, W7rov6, D8rov6, K8rov6, R8rov6, Y8rov6, F9rov6, M9rov6;
wire T9rov6, Aarov6, Harov6, Oarov6, Varov6, Cbrov6, Jbrov6, Qbrov6, Xbrov6, Ecrov6;
wire Lcrov6, Scrov6, Zcrov6, Gdrov6, Ndrov6, Udrov6, Berov6, Ierov6, Perov6, Werov6;
wire Dfrov6, Kfrov6, Rfrov6, Yfrov6, Fgrov6, Mgrov6, Tgrov6, Ahrov6, Hhrov6, Ohrov6;
wire Vhrov6, Cirov6, Jirov6, Qirov6, Xirov6, Ejrov6, Ljrov6, Sjrov6, Zjrov6, Gkrov6;
wire Nkrov6, Ukrov6, Blrov6, Ilrov6, Plrov6, Wlrov6, Dmrov6, Kmrov6, Rmrov6, Ymrov6;
wire Fnrov6, Mnrov6, Tnrov6, Aorov6, Horov6, Oorov6, Vorov6, Cprov6, Jprov6, Qprov6;
wire Xprov6, Eqrov6, Lqrov6, Sqrov6, Zqrov6, Grrov6, Nrrov6, Urrov6, Bsrov6, Isrov6;
wire Psrov6, Wsrov6, Dtrov6, Ktrov6, Rtrov6, Ytrov6, Furov6, Murov6, Turov6, Avrov6;
wire Hvrov6, Ovrov6, Vvrov6, Cwrov6, Jwrov6, Qwrov6, Xwrov6, Exrov6, Lxrov6, Sxrov6;
wire Zxrov6, Gyrov6, Nyrov6, Uyrov6, Bzrov6, Izrov6, Pzrov6, Wzrov6, D0sov6, K0sov6;
wire R0sov6, Y0sov6, F1sov6, M1sov6, T1sov6, A2sov6, H2sov6, O2sov6, V2sov6, C3sov6;
wire J3sov6, Q3sov6, X3sov6, E4sov6, L4sov6, S4sov6, Z4sov6, G5sov6, N5sov6, U5sov6;
wire B6sov6, I6sov6, P6sov6, W6sov6, D7sov6, K7sov6, R7sov6, Y7sov6, F8sov6, M8sov6;
wire T8sov6, A9sov6, H9sov6, O9sov6, V9sov6, Casov6, Jasov6, Qasov6, Xasov6, Ebsov6;
wire Lbsov6, Sbsov6, Zbsov6, Gcsov6, Ncsov6, Ucsov6, Bdsov6, Idsov6, Pdsov6, Wdsov6;
wire Desov6, Kesov6, Resov6, Yesov6, Ffsov6, Mfsov6, Tfsov6, Agsov6, Hgsov6, Ogsov6;
wire Vgsov6, Chsov6, Jhsov6, Qhsov6, Xhsov6, Eisov6, Lisov6, Sisov6, Zisov6, Gjsov6;
wire Njsov6, Ujsov6, Bksov6, Iksov6, Pksov6, Wksov6, Dlsov6, Klsov6, Rlsov6, Ylsov6;
wire Fmsov6, Mmsov6, Tmsov6, Ansov6, Hnsov6, Onsov6, Vnsov6, Cosov6, Josov6, Qosov6;
wire Xosov6, Epsov6, Lpsov6, Spsov6, Zpsov6, Gqsov6, Nqsov6, Uqsov6, Brsov6, Irsov6;
wire Prsov6, Wrsov6, Dssov6, Kssov6, Rssov6, Yssov6, Ftsov6, Mtsov6, Ttsov6, Ausov6;
wire Husov6, Ousov6, Vusov6, Cvsov6, Jvsov6, Qvsov6, Xvsov6, Ewsov6, Lwsov6, Swsov6;
wire Zwsov6, Gxsov6, Nxsov6, Uxsov6, Bysov6, Iysov6, Pysov6, Wysov6, Dzsov6, Kzsov6;
wire Rzsov6, Yzsov6, F0tov6, M0tov6, T0tov6, A1tov6, H1tov6, O1tov6, V1tov6, C2tov6;
wire J2tov6, Q2tov6, X2tov6, E3tov6, L3tov6, S3tov6, Z3tov6, G4tov6, N4tov6, U4tov6;
wire B5tov6, I5tov6, P5tov6, W5tov6, D6tov6, K6tov6, R6tov6, Y6tov6, F7tov6, M7tov6;
wire T7tov6, A8tov6, H8tov6, O8tov6, V8tov6, C9tov6, J9tov6, Q9tov6, X9tov6, Eatov6;
wire Latov6, Satov6, Zatov6, Gbtov6, Nbtov6, Ubtov6, Bctov6, Ictov6, Pctov6, Wctov6;
wire Ddtov6, Kdtov6, Rdtov6, Ydtov6, Fetov6, Metov6, Tetov6, Aftov6, Hftov6, Oftov6;
wire Vftov6, Cgtov6, Jgtov6, Qgtov6, Xgtov6, Ehtov6, Lhtov6, Shtov6, Zhtov6, Gitov6;
wire Nitov6, Uitov6, Bjtov6, Ijtov6, Pjtov6, Wjtov6, Dktov6, Kktov6, Rktov6, Yktov6;
wire Fltov6, Mltov6, Tltov6, Amtov6, Hmtov6, Omtov6, Vmtov6, Cntov6, Jntov6, Mmehw6;
wire Tmehw6, Anehw6, Hnehw6, Onehw6, Vnehw6, Coehw6, Joehw6, Qoehw6, Xoehw6, Epehw6;
wire Lpehw6, Spehw6, Zpehw6, Gqehw6, Nqehw6, Uqehw6, Brehw6, Irehw6, Prehw6, Wrehw6;
wire Dsehw6, Ksehw6, Rsehw6, Ysehw6, Ftehw6, Mtehw6, Ttehw6, Auehw6, Huehw6, Ouehw6;
wire Vuehw6, Cvehw6, Jvehw6, Qvehw6, Xvehw6, Ewehw6, Lwehw6, Swehw6, Zwehw6, Gxehw6;
wire Nxehw6, Uxehw6, Byehw6, Iyehw6, Pyehw6, Wyehw6, Dzehw6, Kzehw6, Rzehw6, Yzehw6;
wire F0fhw6, M0fhw6, T0fhw6, A1fhw6, H1fhw6, O1fhw6, V1fhw6, C2fhw6, J2fhw6, Q2fhw6;
wire X2fhw6, E3fhw6, L3fhw6, S3fhw6, Z3fhw6, G4fhw6, N4fhw6, U4fhw6, B5fhw6, I5fhw6;
wire P5fhw6, W5fhw6, D6fhw6, K6fhw6, R6fhw6, Y6fhw6, F7fhw6, M7fhw6, T7fhw6, A8fhw6;
wire H8fhw6, O8fhw6, V8fhw6, C9fhw6, J9fhw6, Q9fhw6, X9fhw6, Eafhw6, Lafhw6, Safhw6;
wire Zafhw6, Gbfhw6, Nbfhw6, Ubfhw6, Bcfhw6, Icfhw6, Pcfhw6, Wcfhw6, Ddfhw6, Kdfhw6;
wire Rdfhw6, Ydfhw6, Fefhw6, Mefhw6, Tefhw6, Affhw6, Hffhw6, Offhw6, Vffhw6, Cgfhw6;
wire Jgfhw6, Qgfhw6, Xgfhw6, Ehfhw6, Lhfhw6, Shfhw6, Zhfhw6, Gifhw6, Nifhw6, Uifhw6;
wire Bjfhw6, Ijfhw6, Pjfhw6, Wjfhw6, Dkfhw6, Kkfhw6, Rkfhw6, Ykfhw6, Flfhw6, Mlfhw6;
wire Tlfhw6, Amfhw6, Hmfhw6, Omfhw6, Vmfhw6, Cnfhw6, Jnfhw6, Qnfhw6, Xnfhw6, Eofhw6;
wire Lofhw6, Sofhw6, Zofhw6, Gpfhw6, Npfhw6, Upfhw6, Bqfhw6, Iqfhw6, Pqfhw6, Wqfhw6;
wire Drfhw6, Krfhw6, Rrfhw6, Yrfhw6, Fsfhw6, Msfhw6, Tsfhw6, Atfhw6, Htfhw6, Otfhw6;
wire Vtfhw6, Cufhw6, Jufhw6, Qufhw6, Xufhw6, Evfhw6, Lvfhw6, Svfhw6, Zvfhw6, Gwfhw6;
wire Nwfhw6, Uwfhw6, Bxfhw6, Ixfhw6, Pxfhw6, Wxfhw6, Dyfhw6, Kyfhw6, Ryfhw6, Yyfhw6;
wire Fzfhw6, Mzfhw6, Tzfhw6, A0ghw6, H0ghw6, O0ghw6, V0ghw6, C1ghw6, J1ghw6, Q1ghw6;
wire X1ghw6, E2ghw6, L2ghw6, S2ghw6, Z2ghw6, G3ghw6, N3ghw6, U3ghw6, B4ghw6, I4ghw6;
wire P4ghw6, W4ghw6, D5ghw6, K5ghw6, R5ghw6, Y5ghw6, F6ghw6, M6ghw6, T6ghw6, A7ghw6;
wire H7ghw6, O7ghw6, V7ghw6, C8ghw6, J8ghw6, Q8ghw6, X8ghw6, E9ghw6, L9ghw6, S9ghw6;
wire Z9ghw6, Gaghw6, Naghw6, Uaghw6, Bbghw6, Ibghw6, Pbghw6, Wbghw6, Dcghw6, Kcghw6;
wire Rcghw6, Ycghw6, Fdghw6, Mdghw6, Tdghw6, Aeghw6, Heghw6, Oeghw6, Veghw6, Cfghw6;
wire Jfghw6, Qfghw6, Xfghw6, Egghw6, Lgghw6, Sgghw6, Zgghw6, Ghghw6, Nhghw6, Uhghw6;
wire Bighw6, Iighw6, Pighw6, Wighw6, Djghw6, Kjghw6, Rjghw6, Yjghw6, Fkghw6, Mkghw6;
wire Tkghw6, Alghw6, Hlghw6, Olghw6, Vlghw6, Cmghw6, Jmghw6, Qmghw6, Xmghw6, Enghw6;
wire Lnghw6, Snghw6, Znghw6, Goghw6, Noghw6, Uoghw6, Bpghw6, Ipghw6, Ppghw6, Wpghw6;
wire Dqghw6, Kqghw6, Rqghw6, Yqghw6, Frghw6, Mrghw6, Trghw6, Asghw6, Hsghw6, Osghw6;
wire Vsghw6, Ctghw6, Jtghw6, Qtghw6, Xtghw6, Eughw6, Lughw6, Sughw6, Zughw6, Gvghw6;
wire Nvghw6, Uvghw6, Bwghw6, Iwghw6, Pwghw6, Wwghw6, Dxghw6, Kxghw6, Rxghw6, Yxghw6;
wire Fyghw6, Myghw6, Tyghw6, Azghw6, Hzghw6, Ozghw6, Vzghw6, C0hhw6, J0hhw6, Q0hhw6;
wire X0hhw6, E1hhw6, L1hhw6, S1hhw6, Z1hhw6, G2hhw6, N2hhw6, U2hhw6, B3hhw6, I3hhw6;
wire P3hhw6, W3hhw6, D4hhw6, K4hhw6, R4hhw6, Y4hhw6, F5hhw6, M5hhw6, T5hhw6, A6hhw6;
wire H6hhw6, O6hhw6, V6hhw6, C7hhw6, J7hhw6, Q7hhw6, X7hhw6, E8hhw6, L8hhw6, S8hhw6;
wire Z8hhw6, G9hhw6, N9hhw6, U9hhw6, Bahhw6, Iahhw6, Pahhw6, Wahhw6, Dbhhw6, Kbhhw6;
wire Rbhhw6, Ybhhw6, Fchhw6, Mchhw6, Tchhw6, Adhhw6, Hdhhw6, Odhhw6, Vdhhw6, Cehhw6;
wire Jehhw6, Qehhw6, Xehhw6, Efhhw6, Lfhhw6, Sfhhw6, Zfhhw6, Gghhw6, Nghhw6, Ughhw6;
wire Bhhhw6, Ihhhw6, Phhhw6, Whhhw6, Dihhw6, Kihhw6, Rihhw6, Yihhw6, Fjhhw6, Mjhhw6;
wire Tjhhw6, Akhhw6, Hkhhw6, Okhhw6, Vkhhw6, Clhhw6, Jlhhw6, Qlhhw6, Xlhhw6, Emhhw6;
wire Lmhhw6, Smhhw6, Zmhhw6, Gnhhw6, Nnhhw6, Unhhw6, Bohhw6, Iohhw6, Pohhw6, Wohhw6;
wire Dphhw6, Kphhw6, Rphhw6, Yphhw6, Fqhhw6, Mqhhw6, Tqhhw6, Arhhw6, Hrhhw6, Orhhw6;
wire Vrhhw6, Cshhw6, Jshhw6, Qshhw6, Xshhw6, Ethhw6, Lthhw6, Sthhw6, Zthhw6, Guhhw6;
wire Nuhhw6, Uuhhw6, Bvhhw6, Ivhhw6, Pvhhw6, Wvhhw6, Dwhhw6, Kwhhw6, Rwhhw6, Ywhhw6;
wire Fxhhw6, Mxhhw6, Txhhw6, Ayhhw6, Hyhhw6, Oyhhw6, Vyhhw6, Czhhw6, Jzhhw6, Qzhhw6;
wire Xzhhw6, E0ihw6, L0ihw6, S0ihw6, Z0ihw6, G1ihw6, N1ihw6, U1ihw6, B2ihw6, I2ihw6;
wire P2ihw6, W2ihw6, D3ihw6, K3ihw6, R3ihw6, Y3ihw6, F4ihw6, M4ihw6, T4ihw6, A5ihw6;
wire H5ihw6, O5ihw6, V5ihw6, C6ihw6, J6ihw6, Q6ihw6, X6ihw6, E7ihw6, L7ihw6, S7ihw6;
wire Z7ihw6, G8ihw6, N8ihw6, U8ihw6, B9ihw6, I9ihw6, P9ihw6, W9ihw6, Daihw6, Kaihw6;
wire Raihw6, Yaihw6, Fbihw6, Mbihw6, Tbihw6, Acihw6, Hcihw6, Ocihw6, Vcihw6, Cdihw6;
wire Jdihw6, Qdihw6, Xdihw6, Eeihw6, Leihw6, Seihw6, Zeihw6, Gfihw6, Nfihw6, Ufihw6;
wire Bgihw6, Igihw6, Pgihw6, Wgihw6, Dhihw6, Khihw6, Rhihw6, Yhihw6, Fiihw6, Miihw6;
wire Tiihw6, Ajihw6, Hjihw6, Ojihw6, Vjihw6, Ckihw6, Jkihw6, Qkihw6, Xkihw6, Elihw6;
wire Llihw6, Slihw6, Zlihw6, Gmihw6, Nmihw6, Umihw6, Bnihw6, Inihw6, Pnihw6, Wnihw6;
wire Doihw6, Koihw6, Roihw6, Yoihw6, Fpihw6, Mpihw6, Tpihw6, Aqihw6, Hqihw6, Oqihw6;
wire Vqihw6, Crihw6, Jrihw6, Qrihw6, Xrihw6, Esihw6, Lsihw6, Ssihw6, Zsihw6, Gtihw6;
wire Ntihw6, Utihw6, Buihw6, Iuihw6, Puihw6, Wuihw6, Dvihw6, Kvihw6, Rvihw6, Yvihw6;
wire Fwihw6, Mwihw6, Twihw6, Axihw6, Hxihw6, Oxihw6, Vxihw6, Cyihw6, Jyihw6, Qyihw6;
wire Xyihw6, Ezihw6, Lzihw6, Szihw6, Zzihw6, G0jhw6, N0jhw6, U0jhw6, B1jhw6, I1jhw6;
wire P1jhw6, W1jhw6, D2jhw6, K2jhw6, R2jhw6, Y2jhw6, F3jhw6, M3jhw6, T3jhw6, A4jhw6;
wire H4jhw6, O4jhw6, V4jhw6, C5jhw6, J5jhw6, Q5jhw6, X5jhw6, E6jhw6, L6jhw6, S6jhw6;
wire Z6jhw6, G7jhw6, N7jhw6, U7jhw6, B8jhw6, I8jhw6, P8jhw6, W8jhw6, D9jhw6, K9jhw6;
wire R9jhw6, Y9jhw6, Fajhw6, Majhw6, Tajhw6, Abjhw6, Hbjhw6, Objhw6, Vbjhw6, Ccjhw6;
wire Jcjhw6, Qcjhw6, Xcjhw6, Edjhw6, Ldjhw6, Sdjhw6, Zdjhw6, Gejhw6, Nejhw6, Uejhw6;
wire Bfjhw6, Ifjhw6, Pfjhw6, Wfjhw6, Dgjhw6, Kgjhw6, Rgjhw6, Ygjhw6, Fhjhw6, Mhjhw6;
wire Thjhw6, Aijhw6, Hijhw6, Oijhw6, Vijhw6, Cjjhw6, Jjjhw6, Qjjhw6, Xjjhw6, Ekjhw6;
wire Lkjhw6, Skjhw6, Zkjhw6, Gljhw6, Nljhw6, Uljhw6, Bmjhw6, Imjhw6, Pmjhw6, Wmjhw6;
wire Dnjhw6, Knjhw6, Rnjhw6, Ynjhw6, Fojhw6, Mojhw6, Tojhw6, Apjhw6, Hpjhw6, Opjhw6;
wire Vpjhw6, Cqjhw6, Jqjhw6, Qqjhw6, Xqjhw6, Erjhw6, Lrjhw6, Srjhw6, Zrjhw6, Gsjhw6;
wire Nsjhw6, Usjhw6, Btjhw6, Itjhw6, Ptjhw6, Wtjhw6, Dujhw6, Kujhw6, Rujhw6, Yujhw6;
wire Fvjhw6, Mvjhw6, Tvjhw6, Awjhw6, Hwjhw6, Owjhw6, Vwjhw6, Cxjhw6, Jxjhw6, Qxjhw6;
wire Xxjhw6, Eyjhw6, Lyjhw6, Syjhw6, Zyjhw6, Gzjhw6, Nzjhw6, Uzjhw6, B0khw6, I0khw6;
wire P0khw6, W0khw6, D1khw6, K1khw6, R1khw6, Y1khw6, F2khw6, M2khw6, T2khw6, A3khw6;
wire H3khw6, O3khw6, V3khw6, C4khw6, J4khw6, Q4khw6, X4khw6, E5khw6, L5khw6, S5khw6;
wire Z5khw6, G6khw6, N6khw6, U6khw6, B7khw6, I7khw6, P7khw6, W7khw6, D8khw6, K8khw6;
wire R8khw6, Y8khw6, F9khw6, M9khw6, T9khw6, Aakhw6, Hakhw6, Oakhw6, Vakhw6, Cbkhw6;
wire Jbkhw6, Qbkhw6, Xbkhw6, Eckhw6, Lckhw6, Sckhw6, Zckhw6, Gdkhw6, Ndkhw6, Udkhw6;
wire Bekhw6, Iekhw6, Pekhw6, Wekhw6, Dfkhw6, Kfkhw6, Rfkhw6, Yfkhw6, Fgkhw6, Mgkhw6;
wire Tgkhw6, Ahkhw6, Hhkhw6, Ohkhw6, Vhkhw6, Cikhw6, Jikhw6, Qikhw6, Xikhw6, Ejkhw6;
wire Ljkhw6, Sjkhw6, Zjkhw6, Gkkhw6, Nkkhw6, Ukkhw6, Blkhw6, Ilkhw6, Plkhw6, Wlkhw6;
wire Dmkhw6, Kmkhw6, Rmkhw6, Ymkhw6, Fnkhw6, Mnkhw6, Tnkhw6, Aokhw6, Hokhw6, Ookhw6;
wire Vokhw6, Cpkhw6, Jpkhw6, Qpkhw6, Xpkhw6, Eqkhw6, Lqkhw6, Sqkhw6, Zqkhw6, Grkhw6;
wire Nrkhw6, Urkhw6, Bskhw6, Iskhw6, Pskhw6, Wskhw6, Dtkhw6, Ktkhw6, Rtkhw6, Ytkhw6;
wire Fukhw6, Mukhw6, Tukhw6, Avkhw6, Hvkhw6, Ovkhw6, Vvkhw6, Cwkhw6, Jwkhw6, Qwkhw6;
wire Xwkhw6, Exkhw6, Lxkhw6, Sxkhw6, Zxkhw6, Gykhw6, Nykhw6, Uykhw6, Bzkhw6, Izkhw6;
wire Pzkhw6, Wzkhw6, D0lhw6, K0lhw6, R0lhw6, Y0lhw6, F1lhw6, M1lhw6, T1lhw6, A2lhw6;
wire H2lhw6, O2lhw6, V2lhw6, C3lhw6, J3lhw6, Q3lhw6, X3lhw6, E4lhw6, L4lhw6, S4lhw6;
wire Z4lhw6, G5lhw6, N5lhw6, U5lhw6, B6lhw6, I6lhw6, P6lhw6, W6lhw6, D7lhw6, K7lhw6;
wire R7lhw6, Y7lhw6, F8lhw6, M8lhw6, T8lhw6, A9lhw6, H9lhw6, O9lhw6, V9lhw6, Calhw6;
wire Jalhw6, Qalhw6, Xalhw6, Eblhw6, Lblhw6, Sblhw6, Zblhw6, Gclhw6, Nclhw6, Uclhw6;
wire Bdlhw6, Idlhw6, Pdlhw6, Wdlhw6, Delhw6, Kelhw6, Relhw6, Yelhw6, Fflhw6, Mflhw6;
wire Tflhw6, Aglhw6, Hglhw6, Oglhw6, Vglhw6, Chlhw6, Jhlhw6, Qhlhw6, Xhlhw6, Eilhw6;
wire Lilhw6, Silhw6, Zilhw6, Gjlhw6, Njlhw6, Ujlhw6, Bklhw6, Iklhw6, Pklhw6, Wklhw6;
wire Dllhw6, Kllhw6, Rllhw6, Yllhw6, Fmlhw6, Mmlhw6, Tmlhw6, Anlhw6, Hnlhw6, Onlhw6;
wire Vnlhw6, Colhw6, Jolhw6, Qolhw6, Xolhw6, Eplhw6, Lplhw6, Splhw6, Zplhw6, Gqlhw6;
wire Nqlhw6, Uqlhw6, Brlhw6, Irlhw6, Prlhw6, Wrlhw6, Dslhw6, Kslhw6, Rslhw6, Yslhw6;
wire Ftlhw6, Mtlhw6, Ttlhw6, Aulhw6, Hulhw6, Oulhw6, Vulhw6, Cvlhw6, Jvlhw6, Qvlhw6;
wire Xvlhw6, Ewlhw6, Lwlhw6, Swlhw6, Zwlhw6, Gxlhw6, Nxlhw6, Uxlhw6, Bylhw6, Iylhw6;
wire Pylhw6, Wylhw6, Dzlhw6, Kzlhw6, Rzlhw6, Yzlhw6, F0mhw6, M0mhw6, T0mhw6, A1mhw6;
wire H1mhw6, O1mhw6, V1mhw6, C2mhw6, J2mhw6, Q2mhw6, X2mhw6, E3mhw6, L3mhw6, S3mhw6;
wire Z3mhw6, G4mhw6, N4mhw6, U4mhw6, B5mhw6, I5mhw6, P5mhw6, W5mhw6, D6mhw6, K6mhw6;
wire R6mhw6, Y6mhw6, F7mhw6, M7mhw6, T7mhw6, A8mhw6, H8mhw6, O8mhw6, V8mhw6, C9mhw6;
wire J9mhw6, Q9mhw6, X9mhw6, Eamhw6, Lamhw6, Samhw6, Zamhw6, Gbmhw6, Nbmhw6, Ubmhw6;
wire Bcmhw6, Icmhw6, Pcmhw6, Wcmhw6, Ddmhw6, Kdmhw6, Rdmhw6, Ydmhw6, Femhw6, Memhw6;
wire Temhw6, Afmhw6, Hfmhw6, Ofmhw6, Vfmhw6, Cgmhw6, Jgmhw6, Qgmhw6, Xgmhw6, Ehmhw6;
wire Lhmhw6, Shmhw6, Zhmhw6, Gimhw6, Nimhw6, Uimhw6, Bjmhw6, Ijmhw6, Pjmhw6, Wjmhw6;
wire Dkmhw6, Kkmhw6, Rkmhw6, Ykmhw6, Flmhw6, Mlmhw6, Tlmhw6, Ammhw6, Hmmhw6, Ommhw6;
wire Vmmhw6, Cnmhw6, Jnmhw6, Qnmhw6, Xnmhw6, Eomhw6, Lomhw6, Somhw6, Zomhw6, Gpmhw6;
wire Npmhw6, Upmhw6, Bqmhw6, Iqmhw6, Pqmhw6, Wqmhw6, Drmhw6, Krmhw6, Rrmhw6, Yrmhw6;
wire Fsmhw6, Msmhw6, Tsmhw6, Atmhw6, Htmhw6, Otmhw6, Vtmhw6, Cumhw6, Jumhw6, Qumhw6;
wire Xumhw6, Evmhw6, Lvmhw6, Svmhw6, Zvmhw6, Gwmhw6, Nwmhw6, Uwmhw6, Bxmhw6, Ixmhw6;
wire Pxmhw6, Wxmhw6, Dymhw6, Kymhw6, Rymhw6, Yymhw6, Fzmhw6, Mzmhw6, Tzmhw6, A0nhw6;
wire H0nhw6, O0nhw6, V0nhw6, C1nhw6, J1nhw6, Q1nhw6, X1nhw6, E2nhw6, L2nhw6, S2nhw6;
wire Z2nhw6, G3nhw6, N3nhw6, U3nhw6, B4nhw6, I4nhw6, P4nhw6, W4nhw6, D5nhw6, K5nhw6;
wire R5nhw6, Y5nhw6, F6nhw6, M6nhw6, T6nhw6, A7nhw6, H7nhw6, O7nhw6, V7nhw6, C8nhw6;
wire J8nhw6, Q8nhw6, X8nhw6, E9nhw6, L9nhw6, S9nhw6, Z9nhw6, Ganhw6, Nanhw6, Uanhw6;
wire Bbnhw6, Ibnhw6, Pbnhw6, Wbnhw6, Dcnhw6, Kcnhw6, Rcnhw6, Ycnhw6, Fdnhw6, Mdnhw6;
wire Tdnhw6, Aenhw6, Henhw6, Oenhw6, Venhw6, Cfnhw6, Jfnhw6, Qfnhw6, Xfnhw6, Egnhw6;
wire Lgnhw6, Sgnhw6, Zgnhw6, Ghnhw6, Nhnhw6, Uhnhw6, Binhw6, Iinhw6, Pinhw6, Winhw6;
wire Djnhw6, Kjnhw6, Rjnhw6, Yjnhw6, Fknhw6, Mknhw6, Tknhw6, Alnhw6, Hlnhw6, Olnhw6;
wire Vlnhw6, Cmnhw6, Jmnhw6, Qmnhw6, Xmnhw6, Ennhw6, Lnnhw6, Snnhw6, Znnhw6, Gonhw6;
wire Nonhw6, Uonhw6, Bpnhw6, Ipnhw6, Ppnhw6, Wpnhw6, Dqnhw6, Kqnhw6, Rqnhw6, Yqnhw6;
wire Frnhw6, Mrnhw6, Trnhw6, Asnhw6, Hsnhw6, Osnhw6, Vsnhw6, Ctnhw6, Jtnhw6, Qtnhw6;
wire Xtnhw6, Eunhw6, Lunhw6, Sunhw6, Zunhw6, Gvnhw6, Nvnhw6, Uvnhw6, Bwnhw6, Iwnhw6;
wire Pwnhw6, Wwnhw6, Dxnhw6, Kxnhw6, Rxnhw6, Yxnhw6, Fynhw6, Mynhw6, Tynhw6, Aznhw6;
wire Hznhw6, Oznhw6, Vznhw6, C0ohw6, J0ohw6, Q0ohw6, X0ohw6, E1ohw6, L1ohw6, S1ohw6;
wire Z1ohw6, G2ohw6, N2ohw6, U2ohw6, B3ohw6, I3ohw6, P3ohw6, W3ohw6, D4ohw6, K4ohw6;
wire R4ohw6, Y4ohw6, F5ohw6, M5ohw6, T5ohw6, A6ohw6, H6ohw6, O6ohw6, V6ohw6, C7ohw6;
wire J7ohw6, Q7ohw6, X7ohw6, E8ohw6, L8ohw6, S8ohw6, Z8ohw6, G9ohw6, N9ohw6, U9ohw6;
wire Baohw6, Iaohw6, Paohw6, Waohw6, Dbohw6, Kbohw6, Rbohw6, Ybohw6, Fcohw6, Mcohw6;
wire Tcohw6, Adohw6, Hdohw6, Odohw6, Vdohw6, Ceohw6, Jeohw6, Qeohw6, Xeohw6, Efohw6;
wire Lfohw6, Sfohw6, Zfohw6, Ggohw6, Ngohw6, Ugohw6, Bhohw6, Ihohw6, Phohw6, Whohw6;
wire Diohw6, Kiohw6, Riohw6, Yiohw6, Fjohw6, Mjohw6, Tjohw6, Akohw6, Hkohw6, Okohw6;
wire Vkohw6, Clohw6, Jlohw6, Qlohw6, Xlohw6, Emohw6, Lmohw6, Smohw6, Zmohw6, Gnohw6;
wire Nnohw6, Unohw6, Boohw6, Ioohw6, Poohw6, Woohw6, Dpohw6, Kpohw6, Rpohw6, Ypohw6;
wire Fqohw6, Mqohw6, Tqohw6, Arohw6, Hrohw6, Orohw6, Vrohw6, Csohw6, Jsohw6, Qsohw6;
wire Xsohw6, Etohw6, Ltohw6, Stohw6, Ztohw6, Guohw6, Nuohw6, Uuohw6, Bvohw6, Ivohw6;
wire Pvohw6, Wvohw6, Dwohw6, Kwohw6, Rwohw6, Ywohw6, Fxohw6, Mxohw6, Txohw6, Ayohw6;
wire Hyohw6, Oyohw6, Vyohw6, Czohw6, Jzohw6, Qzohw6, Xzohw6, E0phw6, L0phw6, S0phw6;
wire Z0phw6, G1phw6, N1phw6, U1phw6, B2phw6, I2phw6, P2phw6, W2phw6, D3phw6, K3phw6;
wire R3phw6, Y3phw6, F4phw6, M4phw6, T4phw6, A5phw6, H5phw6, O5phw6, V5phw6, C6phw6;
wire J6phw6, Q6phw6, X6phw6, E7phw6, L7phw6, S7phw6, Z7phw6, G8phw6, N8phw6, U8phw6;
wire B9phw6, I9phw6, P9phw6, W9phw6, Daphw6, Kaphw6, Raphw6, Yaphw6, Fbphw6, Mbphw6;
wire Tbphw6, Acphw6, Hcphw6, Ocphw6, Vcphw6, Cdphw6, Jdphw6, Qdphw6, Xdphw6, Eephw6;
wire Lephw6, Sephw6, Zephw6, Gfphw6, Nfphw6, Ufphw6, Bgphw6, Igphw6, Pgphw6, Wgphw6;
wire Dhphw6, Khphw6, Rhphw6, Yhphw6, Fiphw6, Miphw6, Tiphw6, Ajphw6, Hjphw6, Ojphw6;
wire Vjphw6, Ckphw6, Jkphw6, Qkphw6, Xkphw6, Elphw6, Llphw6, Slphw6, Zlphw6, Gmphw6;
wire Nmphw6, Umphw6, Bnphw6, Inphw6, Pnphw6, Wnphw6, Dophw6, Kophw6, Rophw6, Yophw6;
wire Fpphw6, Mpphw6, Tpphw6, Aqphw6, Hqphw6, Oqphw6, Vqphw6, Crphw6, Jrphw6, Qrphw6;
wire Xrphw6, Esphw6, Lsphw6, Ssphw6, Zsphw6, Gtphw6, Ntphw6, Utphw6, Buphw6, Iuphw6;
wire Puphw6, Wuphw6, Dvphw6, Kvphw6, Rvphw6, Yvphw6, Fwphw6, Mwphw6, Twphw6, Axphw6;
wire Hxphw6, Oxphw6, Vxphw6, Cyphw6, Jyphw6, Qyphw6, Xyphw6, Ezphw6, Lzphw6, Szphw6;
wire Zzphw6, G0qhw6, N0qhw6, U0qhw6, B1qhw6, I1qhw6, P1qhw6, W1qhw6, D2qhw6, K2qhw6;
wire R2qhw6, Y2qhw6, F3qhw6, M3qhw6, T3qhw6, A4qhw6, H4qhw6, O4qhw6, V4qhw6, C5qhw6;
wire J5qhw6, Q5qhw6, X5qhw6, E6qhw6, L6qhw6, S6qhw6, Z6qhw6, G7qhw6, N7qhw6, U7qhw6;
wire B8qhw6, I8qhw6, P8qhw6, W8qhw6, D9qhw6, K9qhw6, R9qhw6, Y9qhw6, Faqhw6, Maqhw6;
wire Taqhw6, Abqhw6, Hbqhw6, Obqhw6, Vbqhw6, Ccqhw6, Jcqhw6, Qcqhw6, Xcqhw6, Edqhw6;
wire Ldqhw6, Sdqhw6, Zdqhw6, Geqhw6, Neqhw6, Ueqhw6, Bfqhw6, Ifqhw6, Pfqhw6, Wfqhw6;
wire Dgqhw6, Kgqhw6, Rgqhw6, Ygqhw6, Fhqhw6, Mhqhw6, Thqhw6, Aiqhw6, Hiqhw6, Oiqhw6;
wire Viqhw6, Cjqhw6, Jjqhw6, Qjqhw6, Xjqhw6, Ekqhw6, Lkqhw6, Skqhw6, Zkqhw6, Glqhw6;
wire Nlqhw6, Ulqhw6, Bmqhw6, Imqhw6, Pmqhw6, Wmqhw6, Dnqhw6, Knqhw6, Rnqhw6, Ynqhw6;
wire Foqhw6, Moqhw6, Toqhw6, Apqhw6, Hpqhw6, Opqhw6, Vpqhw6, Cqqhw6, Jqqhw6, Qqqhw6;
wire Xqqhw6, Erqhw6, Lrqhw6, Srqhw6, Zrqhw6, Gsqhw6, Nsqhw6, Usqhw6, Btqhw6, Itqhw6;
wire Ptqhw6, Wtqhw6, Duqhw6, Kuqhw6, Ruqhw6, Yuqhw6, Fvqhw6, Mvqhw6, Tvqhw6, Awqhw6;
wire Hwqhw6, Owqhw6, Vwqhw6, Cxqhw6, Jxqhw6, Qxqhw6, Xxqhw6, Eyqhw6, Lyqhw6, Syqhw6;
wire Zyqhw6, Gzqhw6, Nzqhw6, Uzqhw6, B0rhw6, I0rhw6, P0rhw6, W0rhw6, D1rhw6, K1rhw6;
wire R1rhw6, Y1rhw6, F2rhw6, M2rhw6, T2rhw6, A3rhw6, H3rhw6, O3rhw6, V3rhw6, C4rhw6;
wire J4rhw6, Q4rhw6, X4rhw6, E5rhw6, L5rhw6, S5rhw6, Z5rhw6, G6rhw6, N6rhw6, U6rhw6;
wire B7rhw6, I7rhw6, P7rhw6, W7rhw6, D8rhw6, K8rhw6, R8rhw6, Y8rhw6, F9rhw6, M9rhw6;
wire T9rhw6, Aarhw6, Harhw6, Oarhw6, Varhw6, Cbrhw6, Jbrhw6, Qbrhw6, Xbrhw6, Ecrhw6;
wire Lcrhw6, Scrhw6, Zcrhw6, Gdrhw6, Ndrhw6, Udrhw6, Berhw6, Ierhw6, Perhw6, Werhw6;
wire Dfrhw6, Kfrhw6, Rfrhw6, Yfrhw6, Fgrhw6, Mgrhw6, Tgrhw6, Ahrhw6, Hhrhw6, Ohrhw6;
wire Vhrhw6, Cirhw6, Jirhw6, Qirhw6, Xirhw6, Ejrhw6, Ljrhw6, Sjrhw6, Zjrhw6, Gkrhw6;
wire Nkrhw6, Ukrhw6, Blrhw6, Ilrhw6, Plrhw6, Wlrhw6, Dmrhw6, Kmrhw6, Rmrhw6, Ymrhw6;
wire Fnrhw6, Mnrhw6, Tnrhw6, Aorhw6, Horhw6, Oorhw6, Vorhw6, Cprhw6, Jprhw6, Qprhw6;
wire Xprhw6, Eqrhw6, Lqrhw6, Sqrhw6, Zqrhw6, Grrhw6, Nrrhw6, Urrhw6, Bsrhw6, Isrhw6;
wire Psrhw6, Wsrhw6, Dtrhw6, Ktrhw6, Rtrhw6, Ytrhw6, Furhw6, Murhw6, Turhw6, Avrhw6;
wire Hvrhw6, Ovrhw6, Vvrhw6, Cwrhw6, Jwrhw6, Qwrhw6, Xwrhw6, Exrhw6, Lxrhw6, Sxrhw6;
wire Zxrhw6, Gyrhw6, Nyrhw6, Uyrhw6, Bzrhw6, Izrhw6, Pzrhw6, Wzrhw6, D0shw6, K0shw6;
wire R0shw6, Y0shw6, F1shw6, M1shw6, T1shw6, A2shw6, H2shw6, O2shw6, V2shw6, C3shw6;
wire J3shw6, Q3shw6, X3shw6, E4shw6, L4shw6, S4shw6, Z4shw6, G5shw6, N5shw6, U5shw6;
wire B6shw6, I6shw6, P6shw6, W6shw6, D7shw6, K7shw6, R7shw6, Y7shw6, F8shw6, M8shw6;
wire T8shw6, A9shw6, H9shw6, O9shw6, V9shw6, Cashw6, Jashw6, Qashw6, Xashw6, Ebshw6;
wire Lbshw6, Sbshw6, Zbshw6, Gcshw6, Ncshw6, Ucshw6, Bdshw6, Idshw6, Pdshw6, Wdshw6;
wire Deshw6, Keshw6, Reshw6, Yeshw6, Ffshw6, Mfshw6, Tfshw6, Agshw6, Hgshw6, Ogshw6;
wire Vgshw6, Chshw6, Jhshw6, Qhshw6, Xhshw6, Eishw6, Lishw6, Sishw6, Zishw6, Gjshw6;
wire Njshw6, Ujshw6, Bkshw6, Ikshw6, Pkshw6, Wkshw6, Dlshw6, Klshw6, Rlshw6, Ylshw6;
wire Fmshw6, Mmshw6, Tmshw6, Anshw6, Hnshw6, Onshw6, Vnshw6, Coshw6, Joshw6, Qoshw6;
wire Xoshw6, Epshw6, Lpshw6, Spshw6, Zpshw6, Gqshw6, Nqshw6, Uqshw6, Brshw6, Irshw6;
wire Prshw6, Wrshw6, Dsshw6, Ksshw6, Rsshw6, Ysshw6, Ftshw6, Mtshw6, Ttshw6, Aushw6;
wire Hushw6, Oushw6, Vushw6, Cvshw6, Jvshw6, Qvshw6, Xvshw6, Ewshw6, Lwshw6, Swshw6;
wire Zwshw6, Gxshw6, Nxshw6, Uxshw6, Byshw6, Iyshw6, Pyshw6, Wyshw6, Dzshw6, Kzshw6;
wire Rzshw6, Yzshw6, F0thw6, M0thw6, T0thw6, A1thw6, H1thw6, O1thw6, V1thw6, C2thw6;
wire J2thw6, Q2thw6, X2thw6, E3thw6, L3thw6, S3thw6, Z3thw6, G4thw6, N4thw6, U4thw6;
wire B5thw6, I5thw6, P5thw6, W5thw6, D6thw6, K6thw6, R6thw6, Y6thw6, F7thw6, M7thw6;
wire T7thw6, A8thw6, H8thw6, O8thw6, V8thw6, C9thw6, J9thw6, Q9thw6, X9thw6, Eathw6;
wire Lathw6, Sathw6, Zathw6, Gbthw6, Nbthw6, Ubthw6, Bcthw6, Icthw6, Pcthw6, Wcthw6;
wire Ddthw6, Kdthw6, Rdthw6, Ydthw6, Fethw6, Methw6, Tethw6, Afthw6, Hfthw6, Ofthw6;
wire Vfthw6, Cgthw6, Jgthw6, Qgthw6, Xgthw6, Ehthw6, Lhthw6, Shthw6, Zhthw6, Githw6;
wire Nithw6, Uithw6, Bjthw6, Ijthw6, Pjthw6, Wjthw6, Dkthw6, Kkthw6, Rkthw6, Ykthw6;
wire Flthw6, Mlthw6, Tlthw6, Amthw6, Hmthw6, Omthw6, Vmthw6, Cnthw6, Jnthw6, Qnthw6;
wire Xnthw6, Eothw6, Lothw6, Sothw6, Zothw6, Gpthw6, Npthw6, Upthw6, Bqthw6, Iqthw6;
wire Pqthw6, Wqthw6, Drthw6, Krthw6, Rrthw6, Yrthw6, Fsthw6, Msthw6, Tsthw6, Atthw6;
wire Htthw6, Otthw6, Vtthw6, Cuthw6, Juthw6, Quthw6, Xuthw6, Evthw6, Lvthw6, Svthw6;
wire Zvthw6, Gwthw6, Nwthw6, Uwthw6, Bxthw6, Ixthw6, Pxthw6, Wxthw6, Dythw6, Kythw6;
wire Rythw6, Yythw6, Fzthw6, Mzthw6, Tzthw6, A0uhw6, H0uhw6, O0uhw6, V0uhw6, C1uhw6;
wire J1uhw6, Q1uhw6, X1uhw6, E2uhw6, L2uhw6, S2uhw6, Z2uhw6, G3uhw6, N3uhw6, U3uhw6;
wire B4uhw6, I4uhw6, P4uhw6, W4uhw6, D5uhw6, K5uhw6, R5uhw6, Y5uhw6, F6uhw6, M6uhw6;
wire T6uhw6, A7uhw6, H7uhw6, O7uhw6, V7uhw6, C8uhw6, J8uhw6, Q8uhw6, X8uhw6, E9uhw6;
wire L9uhw6, S9uhw6, Z9uhw6, Gauhw6, Nauhw6, Uauhw6, Bbuhw6, Ibuhw6, Pbuhw6, Wbuhw6;
wire Dcuhw6, Kcuhw6, Rcuhw6, Ycuhw6, Fduhw6, Mduhw6, Tduhw6, Aeuhw6, Heuhw6, Oeuhw6;
wire Veuhw6, Cfuhw6, Jfuhw6, Qfuhw6, Xfuhw6, Eguhw6, Lguhw6, Sguhw6, Zguhw6, Ghuhw6;
wire Nhuhw6, Uhuhw6, Biuhw6, Iiuhw6, Piuhw6, Wiuhw6, Djuhw6, Kjuhw6, Rjuhw6, Yjuhw6;
wire Fkuhw6, Mkuhw6, Tkuhw6, Aluhw6, Hluhw6, Oluhw6, Vluhw6, Cmuhw6, Jmuhw6, Qmuhw6;
wire Xmuhw6, Enuhw6, Lnuhw6, Snuhw6, Znuhw6, Gouhw6, Nouhw6, Uouhw6, Bpuhw6, Ipuhw6;
wire Ppuhw6, Wpuhw6, Dquhw6, Kquhw6, Rquhw6, Yquhw6, Fruhw6, Mruhw6, Truhw6, Asuhw6;
wire Hsuhw6, Osuhw6, Vsuhw6, Ctuhw6, Jtuhw6, Qtuhw6, Xtuhw6, Euuhw6, Luuhw6, Suuhw6;
wire Zuuhw6, Gvuhw6, Nvuhw6, Uvuhw6, Bwuhw6, Iwuhw6, Pwuhw6, Wwuhw6, Dxuhw6, Kxuhw6;
wire Rxuhw6, Yxuhw6, Fyuhw6, Myuhw6, Tyuhw6, Azuhw6, Hzuhw6, Ozuhw6, Vzuhw6, C0vhw6;
wire J0vhw6, Q0vhw6, X0vhw6, E1vhw6, L1vhw6, S1vhw6, Z1vhw6, G2vhw6, N2vhw6, U2vhw6;
wire B3vhw6, I3vhw6, P3vhw6, W3vhw6, D4vhw6, K4vhw6, R4vhw6, Y4vhw6, F5vhw6, M5vhw6;
wire T5vhw6, A6vhw6, H6vhw6, O6vhw6, V6vhw6, C7vhw6, J7vhw6, Q7vhw6, X7vhw6, E8vhw6;
wire L8vhw6, S8vhw6, Z8vhw6, G9vhw6, N9vhw6, U9vhw6, Bavhw6, Iavhw6, Pavhw6, Wavhw6;
wire Dbvhw6, Kbvhw6, Rbvhw6, Ybvhw6, Fcvhw6, Mcvhw6, Tcvhw6, Advhw6, Hdvhw6, Odvhw6;
wire Vdvhw6, Cevhw6, Jevhw6, Qevhw6, Xevhw6, Efvhw6, Lfvhw6, Sfvhw6, Zfvhw6, Ggvhw6;
wire Ngvhw6, Ugvhw6, Bhvhw6, Ihvhw6, Phvhw6, Whvhw6, Divhw6, Kivhw6, Rivhw6, Yivhw6;
wire Fjvhw6, Mjvhw6, Tjvhw6, Akvhw6, Hkvhw6, Okvhw6, Vkvhw6, Clvhw6, Jlvhw6, Qlvhw6;
wire Xlvhw6, Emvhw6, Lmvhw6, Smvhw6, Zmvhw6, Gnvhw6, Nnvhw6, Unvhw6, Bovhw6, Iovhw6;
wire Povhw6, Wovhw6, Dpvhw6, Kpvhw6, Rpvhw6, Ypvhw6, Fqvhw6, Mqvhw6, Tqvhw6, Arvhw6;
wire Hrvhw6, Orvhw6, Vrvhw6, Csvhw6, Jsvhw6, Qsvhw6, Xsvhw6, Etvhw6, Ltvhw6, Stvhw6;
wire Ztvhw6, Guvhw6, Nuvhw6, Uuvhw6, Bvvhw6, Ivvhw6, Pvvhw6, Wvvhw6, Dwvhw6, Kwvhw6;
wire Rwvhw6, Ywvhw6, Fxvhw6, Mxvhw6, Txvhw6, Ayvhw6, Hyvhw6, Oyvhw6, Vyvhw6, Czvhw6;
wire Jzvhw6, Qzvhw6, Xzvhw6, E0whw6, L0whw6, S0whw6, Z0whw6, G1whw6, N1whw6, U1whw6;
wire B2whw6, I2whw6, P2whw6, W2whw6, D3whw6, K3whw6, R3whw6, Y3whw6, F4whw6, M4whw6;
wire T4whw6, A5whw6, H5whw6, O5whw6, V5whw6, C6whw6, J6whw6, Q6whw6, X6whw6, E7whw6;
wire L7whw6, S7whw6, Z7whw6, G8whw6, N8whw6, U8whw6, B9whw6, I9whw6, P9whw6, W9whw6;
wire Dawhw6, Kawhw6, Rawhw6, Yawhw6, Fbwhw6, Mbwhw6, Tbwhw6, Acwhw6, Hcwhw6, Ocwhw6;
wire Vcwhw6, Cdwhw6, Jdwhw6, Qdwhw6, Xdwhw6, Eewhw6, Lewhw6, Sewhw6, Zewhw6, Gfwhw6;
wire Nfwhw6, Ufwhw6, Bgwhw6, Igwhw6, Pgwhw6, Wgwhw6, Dhwhw6, Khwhw6, Rhwhw6, Yhwhw6;
wire Fiwhw6, Miwhw6, Tiwhw6, Ajwhw6, Hjwhw6, Ojwhw6, Vjwhw6, Ckwhw6, Jkwhw6, Qkwhw6;
wire Xkwhw6, Elwhw6, Llwhw6, Slwhw6, Zlwhw6, Gmwhw6, Nmwhw6, Umwhw6, Bnwhw6, Inwhw6;
wire Pnwhw6, Wnwhw6, Dowhw6, Kowhw6, Rowhw6, Yowhw6, Fpwhw6, Mpwhw6, Tpwhw6, Aqwhw6;
wire Hqwhw6, Oqwhw6, Vqwhw6, Crwhw6, Jrwhw6, Qrwhw6, Xrwhw6, Eswhw6, Lswhw6, Sswhw6;
wire Zswhw6, Gtwhw6, Ntwhw6, Utwhw6, Buwhw6, Iuwhw6, Puwhw6, Wuwhw6, Dvwhw6, Kvwhw6;
wire Rvwhw6, Yvwhw6, Fwwhw6, Mwwhw6, Twwhw6, Axwhw6, Hxwhw6, Oxwhw6, Vxwhw6, Cywhw6;
wire Jywhw6, Qywhw6, Xywhw6, Ezwhw6, Lzwhw6, Szwhw6, Zzwhw6, G0xhw6, N0xhw6, U0xhw6;
wire B1xhw6, I1xhw6, P1xhw6, W1xhw6, D2xhw6, K2xhw6, R2xhw6, Y2xhw6, F3xhw6, M3xhw6;
wire T3xhw6, A4xhw6, H4xhw6, O4xhw6, V4xhw6, C5xhw6, J5xhw6, Q5xhw6, X5xhw6, E6xhw6;
wire L6xhw6, S6xhw6, Z6xhw6, G7xhw6, N7xhw6, U7xhw6, B8xhw6, I8xhw6, P8xhw6, W8xhw6;
wire D9xhw6, K9xhw6, R9xhw6, Y9xhw6, Faxhw6, Maxhw6, Taxhw6, Abxhw6, Hbxhw6, Obxhw6;
wire Vbxhw6, Ccxhw6, Jcxhw6, Qcxhw6, Xcxhw6, Edxhw6, Ldxhw6, Sdxhw6, Zdxhw6, Gexhw6;
wire Nexhw6, Uexhw6, Bfxhw6, Ifxhw6, Pfxhw6, Wfxhw6, Dgxhw6, Kgxhw6, Rgxhw6, Ygxhw6;
wire Fhxhw6, Mhxhw6, Thxhw6, Aixhw6, Hixhw6, Oixhw6, Vixhw6, Cjxhw6, Jjxhw6, Qjxhw6;
wire Xjxhw6, Ekxhw6, Lkxhw6, Skxhw6, Zkxhw6, Glxhw6, Nlxhw6, Ulxhw6, Bmxhw6, Imxhw6;
wire Pmxhw6, Wmxhw6, Dnxhw6, Knxhw6, Rnxhw6, Ynxhw6, Foxhw6, Moxhw6, Toxhw6, Apxhw6;
wire Hpxhw6, Opxhw6, Vpxhw6, Cqxhw6, Jqxhw6, Qqxhw6, Xqxhw6, Erxhw6, Lrxhw6, Srxhw6;
wire Zrxhw6, Gsxhw6, Nsxhw6, Usxhw6, Btxhw6, Itxhw6, Ptxhw6, Wtxhw6, Duxhw6, Kuxhw6;
wire Ruxhw6, Yuxhw6, Fvxhw6, Mvxhw6, Tvxhw6, Awxhw6, Hwxhw6, Owxhw6, Vwxhw6, Cxxhw6;
wire Jxxhw6, Qxxhw6, Xxxhw6, Eyxhw6, Lyxhw6, Syxhw6, Zyxhw6, Gzxhw6, Nzxhw6, Uzxhw6;
wire B0yhw6, I0yhw6, P0yhw6, W0yhw6, D1yhw6, K1yhw6, R1yhw6, Y1yhw6, F2yhw6, M2yhw6;
wire T2yhw6, A3yhw6, H3yhw6, O3yhw6, V3yhw6, C4yhw6, J4yhw6, Q4yhw6, X4yhw6, E5yhw6;
wire L5yhw6, S5yhw6, Z5yhw6, G6yhw6, N6yhw6, U6yhw6, B7yhw6, I7yhw6, P7yhw6, W7yhw6;
wire D8yhw6, K8yhw6, R8yhw6, Y8yhw6, F9yhw6, M9yhw6, T9yhw6, Aayhw6, Hayhw6, Oayhw6;
wire Vayhw6, Cbyhw6, Jbyhw6, Qbyhw6, Xbyhw6, Ecyhw6, Lcyhw6, Scyhw6, Zcyhw6, Gdyhw6;
wire Ndyhw6, Udyhw6, Beyhw6, Ieyhw6, Peyhw6, Weyhw6, Dfyhw6, Kfyhw6, Rfyhw6, Yfyhw6;
wire Fgyhw6, Mgyhw6, Tgyhw6, Ahyhw6, Hhyhw6, Ohyhw6, Vhyhw6, Ciyhw6, Jiyhw6, Qiyhw6;
wire Xiyhw6, Ejyhw6, Ljyhw6, Sjyhw6, Zjyhw6, Gkyhw6, Nkyhw6, Ukyhw6, Blyhw6, Ilyhw6;
wire Plyhw6, Wlyhw6, Dmyhw6, Kmyhw6, Rmyhw6, Ymyhw6, Fnyhw6, Mnyhw6, Tnyhw6, Aoyhw6;
wire Hoyhw6, Ooyhw6, Voyhw6, Cpyhw6, Jpyhw6, Qpyhw6, Xpyhw6, Eqyhw6, Lqyhw6, Sqyhw6;
wire Zqyhw6, Gryhw6, Nryhw6, Uryhw6, Bsyhw6, Isyhw6, Psyhw6, Wsyhw6, Dtyhw6, Ktyhw6;
wire Rtyhw6, Ytyhw6, Fuyhw6, Muyhw6, Tuyhw6, Avyhw6, Hvyhw6, Ovyhw6, Vvyhw6, Cwyhw6;
wire Jwyhw6, Qwyhw6, Xwyhw6, Exyhw6, Lxyhw6, Sxyhw6, Zxyhw6, Gyyhw6, Nyyhw6, Uyyhw6;
wire Bzyhw6, Izyhw6, Pzyhw6, Wzyhw6, D0zhw6, K0zhw6, R0zhw6, Y0zhw6, F1zhw6, M1zhw6;
wire T1zhw6, A2zhw6, H2zhw6, O2zhw6, V2zhw6, C3zhw6, J3zhw6, Q3zhw6, X3zhw6, E4zhw6;
wire L4zhw6, S4zhw6, Z4zhw6, G5zhw6, N5zhw6, U5zhw6, B6zhw6, I6zhw6, P6zhw6, W6zhw6;
wire D7zhw6, K7zhw6, R7zhw6, Y7zhw6, F8zhw6, M8zhw6, T8zhw6, A9zhw6, H9zhw6, O9zhw6;
wire V9zhw6, Cazhw6, Jazhw6, Qazhw6, Xazhw6, Ebzhw6, Lbzhw6, Sbzhw6, Zbzhw6, Gczhw6;
wire Nczhw6, Uczhw6, Bdzhw6, Idzhw6, Pdzhw6, Wdzhw6, Dezhw6, Kezhw6, Rezhw6, Yezhw6;
wire Ffzhw6, Mfzhw6, Tfzhw6, Agzhw6, Hgzhw6, Ogzhw6, Vgzhw6, Chzhw6, Jhzhw6, Qhzhw6;
wire Xhzhw6, Eizhw6, Lizhw6, Sizhw6, Zizhw6, Gjzhw6, Njzhw6, Ujzhw6, Bkzhw6, Ikzhw6;
wire Pkzhw6, Wkzhw6, Dlzhw6, Klzhw6, Rlzhw6, Ylzhw6, Fmzhw6, Mmzhw6, Tmzhw6, Anzhw6;
wire Hnzhw6, Onzhw6, Vnzhw6, Cozhw6, Jozhw6, Qozhw6, Xozhw6, Epzhw6, Lpzhw6, Spzhw6;
wire Zpzhw6, Gqzhw6, Nqzhw6, Uqzhw6, Brzhw6, Irzhw6, Przhw6, Wrzhw6, Dszhw6, Kszhw6;
wire Rszhw6, Yszhw6, Ftzhw6, Mtzhw6, Ttzhw6, Auzhw6, Huzhw6, Ouzhw6, Vuzhw6, Cvzhw6;
wire Jvzhw6, Qvzhw6, Xvzhw6, Ewzhw6, Lwzhw6, Swzhw6, Zwzhw6, Gxzhw6, Nxzhw6, Uxzhw6;
wire Byzhw6, Iyzhw6, Pyzhw6, Wyzhw6, Dzzhw6, Kzzhw6, Rzzhw6, Yzzhw6, F00iw6, M00iw6;
wire T00iw6, A10iw6, H10iw6, O10iw6, V10iw6, C20iw6, J20iw6, Q20iw6, X20iw6, E30iw6;
wire L30iw6, S30iw6, Z30iw6, G40iw6, N40iw6, U40iw6, B50iw6, I50iw6, P50iw6, W50iw6;
wire D60iw6, K60iw6, R60iw6, Y60iw6, F70iw6, M70iw6, T70iw6, A80iw6, H80iw6, O80iw6;
wire V80iw6, C90iw6, J90iw6, Q90iw6, X90iw6, Ea0iw6, La0iw6, Sa0iw6, Za0iw6, Gb0iw6;
wire Nb0iw6, Ub0iw6, Bc0iw6, Ic0iw6, Pc0iw6, Wc0iw6, Dd0iw6, Kd0iw6, Rd0iw6, Yd0iw6;
wire Fe0iw6, Me0iw6, Te0iw6, Af0iw6, Hf0iw6, Of0iw6, Vf0iw6, Cg0iw6, Jg0iw6, Qg0iw6;
wire Xg0iw6, Eh0iw6, Lh0iw6, Sh0iw6, Zh0iw6, Gi0iw6, Ni0iw6, Ui0iw6, Bj0iw6, Ij0iw6;
wire Pj0iw6, Wj0iw6, Dk0iw6, Kk0iw6, Rk0iw6, Yk0iw6, Fl0iw6, Ml0iw6, Tl0iw6, Am0iw6;
wire Hm0iw6, Om0iw6, Vm0iw6, Cn0iw6, Jn0iw6, Qn0iw6, Xn0iw6, Eo0iw6, Lo0iw6, So0iw6;
wire Zo0iw6, Gp0iw6, Np0iw6, Up0iw6, Bq0iw6, Iq0iw6, Pq0iw6, Wq0iw6, Dr0iw6, Kr0iw6;
wire Rr0iw6, Yr0iw6, Fs0iw6, Ms0iw6, Ts0iw6, At0iw6, Ht0iw6, Ot0iw6, Vt0iw6, Cu0iw6;
wire Ju0iw6, Qu0iw6, Xu0iw6, Ev0iw6, Lv0iw6, Sv0iw6, Zv0iw6, Gw0iw6, Nw0iw6, Uw0iw6;
wire Bx0iw6, Ix0iw6, Px0iw6, Wx0iw6, Dy0iw6, Ky0iw6, Ry0iw6, Yy0iw6, Fz0iw6, Mz0iw6;
wire Tz0iw6, A01iw6, H01iw6, O01iw6, V01iw6, C11iw6, J11iw6, Q11iw6, X11iw6, E21iw6;
wire L21iw6, S21iw6, Z21iw6, G31iw6, N31iw6, U31iw6, B41iw6, I41iw6, P41iw6, W41iw6;
wire D51iw6, K51iw6, R51iw6, Y51iw6, F61iw6, M61iw6, T61iw6, A71iw6, H71iw6, O71iw6;
wire V71iw6, C81iw6, J81iw6, Q81iw6, X81iw6, E91iw6, L91iw6, S91iw6, Z91iw6, Ga1iw6;
wire Na1iw6, Ua1iw6, Bb1iw6, Ib1iw6, Pb1iw6, Wb1iw6, Dc1iw6, Kc1iw6, Rc1iw6, Yc1iw6;
wire Fd1iw6, Md1iw6, Td1iw6, Ae1iw6, He1iw6, Oe1iw6, Ve1iw6, Cf1iw6, Jf1iw6, Qf1iw6;
wire Xf1iw6, Eg1iw6, Lg1iw6, Sg1iw6, Zg1iw6, Gh1iw6, Nh1iw6, Uh1iw6, Bi1iw6, Ii1iw6;
wire Pi1iw6, Wi1iw6, Dj1iw6, Kj1iw6, Rj1iw6, Yj1iw6, Fk1iw6, Mk1iw6, Tk1iw6, Al1iw6;
wire Hl1iw6, Ol1iw6, Vl1iw6, Cm1iw6, Jm1iw6, Qm1iw6, Xm1iw6, En1iw6, Ln1iw6, Sn1iw6;
wire Zn1iw6, Go1iw6, No1iw6, Uo1iw6, Bp1iw6, Ip1iw6, Pp1iw6, Wp1iw6, Dq1iw6, Kq1iw6;
wire Rq1iw6, Yq1iw6, Fr1iw6, Mr1iw6, Tr1iw6, As1iw6, Hs1iw6, Os1iw6, Vs1iw6, Ct1iw6;
wire Jt1iw6, Qt1iw6, Xt1iw6, Eu1iw6, Lu1iw6, Su1iw6, Zu1iw6, Gv1iw6, Nv1iw6, Uv1iw6;
wire Bw1iw6, Iw1iw6, Pw1iw6, Ww1iw6, Dx1iw6, Kx1iw6, Rx1iw6, Yx1iw6, Fy1iw6, My1iw6;
wire Ty1iw6, Az1iw6, Hz1iw6, Oz1iw6, Vz1iw6, C02iw6, J02iw6, Q02iw6, X02iw6, E12iw6;
wire L12iw6, S12iw6, Z12iw6, G22iw6, N22iw6, U22iw6, B32iw6, I32iw6, P32iw6, W32iw6;
wire D42iw6, K42iw6, R42iw6, Y42iw6, F52iw6, M52iw6, T52iw6, A62iw6, H62iw6, O62iw6;
wire V62iw6, C72iw6, J72iw6, Q72iw6, X72iw6, E82iw6, L82iw6, S82iw6, Z82iw6, G92iw6;
wire N92iw6, U92iw6, Ba2iw6, Ia2iw6, Pa2iw6, Wa2iw6, Db2iw6, Kb2iw6, Rb2iw6, Yb2iw6;
wire Fc2iw6, Mc2iw6, Tc2iw6, Ad2iw6, Hd2iw6, Od2iw6, Vd2iw6, Ce2iw6, Je2iw6, Qe2iw6;
wire Xe2iw6, Ef2iw6, Lf2iw6, Sf2iw6, Zf2iw6, Gg2iw6, Ng2iw6, Ug2iw6, Bh2iw6, Ih2iw6;
wire Ph2iw6, Wh2iw6, Di2iw6, Ki2iw6, Ri2iw6, Yi2iw6, Fj2iw6, Mj2iw6, Tj2iw6, Ak2iw6;
wire Hk2iw6, Ok2iw6, Vk2iw6, Cl2iw6, Jl2iw6, Ql2iw6, Xl2iw6, Em2iw6, Lm2iw6, Sm2iw6;
wire Zm2iw6, Gn2iw6, Nn2iw6, Un2iw6, Bo2iw6, Io2iw6, Po2iw6, Wo2iw6, Dp2iw6, Kp2iw6;
wire Rp2iw6, Yp2iw6, Fq2iw6, Mq2iw6, Tq2iw6, Ar2iw6, Hr2iw6, Or2iw6, Vr2iw6, Cs2iw6;
wire Js2iw6, Qs2iw6, Xs2iw6, Et2iw6, Lt2iw6, St2iw6, Zt2iw6, Gu2iw6, Nu2iw6, Uu2iw6;
wire Bv2iw6, Iv2iw6, Pv2iw6, Wv2iw6, Dw2iw6, Kw2iw6, Rw2iw6, Yw2iw6, Fx2iw6, Mx2iw6;
wire Tx2iw6, Ay2iw6, Hy2iw6, Oy2iw6, Vy2iw6, Cz2iw6, Jz2iw6, Qz2iw6, Xz2iw6, E03iw6;
wire L03iw6, S03iw6, Z03iw6, G13iw6, N13iw6, U13iw6, B23iw6, I23iw6, P23iw6, W23iw6;
wire D33iw6, K33iw6, R33iw6, Y33iw6, F43iw6, M43iw6, T43iw6, A53iw6, H53iw6, O53iw6;
wire V53iw6, C63iw6, J63iw6, Q63iw6, X63iw6, E73iw6, L73iw6, S73iw6, Z73iw6, G83iw6;
wire N83iw6, U83iw6, B93iw6, I93iw6, P93iw6, W93iw6, Da3iw6, Ka3iw6, Ra3iw6, Ya3iw6;
wire Fb3iw6, Mb3iw6, Tb3iw6, Ac3iw6, Hc3iw6, Oc3iw6, Vc3iw6, Cd3iw6, Jd3iw6, Qd3iw6;
wire Xd3iw6, Ee3iw6, Le3iw6, Se3iw6, Ze3iw6, Gf3iw6, Nf3iw6, Uf3iw6, Bg3iw6, Ig3iw6;
wire Pg3iw6, Wg3iw6, Dh3iw6, Kh3iw6, Rh3iw6, Yh3iw6, Fi3iw6, Mi3iw6, Ti3iw6, Aj3iw6;
wire Hj3iw6, Oj3iw6, Vj3iw6, Ck3iw6, Jk3iw6, Qk3iw6, Xk3iw6, El3iw6, Ll3iw6, Sl3iw6;
wire Zl3iw6, Gm3iw6, Nm3iw6, Um3iw6, Bn3iw6, In3iw6, Pn3iw6, Wn3iw6, Do3iw6, Ko3iw6;
wire Ro3iw6, Yo3iw6, Fp3iw6, Mp3iw6, Tp3iw6, Aq3iw6, Hq3iw6, Oq3iw6, Vq3iw6, Cr3iw6;
wire Jr3iw6, Qr3iw6, Xr3iw6, Es3iw6, Ls3iw6, Ss3iw6, Zs3iw6, Gt3iw6, Nt3iw6, Ut3iw6;
wire Bu3iw6, Iu3iw6, Pu3iw6, Wu3iw6, Dv3iw6, Kv3iw6, Rv3iw6, Yv3iw6, Fw3iw6, Mw3iw6;
wire Tw3iw6, Ax3iw6, Hx3iw6, Ox3iw6, Vx3iw6, Cy3iw6, Jy3iw6, Qy3iw6, Xy3iw6, Ez3iw6;
wire Lz3iw6, Sz3iw6, Zz3iw6, G04iw6, N04iw6, U04iw6, B14iw6, I14iw6, P14iw6, W14iw6;
wire D24iw6, K24iw6, R24iw6, Y24iw6, F34iw6, M34iw6, T34iw6, A44iw6, H44iw6, O44iw6;
wire V44iw6, C54iw6, J54iw6, Q54iw6, X54iw6, E64iw6, L64iw6, S64iw6, Z64iw6, G74iw6;
wire N74iw6, U74iw6, B84iw6, I84iw6, P84iw6, W84iw6, D94iw6, K94iw6, R94iw6, Y94iw6;
wire Fa4iw6, Ma4iw6, Ta4iw6, Ab4iw6, Hb4iw6, Ob4iw6, Vb4iw6, Cc4iw6, Jc4iw6, Qc4iw6;
wire Xc4iw6, Ed4iw6, Ld4iw6, Sd4iw6, Zd4iw6, Ge4iw6, Ne4iw6, Ue4iw6, Bf4iw6, If4iw6;
wire Pf4iw6, Wf4iw6, Dg4iw6, Kg4iw6, Rg4iw6, Yg4iw6, Fh4iw6, Mh4iw6, Th4iw6, Ai4iw6;
wire Hi4iw6, Oi4iw6, Vi4iw6, Cj4iw6, Jj4iw6, Qj4iw6, Xj4iw6, Ek4iw6, Lk4iw6, Sk4iw6;
wire Zk4iw6, Gl4iw6, Nl4iw6, Ul4iw6, Bm4iw6, Im4iw6, Pm4iw6, Wm4iw6, Dn4iw6, Kn4iw6;
wire Rn4iw6, Yn4iw6, Fo4iw6, Mo4iw6, To4iw6, Ap4iw6, Hp4iw6, Op4iw6, Vp4iw6, Cq4iw6;
wire Jq4iw6, Qq4iw6, Xq4iw6, Er4iw6, Lr4iw6, Sr4iw6, Zr4iw6, Gs4iw6, Ns4iw6, Us4iw6;
wire Bt4iw6, It4iw6, Pt4iw6, Wt4iw6, Du4iw6, Ku4iw6, Ru4iw6, Yu4iw6, Fv4iw6, Mv4iw6;
wire Tv4iw6, Aw4iw6, Hw4iw6, Ow4iw6, Vw4iw6, Cx4iw6, Jx4iw6, Qx4iw6, Xx4iw6, Ey4iw6;
wire Ly4iw6, Sy4iw6, Zy4iw6, Gz4iw6, Nz4iw6, Uz4iw6, B05iw6, I05iw6, P05iw6, W05iw6;
wire D15iw6, K15iw6, R15iw6, Y15iw6, F25iw6, M25iw6, T25iw6, A35iw6, H35iw6, O35iw6;
wire V35iw6, C45iw6, J45iw6, Q45iw6, X45iw6, E55iw6, L55iw6, S55iw6, Z55iw6, G65iw6;
wire N65iw6, U65iw6, B75iw6, I75iw6, P75iw6, W75iw6, D85iw6, K85iw6, R85iw6, Y85iw6;
wire F95iw6, M95iw6, T95iw6, Aa5iw6, Ha5iw6, Oa5iw6, Va5iw6, Cb5iw6, Jb5iw6, Qb5iw6;
wire Xb5iw6, Ec5iw6, Lc5iw6, Sc5iw6, Zc5iw6, Gd5iw6, Nd5iw6, Ud5iw6, Be5iw6, Ie5iw6;
wire Pe5iw6, We5iw6, Df5iw6, Kf5iw6, Rf5iw6, Yf5iw6, Fg5iw6, Mg5iw6, Tg5iw6, Ah5iw6;
wire Hh5iw6, Oh5iw6, Vh5iw6, Ci5iw6, Ji5iw6, Qi5iw6, Xi5iw6, Ej5iw6, Lj5iw6, Sj5iw6;
wire Zj5iw6, Gk5iw6, Nk5iw6, Uk5iw6, Bl5iw6, Il5iw6, Pl5iw6, Wl5iw6, Dm5iw6, Km5iw6;
wire Rm5iw6, Ym5iw6, Fn5iw6, Mn5iw6, Tn5iw6, Ao5iw6, Ho5iw6, Oo5iw6, Vo5iw6, Cp5iw6;
wire Jp5iw6, Qp5iw6, Xp5iw6, Eq5iw6, Lq5iw6, Sq5iw6, Zq5iw6, Gr5iw6, Nr5iw6, Ur5iw6;
wire Bs5iw6, Is5iw6, Ps5iw6, Ws5iw6, Dt5iw6, Kt5iw6, Rt5iw6, Yt5iw6, Fu5iw6, Mu5iw6;
wire Tu5iw6, Av5iw6, Hv5iw6, Ov5iw6, Vv5iw6, Cw5iw6, Jw5iw6, Qw5iw6, Xw5iw6, Ex5iw6;
wire Lx5iw6, Sx5iw6, Zx5iw6, Gy5iw6, Ny5iw6, Uy5iw6, Bz5iw6, Iz5iw6, Pz5iw6, Wz5iw6;
wire D06iw6, K06iw6, R06iw6, Y06iw6, F16iw6, M16iw6, T16iw6, A26iw6, H26iw6, O26iw6;
wire V26iw6, C36iw6, J36iw6, Q36iw6, X36iw6, E46iw6, L46iw6, S46iw6, Z46iw6, G56iw6;
wire N56iw6, U56iw6, B66iw6, I66iw6, P66iw6, W66iw6, D76iw6, K76iw6, R76iw6, Y76iw6;
wire F86iw6, M86iw6, T86iw6, A96iw6, H96iw6, O96iw6, V96iw6, Ca6iw6, Ja6iw6, Qa6iw6;
wire Xa6iw6, Eb6iw6, Lb6iw6, Sb6iw6, Zb6iw6, Gc6iw6, Nc6iw6, Uc6iw6, Bd6iw6, Id6iw6;
wire Pd6iw6, Wd6iw6, De6iw6, Ke6iw6, Re6iw6, Ye6iw6, Ff6iw6, Mf6iw6, Tf6iw6, Ag6iw6;
wire Hg6iw6, Og6iw6, Vg6iw6, Ch6iw6, Jh6iw6, Qh6iw6, Xh6iw6, Ei6iw6, Li6iw6, Si6iw6;
wire Zi6iw6, Gj6iw6, Nj6iw6, Uj6iw6, Bk6iw6, Ik6iw6, Pk6iw6, Wk6iw6, Dl6iw6, Kl6iw6;
wire Rl6iw6, Yl6iw6, Fm6iw6, Mm6iw6, Tm6iw6, An6iw6, Hn6iw6, On6iw6, Vn6iw6, Co6iw6;
wire Jo6iw6, Qo6iw6, Xo6iw6, Ep6iw6, Lp6iw6, Sp6iw6, Zp6iw6, Gq6iw6, Nq6iw6, Uq6iw6;
wire Br6iw6, Ir6iw6, Pr6iw6, Wr6iw6, Ds6iw6, Ks6iw6, Rs6iw6, Ys6iw6, Ft6iw6, Mt6iw6;
wire Tt6iw6, Au6iw6, Hu6iw6, Ou6iw6, Vu6iw6, Cv6iw6, Jv6iw6, Qv6iw6, Xv6iw6, Ew6iw6;
wire Lw6iw6, Sw6iw6, Zw6iw6, Gx6iw6, Nx6iw6, Ux6iw6, By6iw6, Iy6iw6, Py6iw6, Wy6iw6;
wire Dz6iw6, Kz6iw6, Rz6iw6, Yz6iw6, F07iw6, M07iw6, T07iw6, A17iw6, H17iw6, O17iw6;
wire V17iw6, C27iw6, J27iw6, Q27iw6, X27iw6, E37iw6, L37iw6, S37iw6, Z37iw6, G47iw6;
wire N47iw6, U47iw6, B57iw6, I57iw6, P57iw6, W57iw6, D67iw6, K67iw6, R67iw6, Y67iw6;
wire F77iw6, M77iw6, T77iw6, A87iw6, H87iw6, O87iw6, V87iw6, C97iw6, J97iw6, Q97iw6;
wire X97iw6, Ea7iw6, La7iw6, Sa7iw6, Za7iw6, Gb7iw6, Nb7iw6, Ub7iw6, Bc7iw6, Ic7iw6;
wire Pc7iw6, Wc7iw6, Dd7iw6, Kd7iw6, Rd7iw6, Yd7iw6, Fe7iw6, Me7iw6, Te7iw6, Af7iw6;
wire Hf7iw6, Of7iw6, Vf7iw6, Cg7iw6, Jg7iw6, Qg7iw6, Xg7iw6, Eh7iw6, Lh7iw6, Sh7iw6;
wire Zh7iw6, Gi7iw6, Ni7iw6, Ui7iw6, Bj7iw6, Ij7iw6, Pj7iw6, Wj7iw6, Dk7iw6, Kk7iw6;
wire Rk7iw6, Yk7iw6, Fl7iw6, Ml7iw6, Tl7iw6, Am7iw6, Hm7iw6, Om7iw6, Vm7iw6, Cn7iw6;
wire Jn7iw6, Qn7iw6, Xn7iw6, Eo7iw6, Lo7iw6, So7iw6, Zo7iw6, Gp7iw6, Np7iw6, Up7iw6;
wire Bq7iw6, Iq7iw6, Pq7iw6, Wq7iw6, Dr7iw6, Kr7iw6, Rr7iw6, Yr7iw6, Fs7iw6, Ms7iw6;
wire Ts7iw6, At7iw6, Ht7iw6, Ot7iw6, Vt7iw6, Cu7iw6, Ju7iw6, Qu7iw6, Xu7iw6, Ev7iw6;
wire Lv7iw6, Sv7iw6, Zv7iw6, Gw7iw6, Nw7iw6, Uw7iw6, Bx7iw6, Ix7iw6, Px7iw6, Wx7iw6;
wire Dy7iw6, Ky7iw6, Ry7iw6, Yy7iw6, Fz7iw6, Mz7iw6, Tz7iw6, A08iw6, H08iw6, O08iw6;
wire V08iw6, C18iw6, J18iw6, Q18iw6, X18iw6, E28iw6, L28iw6, S28iw6, Z28iw6, G38iw6;
wire N38iw6, U38iw6, B48iw6, I48iw6, P48iw6, W48iw6, D58iw6, K58iw6, R58iw6, Y58iw6;
wire F68iw6, M68iw6, T68iw6, A78iw6, H78iw6, O78iw6, V78iw6, C88iw6, J88iw6, Q88iw6;
wire X88iw6, E98iw6, L98iw6, S98iw6, Z98iw6, Ga8iw6, Na8iw6, Ua8iw6, Bb8iw6, Ib8iw6;
wire Pb8iw6, Wb8iw6, Dc8iw6, Kc8iw6, Rc8iw6, Yc8iw6, Fd8iw6, Md8iw6, Td8iw6, Ae8iw6;
wire He8iw6, Oe8iw6, Ve8iw6, Cf8iw6, Jf8iw6, Qf8iw6, Xf8iw6, Eg8iw6, Lg8iw6, Sg8iw6;
wire Zg8iw6, Gh8iw6, Nh8iw6, Uh8iw6, Bi8iw6, Ii8iw6, Pi8iw6, Wi8iw6, Dj8iw6, Kj8iw6;
wire Rj8iw6, Yj8iw6, Fk8iw6, Mk8iw6, Tk8iw6, Al8iw6, Hl8iw6, Ol8iw6, Vl8iw6, Cm8iw6;
wire Jm8iw6, Qm8iw6, Xm8iw6, En8iw6, Ln8iw6, Sn8iw6, Zn8iw6, Go8iw6, No8iw6, Uo8iw6;
wire Bp8iw6, Ip8iw6, Pp8iw6, Wp8iw6, Dq8iw6, Kq8iw6, Rq8iw6, Yq8iw6, Fr8iw6, Mr8iw6;
wire Tr8iw6, As8iw6, Hs8iw6, Os8iw6, Vs8iw6, Ct8iw6, Jt8iw6, Qt8iw6, Xt8iw6, Eu8iw6;
wire Lu8iw6, Su8iw6, Zu8iw6, Gv8iw6, Nv8iw6, Uv8iw6, Bw8iw6, Iw8iw6, Pw8iw6, Ww8iw6;
wire Dx8iw6, Kx8iw6, Rx8iw6, Yx8iw6, Fy8iw6, My8iw6, Ty8iw6, Az8iw6, Hz8iw6, Oz8iw6;
wire Vz8iw6, C09iw6, J09iw6, Q09iw6, X09iw6, E19iw6, L19iw6, S19iw6, Z19iw6, G29iw6;
wire N29iw6, U29iw6, B39iw6, I39iw6, P39iw6, W39iw6, D49iw6, K49iw6, R49iw6, Y49iw6;
wire F59iw6, M59iw6, T59iw6, A69iw6, H69iw6, O69iw6, V69iw6, C79iw6, J79iw6, Q79iw6;
wire X79iw6, E89iw6, L89iw6, S89iw6, Z89iw6, G99iw6, N99iw6, U99iw6, Ba9iw6, Ia9iw6;
wire Pa9iw6, Wa9iw6, Db9iw6, Kb9iw6, Rb9iw6, Yb9iw6, Fc9iw6, Mc9iw6, Tc9iw6, Ad9iw6;
wire Hd9iw6, Od9iw6, Vd9iw6, Ce9iw6, Je9iw6, Qe9iw6, Xe9iw6, Ef9iw6, Lf9iw6, Sf9iw6;
wire Zf9iw6, Gg9iw6, Ng9iw6, Ug9iw6, Bh9iw6, Ih9iw6, Ph9iw6, Wh9iw6, Di9iw6, Ki9iw6;
wire Ri9iw6, Yi9iw6, Fj9iw6, Mj9iw6, Tj9iw6, Ak9iw6, Hk9iw6, Ok9iw6, Vk9iw6, Cl9iw6;
wire Jl9iw6, Ql9iw6, Xl9iw6, Em9iw6, Lm9iw6, Sm9iw6, Zm9iw6, Gn9iw6, Nn9iw6, Un9iw6;
wire Bo9iw6, Io9iw6, Po9iw6, Wo9iw6, Dp9iw6, Kp9iw6, Rp9iw6, Yp9iw6, Fq9iw6, Mq9iw6;
wire Tq9iw6, Ar9iw6, Hr9iw6, Or9iw6, Vr9iw6, Cs9iw6, Js9iw6, Qs9iw6, Xs9iw6, Et9iw6;
wire Lt9iw6, St9iw6, Zt9iw6, Gu9iw6, Nu9iw6, Uu9iw6, Bv9iw6, Iv9iw6, Pv9iw6, Wv9iw6;
wire Dw9iw6, Kw9iw6, Rw9iw6, Yw9iw6, Fx9iw6, Mx9iw6, Tx9iw6, Ay9iw6, Hy9iw6, Oy9iw6;
wire Vy9iw6, Cz9iw6, Jz9iw6, Qz9iw6, Xz9iw6, E0aiw6, L0aiw6, S0aiw6, Z0aiw6, G1aiw6;
wire N1aiw6, U1aiw6, B2aiw6, I2aiw6, P2aiw6, W2aiw6, D3aiw6, K3aiw6, R3aiw6, Y3aiw6;
wire F4aiw6, M4aiw6, T4aiw6, A5aiw6, H5aiw6, O5aiw6, V5aiw6, C6aiw6, J6aiw6, Q6aiw6;
wire X6aiw6, E7aiw6, L7aiw6, S7aiw6, Z7aiw6, G8aiw6, N8aiw6, U8aiw6, B9aiw6, I9aiw6;
wire P9aiw6, W9aiw6, Daaiw6, Kaaiw6, Raaiw6, Yaaiw6, Fbaiw6, Mbaiw6, Tbaiw6, Acaiw6;
wire Hcaiw6, Ocaiw6, Vcaiw6, Cdaiw6, Jdaiw6, Qdaiw6, Xdaiw6, Eeaiw6, Leaiw6, Seaiw6;
wire Zeaiw6, Gfaiw6, Nfaiw6, Ufaiw6, Bgaiw6, Igaiw6, Pgaiw6, Wgaiw6, Dhaiw6, Khaiw6;
wire Rhaiw6, Yhaiw6, Fiaiw6, Miaiw6, Tiaiw6, Ajaiw6, Hjaiw6, Ojaiw6, Vjaiw6, Ckaiw6;
wire Jkaiw6, Qkaiw6, Xkaiw6, Elaiw6, Llaiw6, Slaiw6, Zlaiw6, Gmaiw6, Nmaiw6, Umaiw6;
wire Bnaiw6, Inaiw6, Pnaiw6, Wnaiw6, Doaiw6, Koaiw6, Roaiw6, Yoaiw6, Fpaiw6, Mpaiw6;
wire Tpaiw6, Aqaiw6, Hqaiw6, Oqaiw6, Vqaiw6, Craiw6, Jraiw6, Qraiw6, Xraiw6, Esaiw6;
wire Lsaiw6, Ssaiw6, Zsaiw6, Gtaiw6, Ntaiw6, Utaiw6, Buaiw6, Iuaiw6, Puaiw6, Wuaiw6;
wire Dvaiw6, Kvaiw6, Rvaiw6, Yvaiw6, Fwaiw6, Mwaiw6, Twaiw6, Axaiw6, Hxaiw6, Oxaiw6;
wire Vxaiw6, Cyaiw6, Jyaiw6, Qyaiw6, Xyaiw6, Ezaiw6, Lzaiw6, Szaiw6, Zzaiw6, G0biw6;
wire N0biw6, U0biw6, B1biw6, I1biw6, P1biw6, W1biw6, D2biw6, K2biw6, R2biw6, Y2biw6;
wire F3biw6, M3biw6, T3biw6, A4biw6, H4biw6, O4biw6, V4biw6, C5biw6, J5biw6, Q5biw6;
wire X5biw6, E6biw6, L6biw6, S6biw6, Z6biw6, G7biw6, N7biw6, U7biw6, B8biw6, I8biw6;
wire P8biw6, W8biw6, D9biw6, K9biw6, R9biw6, Y9biw6, Fabiw6, Mabiw6, Tabiw6, Abbiw6;
wire Hbbiw6, Obbiw6, Vbbiw6, Ccbiw6, Jcbiw6, Qcbiw6, Xcbiw6, Edbiw6, Ldbiw6, Sdbiw6;
wire Zdbiw6, Gebiw6, Nebiw6, Uebiw6, Bfbiw6, Ifbiw6, Pfbiw6, Wfbiw6, Dgbiw6, Kgbiw6;
wire Rgbiw6, Ygbiw6, Fhbiw6, Mhbiw6, Thbiw6, Aibiw6, Hibiw6, Oibiw6, Vibiw6, Cjbiw6;
wire Jjbiw6, Qjbiw6, Xjbiw6, Ekbiw6, Lkbiw6, Skbiw6, Zkbiw6, Glbiw6, Nlbiw6, Ulbiw6;
wire Bmbiw6, Imbiw6, Pmbiw6, Wmbiw6, Dnbiw6, Knbiw6, Rnbiw6, Ynbiw6, Fobiw6, Mobiw6;
wire Tobiw6, Apbiw6, Hpbiw6, Opbiw6, Vpbiw6, Cqbiw6, Jqbiw6, Qqbiw6, Xqbiw6, Erbiw6;
wire Lrbiw6, Srbiw6, Zrbiw6, Gsbiw6, Nsbiw6, Usbiw6, Btbiw6, Itbiw6, Ptbiw6, Wtbiw6;
wire Dubiw6, Kubiw6, Rubiw6, Yubiw6, Fvbiw6, Mvbiw6, Tvbiw6, Awbiw6, Hwbiw6, Owbiw6;
wire Vwbiw6, Cxbiw6, Jxbiw6, Qxbiw6, Xxbiw6, Eybiw6, Lybiw6, Sybiw6, Zybiw6, Gzbiw6;
wire Nzbiw6, Uzbiw6, B0ciw6, I0ciw6, P0ciw6, W0ciw6, D1ciw6, K1ciw6, R1ciw6, Y1ciw6;
wire F2ciw6, M2ciw6, T2ciw6, A3ciw6, H3ciw6, O3ciw6, V3ciw6, C4ciw6, J4ciw6, Q4ciw6;
wire X4ciw6, E5ciw6, L5ciw6, S5ciw6, Z5ciw6, G6ciw6, N6ciw6, U6ciw6, B7ciw6, I7ciw6;
wire P7ciw6, W7ciw6, D8ciw6, K8ciw6, R8ciw6, Y8ciw6, F9ciw6, M9ciw6, T9ciw6, Aaciw6;
wire Haciw6, Oaciw6, Vaciw6, Cbciw6, Jbciw6, Qbciw6, Xbciw6, Ecciw6, Lcciw6, Scciw6;
wire Zcciw6, Gdciw6, Ndciw6, Udciw6, Beciw6, Ieciw6, Peciw6, Weciw6, Dfciw6, Kfciw6;
wire Rfciw6, Yfciw6, Fgciw6, Mgciw6, Tgciw6, Ahciw6, Hhciw6, Ohciw6, Vhciw6, Ciciw6;
wire Jiciw6, Qiciw6, Xiciw6, Ejciw6, Ljciw6, Sjciw6, Zjciw6, Gkciw6, Nkciw6, Ukciw6;
wire Blciw6, Ilciw6, Plciw6, Wlciw6, Dmciw6, Kmciw6, Rmciw6, Ymciw6, Fnciw6, Mnciw6;
wire Tnciw6, Aociw6, Hociw6, Oociw6, Vociw6, Cpciw6, Jpciw6, Qpciw6, Xpciw6, Eqciw6;
wire Lqciw6, Sqciw6, Zqciw6, Grciw6, Nrciw6, Urciw6, Bsciw6, Isciw6, Psciw6, Wsciw6;
wire Dtciw6, Ktciw6, Rtciw6, Ytciw6, Fuciw6, Muciw6, Tuciw6, Avciw6, Hvciw6, Ovciw6;
wire Vvciw6, Cwciw6, Jwciw6, Qwciw6, Xwciw6, Exciw6, Lxciw6, Sxciw6, Zxciw6, Gyciw6;
wire Nyciw6, Uyciw6, Bzciw6, Izciw6, Pzciw6, Wzciw6, D0diw6, K0diw6, R0diw6, Y0diw6;
wire F1diw6, M1diw6, T1diw6, A2diw6, H2diw6, O2diw6, V2diw6, C3diw6, J3diw6, Q3diw6;
wire X3diw6, E4diw6, L4diw6, S4diw6, Z4diw6, G5diw6, N5diw6, U5diw6, B6diw6, I6diw6;
wire P6diw6, W6diw6, D7diw6, K7diw6, R7diw6, Y7diw6, F8diw6, M8diw6, T8diw6, A9diw6;
wire H9diw6, O9diw6, V9diw6, Cadiw6, Jadiw6, Qadiw6, Xadiw6, Ebdiw6, Lbdiw6, Sbdiw6;
wire Zbdiw6, Gcdiw6, Ncdiw6, Ucdiw6, Bddiw6, Iddiw6, Pddiw6, Wddiw6, Dediw6, Kediw6;
wire Rediw6, Yediw6, Ffdiw6, Mfdiw6, Tfdiw6, Agdiw6, Hgdiw6, Ogdiw6, Vgdiw6, Chdiw6;
wire Jhdiw6, Qhdiw6, Xhdiw6, Eidiw6, Lidiw6, Sidiw6, Zidiw6, Gjdiw6, Njdiw6, Ujdiw6;
wire Bkdiw6, Ikdiw6, Pkdiw6, Wkdiw6, Dldiw6, Kldiw6, Rldiw6, Yldiw6, Fmdiw6, Mmdiw6;
wire Tmdiw6, Andiw6, Hndiw6, Ondiw6, Vndiw6, Codiw6, Jodiw6, Qodiw6, Xodiw6, Epdiw6;
wire Lpdiw6, Spdiw6, Zpdiw6, Gqdiw6, Nqdiw6, Uqdiw6, Brdiw6, Irdiw6, Prdiw6, Wrdiw6;
wire Dsdiw6, Ksdiw6, Rsdiw6, Ysdiw6, Ftdiw6, Mtdiw6, Ttdiw6, Audiw6, Hudiw6, Oudiw6;
wire Vudiw6, Cvdiw6, Jvdiw6, Qvdiw6, Xvdiw6, Ewdiw6, Lwdiw6, Swdiw6, Zwdiw6, Gxdiw6;
wire Nxdiw6, Uxdiw6, Bydiw6, Iydiw6, Pydiw6, Wydiw6, Dzdiw6, Kzdiw6, Rzdiw6, Yzdiw6;
wire F0eiw6, M0eiw6, T0eiw6, A1eiw6, H1eiw6, O1eiw6, V1eiw6, C2eiw6, J2eiw6, Q2eiw6;
wire X2eiw6, E3eiw6, L3eiw6, S3eiw6, Z3eiw6, G4eiw6, N4eiw6, U4eiw6, B5eiw6, I5eiw6;
wire P5eiw6, W5eiw6, D6eiw6, K6eiw6, R6eiw6, Y6eiw6, F7eiw6, M7eiw6, T7eiw6, A8eiw6;
wire H8eiw6, O8eiw6, V8eiw6, C9eiw6, J9eiw6, Q9eiw6, X9eiw6, Eaeiw6, Laeiw6, Saeiw6;
wire Zaeiw6, Gbeiw6, Nbeiw6, Ubeiw6, Bceiw6, Iceiw6, Pceiw6, Wceiw6, Ddeiw6, Kdeiw6;
wire Rdeiw6, Ydeiw6, Feeiw6, Meeiw6, Teeiw6, Afeiw6, Hfeiw6, Ofeiw6, Vfeiw6, Cgeiw6;
wire Jgeiw6, Qgeiw6, Xgeiw6, Eheiw6, Lheiw6, Sheiw6, Zheiw6, Gieiw6, Nieiw6, Uieiw6;
wire Bjeiw6, Ijeiw6, Pjeiw6, Wjeiw6, Dkeiw6, Kkeiw6, Rkeiw6, Ykeiw6, Fleiw6, Mleiw6;
wire Tleiw6, Ameiw6, Hmeiw6, Omeiw6, Vmeiw6, Cneiw6, Jneiw6, Qneiw6, Xneiw6, Eoeiw6;
wire Loeiw6, Soeiw6, Zoeiw6, Gpeiw6, Npeiw6, Upeiw6, Bqeiw6, Iqeiw6, Pqeiw6, Wqeiw6;
wire Dreiw6, Kreiw6, Rreiw6, Yreiw6, Fseiw6, Mseiw6, Tseiw6, Ateiw6, Hteiw6, Oteiw6;
wire Vteiw6, Cueiw6, Jueiw6, Queiw6, Xueiw6, Eveiw6, Lveiw6, Sveiw6, Zveiw6, Gweiw6;
wire Nweiw6, Uweiw6, Bxeiw6, Ixeiw6, Pxeiw6, Wxeiw6, Dyeiw6, Kyeiw6, Ryeiw6, Yyeiw6;
wire Fzeiw6, Mzeiw6, Tzeiw6, A0fiw6, H0fiw6, O0fiw6, V0fiw6, C1fiw6, J1fiw6, Q1fiw6;
wire X1fiw6, E2fiw6, L2fiw6, S2fiw6, Z2fiw6, G3fiw6, N3fiw6, U3fiw6, B4fiw6, I4fiw6;
wire P4fiw6, W4fiw6, D5fiw6, K5fiw6, R5fiw6, Y5fiw6, F6fiw6, M6fiw6, T6fiw6, A7fiw6;
wire H7fiw6, O7fiw6, V7fiw6, C8fiw6, J8fiw6, Q8fiw6, X8fiw6, E9fiw6, L9fiw6, S9fiw6;
wire Z9fiw6, Gafiw6, Nafiw6, Uafiw6, Bbfiw6, Ibfiw6, Pbfiw6, Wbfiw6, Dcfiw6, Kcfiw6;
wire Rcfiw6, Ycfiw6, Fdfiw6, Mdfiw6, Tdfiw6, Aefiw6, Hefiw6, Oefiw6, Vefiw6, Cffiw6;
wire Jffiw6, Qffiw6, Xffiw6, Egfiw6, Lgfiw6, Sgfiw6, Zgfiw6, Ghfiw6, Nhfiw6, Uhfiw6;
wire Bifiw6, Iifiw6, Pifiw6, Wifiw6, Djfiw6, Kjfiw6, Rjfiw6, Yjfiw6, Fkfiw6, Mkfiw6;
wire Tkfiw6, Alfiw6, Hlfiw6, Olfiw6, Vlfiw6, Cmfiw6, Jmfiw6, Qmfiw6, Xmfiw6, Enfiw6;
wire Lnfiw6, Snfiw6, Znfiw6, Gofiw6, Nofiw6, Uofiw6, Bpfiw6, Ipfiw6, Ppfiw6, Wpfiw6;
wire Dqfiw6, Kqfiw6, Rqfiw6, Yqfiw6, Frfiw6, Mrfiw6, Trfiw6, Asfiw6, Hsfiw6, Osfiw6;
wire Vsfiw6, Ctfiw6, Jtfiw6, Qtfiw6, Xtfiw6, Eufiw6, Lufiw6, Sufiw6, Zufiw6, Gvfiw6;
wire Nvfiw6, Uvfiw6, Bwfiw6, Iwfiw6, Pwfiw6, Wwfiw6, Dxfiw6, Kxfiw6, Rxfiw6, Yxfiw6;
wire Fyfiw6, Myfiw6, Tyfiw6, Azfiw6, Hzfiw6, Ozfiw6, Vzfiw6, C0giw6, J0giw6, Q0giw6;
wire X0giw6, E1giw6, L1giw6, S1giw6, Z1giw6, G2giw6, N2giw6, U2giw6, B3giw6, I3giw6;
wire P3giw6, W3giw6, D4giw6, K4giw6, R4giw6, Y4giw6, F5giw6, M5giw6, T5giw6, A6giw6;
wire H6giw6, O6giw6, V6giw6, C7giw6, J7giw6, Q7giw6, X7giw6, E8giw6, L8giw6, S8giw6;
wire Z8giw6, G9giw6, N9giw6, U9giw6, Bagiw6, Iagiw6, Pagiw6, Wagiw6, Dbgiw6, Kbgiw6;
wire Rbgiw6, Ybgiw6, Fcgiw6, Mcgiw6, Tcgiw6, Adgiw6, Hdgiw6, Odgiw6, Vdgiw6, Cegiw6;
wire Jegiw6, Qegiw6, Xegiw6, Efgiw6, Lfgiw6, Sfgiw6, Zfgiw6, Gggiw6, Nggiw6, Uggiw6;
wire Bhgiw6, Ihgiw6, Phgiw6, Whgiw6, Digiw6, Kigiw6, Rigiw6, Yigiw6, Fjgiw6, Mjgiw6;
wire Tjgiw6, Akgiw6, Hkgiw6, Okgiw6, Vkgiw6, Clgiw6, Jlgiw6, Qlgiw6, Xlgiw6, Emgiw6;
wire Lmgiw6, Smgiw6, Zmgiw6, Gngiw6, Nngiw6, Ungiw6, Bogiw6, Iogiw6, Pogiw6, Wogiw6;
wire Dpgiw6, Kpgiw6, Rpgiw6, Ypgiw6, Fqgiw6, Mqgiw6, Tqgiw6, Argiw6, Hrgiw6, Orgiw6;
wire Vrgiw6, Csgiw6, Jsgiw6, Qsgiw6, Xsgiw6, Etgiw6, Ltgiw6, Stgiw6, Ztgiw6, Gugiw6;
wire Nugiw6, Uugiw6, Bvgiw6, Ivgiw6, Pvgiw6, Wvgiw6, Dwgiw6, Kwgiw6, Rwgiw6, Ywgiw6;
wire Fxgiw6, Mxgiw6, Txgiw6, Aygiw6, Hygiw6, Oygiw6, Vygiw6, Czgiw6, Jzgiw6, Qzgiw6;
wire Xzgiw6, E0hiw6, L0hiw6, S0hiw6, Z0hiw6, G1hiw6, N1hiw6, U1hiw6, B2hiw6, I2hiw6;
wire P2hiw6, W2hiw6, D3hiw6, K3hiw6, R3hiw6, Y3hiw6, F4hiw6, M4hiw6, T4hiw6, A5hiw6;
wire H5hiw6, O5hiw6, V5hiw6, C6hiw6, J6hiw6, Q6hiw6, X6hiw6, E7hiw6, L7hiw6, S7hiw6;
wire Z7hiw6, G8hiw6, N8hiw6, U8hiw6, B9hiw6, I9hiw6, P9hiw6, W9hiw6, Dahiw6, Kahiw6;
wire Rahiw6, Yahiw6, Fbhiw6, Mbhiw6, Tbhiw6, Achiw6, Hchiw6, Ochiw6, Vchiw6, Cdhiw6;
wire Jdhiw6, Qdhiw6, Xdhiw6, Eehiw6, Lehiw6, Sehiw6, Zehiw6, Gfhiw6, Nfhiw6, Ufhiw6;
wire Bghiw6, Ighiw6, Pghiw6, Wghiw6, Dhhiw6, Khhiw6, Rhhiw6, Yhhiw6, Fihiw6, Mihiw6;
wire Tihiw6, Ajhiw6, Hjhiw6, Ojhiw6, Vjhiw6, Ckhiw6, Jkhiw6, Qkhiw6, Xkhiw6, Elhiw6;
wire Llhiw6, Slhiw6, Zlhiw6, Gmhiw6, Nmhiw6, Umhiw6, Bnhiw6, Inhiw6, Pnhiw6, Wnhiw6;
wire Dohiw6, Kohiw6, Rohiw6, Yohiw6, Fphiw6, Mphiw6, Tphiw6, Aqhiw6, Hqhiw6, Oqhiw6;
wire Vqhiw6, Crhiw6, Jrhiw6, Qrhiw6, Xrhiw6, Eshiw6, Lshiw6, Sshiw6, Zshiw6, Gthiw6;
wire Nthiw6, Uthiw6, Buhiw6, Iuhiw6, Puhiw6, Wuhiw6, Dvhiw6, Kvhiw6, Rvhiw6, Yvhiw6;
wire Fwhiw6, Mwhiw6, Twhiw6, Axhiw6, Hxhiw6, Oxhiw6, Vxhiw6, Cyhiw6, Jyhiw6, Qyhiw6;
wire Xyhiw6, Ezhiw6, Lzhiw6, Szhiw6, Zzhiw6, G0iiw6, N0iiw6, U0iiw6, B1iiw6, I1iiw6;
wire P1iiw6, W1iiw6, D2iiw6, K2iiw6, R2iiw6, Y2iiw6, F3iiw6, M3iiw6, T3iiw6, A4iiw6;
wire H4iiw6, O4iiw6, V4iiw6, C5iiw6, J5iiw6, Q5iiw6, X5iiw6, E6iiw6, L6iiw6, S6iiw6;
wire Z6iiw6, G7iiw6, N7iiw6, U7iiw6, B8iiw6, I8iiw6, P8iiw6, W8iiw6, D9iiw6, K9iiw6;
wire R9iiw6, Y9iiw6, Faiiw6, Maiiw6, Taiiw6, Abiiw6, Hbiiw6, Obiiw6, Vbiiw6, Cciiw6;
wire Jciiw6, Qciiw6, Xciiw6, Ediiw6, Ldiiw6, Sdiiw6, Zdiiw6, Geiiw6, Neiiw6, Ueiiw6;
wire Bfiiw6, Ifiiw6, Pfiiw6, Wfiiw6, Dgiiw6, Kgiiw6, Rgiiw6, Ygiiw6, Fhiiw6, Mhiiw6;
wire Thiiw6, Aiiiw6, Hiiiw6, Oiiiw6, Viiiw6, Cjiiw6, Jjiiw6, Qjiiw6, Xjiiw6, Ekiiw6;
wire Lkiiw6, Skiiw6, Zkiiw6, Gliiw6, Nliiw6, Uliiw6, Bmiiw6, Imiiw6, Pmiiw6, Wmiiw6;
wire Dniiw6, Kniiw6, Rniiw6, Yniiw6, Foiiw6, Moiiw6, Toiiw6, Apiiw6, Hpiiw6, Opiiw6;
wire Vpiiw6, Cqiiw6, Jqiiw6, Qqiiw6, Xqiiw6, Eriiw6, Lriiw6, Sriiw6, Zriiw6, Gsiiw6;
wire Nsiiw6, Usiiw6, Btiiw6, Itiiw6, Ptiiw6, Wtiiw6, Duiiw6, Kuiiw6, Ruiiw6, Yuiiw6;
wire Fviiw6, Mviiw6, Tviiw6, Awiiw6, Hwiiw6, Owiiw6, Vwiiw6, Cxiiw6, Jxiiw6, Qxiiw6;
wire Xxiiw6, Eyiiw6, Lyiiw6, Syiiw6, Zyiiw6, Gziiw6, Nziiw6, Uziiw6, B0jiw6, I0jiw6;
wire P0jiw6, W0jiw6, D1jiw6, K1jiw6, R1jiw6, Y1jiw6, F2jiw6, M2jiw6, T2jiw6, A3jiw6;
wire H3jiw6, O3jiw6, V3jiw6, C4jiw6, J4jiw6, Q4jiw6, X4jiw6, E5jiw6, L5jiw6, S5jiw6;
wire Z5jiw6, G6jiw6, N6jiw6, U6jiw6, B7jiw6, I7jiw6, P7jiw6, W7jiw6, D8jiw6, K8jiw6;
wire R8jiw6, Y8jiw6, F9jiw6, M9jiw6, T9jiw6, Aajiw6, Hajiw6, Oajiw6, Vajiw6, Cbjiw6;
wire Jbjiw6, Qbjiw6, Xbjiw6, Ecjiw6, Lcjiw6, Scjiw6, Zcjiw6, Gdjiw6, Ndjiw6, Udjiw6;
wire Bejiw6, Iejiw6, Pejiw6, Wejiw6, Dfjiw6, Kfjiw6, Rfjiw6, Yfjiw6, Fgjiw6, Mgjiw6;
wire Tgjiw6, Ahjiw6, Hhjiw6, Ohjiw6, Vhjiw6, Cijiw6, Jijiw6, Qijiw6, Xijiw6, Ejjiw6;
wire Ljjiw6, Sjjiw6, Zjjiw6, Gkjiw6, Nkjiw6, Ukjiw6, Bljiw6, Iljiw6, Pljiw6, Wljiw6;
wire Dmjiw6, Kmjiw6, Rmjiw6, Ymjiw6, Fnjiw6, Mnjiw6, Tnjiw6, Aojiw6, Hojiw6, Oojiw6;
wire Vojiw6, Cpjiw6, Jpjiw6, Qpjiw6, Xpjiw6, Eqjiw6, Lqjiw6, Sqjiw6, Zqjiw6, Grjiw6;
wire Nrjiw6, Urjiw6, Bsjiw6, Isjiw6, Psjiw6, Wsjiw6, Dtjiw6, Ktjiw6, Rtjiw6, Ytjiw6;
wire Fujiw6, Mujiw6, Tujiw6, Avjiw6, Hvjiw6, Ovjiw6, Vvjiw6, Cwjiw6, Jwjiw6, Qwjiw6;
wire Xwjiw6, Exjiw6, Lxjiw6, Sxjiw6, Zxjiw6, Gyjiw6, Nyjiw6, Uyjiw6, Bzjiw6, Izjiw6;
wire Pzjiw6, Wzjiw6, D0kiw6, K0kiw6, R0kiw6, Y0kiw6, F1kiw6, M1kiw6, T1kiw6, A2kiw6;
wire H2kiw6, O2kiw6, V2kiw6, C3kiw6, J3kiw6, Q3kiw6, X3kiw6, E4kiw6, L4kiw6, S4kiw6;
wire Z4kiw6, G5kiw6, N5kiw6, U5kiw6, B6kiw6, I6kiw6, P6kiw6, W6kiw6, D7kiw6, K7kiw6;
wire R7kiw6, Y7kiw6, F8kiw6, M8kiw6, T8kiw6, A9kiw6, H9kiw6, O9kiw6, V9kiw6, Cakiw6;
wire Jakiw6, Qakiw6, Xakiw6, Ebkiw6, Lbkiw6, Sbkiw6, Zbkiw6, Gckiw6, Nckiw6, Uckiw6;
wire Bdkiw6, Idkiw6, Pdkiw6, Wdkiw6, Dekiw6, Kekiw6, Rekiw6, Yekiw6, Ffkiw6, Mfkiw6;
wire Tfkiw6, Agkiw6, Hgkiw6, Ogkiw6, Vgkiw6, Chkiw6, Jhkiw6, Qhkiw6, Xhkiw6, Eikiw6;
wire Likiw6, Sikiw6, Zikiw6, Gjkiw6, Njkiw6, Ujkiw6, Bkkiw6, Ikkiw6, Pkkiw6, Wkkiw6;
wire Dlkiw6, Klkiw6, Rlkiw6, Ylkiw6, Fmkiw6, Mmkiw6, Tmkiw6, Ankiw6, Hnkiw6, Onkiw6;
wire Vnkiw6, Cokiw6, Jokiw6, Qokiw6, Xokiw6, Epkiw6, Lpkiw6, Spkiw6, Zpkiw6, Gqkiw6;
wire Nqkiw6, Uqkiw6, Brkiw6, Irkiw6, Prkiw6, Wrkiw6, Dskiw6, Kskiw6, Rskiw6, Yskiw6;
wire Ftkiw6, Mtkiw6, Ttkiw6, Aukiw6, Hukiw6, Oukiw6, Vukiw6, Cvkiw6, Jvkiw6, Qvkiw6;
wire Xvkiw6, Ewkiw6, Lwkiw6, Swkiw6, Zwkiw6, Gxkiw6, Nxkiw6, Uxkiw6, Bykiw6, Iykiw6;
wire Pykiw6, Wykiw6, Dzkiw6, Kzkiw6, Rzkiw6, Yzkiw6, F0liw6, M0liw6, T0liw6, A1liw6;
wire H1liw6, O1liw6, V1liw6, C2liw6, J2liw6, Q2liw6, X2liw6, E3liw6, L3liw6, S3liw6;
wire Z3liw6, G4liw6, N4liw6, U4liw6, B5liw6, I5liw6, P5liw6, W5liw6, D6liw6, K6liw6;
wire R6liw6, Y6liw6, F7liw6, M7liw6, T7liw6, A8liw6, H8liw6, O8liw6, V8liw6, C9liw6;
wire J9liw6, Q9liw6, X9liw6, Ealiw6, Laliw6, Saliw6, Zaliw6, Gbliw6, Nbliw6, Ubliw6;
wire Bcliw6, Icliw6, Pcliw6, Wcliw6, Ddliw6, Kdliw6, Rdliw6, Ydliw6, Feliw6, Meliw6;
wire Teliw6, Afliw6, Hfliw6, Ofliw6, Vfliw6, Cgliw6, Jgliw6, Qgliw6, Xgliw6, Ehliw6;
wire Lhliw6, Shliw6, Zhliw6, Giliw6, Niliw6, Uiliw6, Bjliw6, Ijliw6, Pjliw6, Wjliw6;
wire Dkliw6, Kkliw6, Rkliw6, Ykliw6, Flliw6, Mlliw6, Tlliw6, Amliw6, Hmliw6, Omliw6;
wire Vmliw6, Cnliw6, Jnliw6, Qnliw6, Xnliw6, Eoliw6, Loliw6, Soliw6, Zoliw6, Gpliw6;
wire Npliw6, Upliw6, Bqliw6, Iqliw6, Pqliw6, Wqliw6, Drliw6, Krliw6, Rrliw6, Yrliw6;
wire Fsliw6, Msliw6, Tsliw6, Atliw6, Htliw6, Otliw6, Vtliw6, Culiw6, Juliw6, Quliw6;
wire Xuliw6, Evliw6, Lvliw6, Svliw6, Zvliw6, Gwliw6, Nwliw6, Uwliw6, Bxliw6, Ixliw6;
wire Pxliw6, Wxliw6, Dyliw6, Kyliw6, Ryliw6, Yyliw6, Fzliw6, Mzliw6, Tzliw6, A0miw6;
wire H0miw6, O0miw6, V0miw6, C1miw6, J1miw6, Q1miw6, X1miw6, E2miw6, L2miw6, S2miw6;
wire Z2miw6, G3miw6, N3miw6, U3miw6, B4miw6, I4miw6, P4miw6, W4miw6, D5miw6, K5miw6;
wire R5miw6, Y5miw6, F6miw6, M6miw6, T6miw6, A7miw6, H7miw6, O7miw6, V7miw6, C8miw6;
wire J8miw6, Q8miw6, X8miw6, E9miw6, L9miw6, S9miw6, Z9miw6, Gamiw6, Namiw6, Uamiw6;
wire Bbmiw6, Ibmiw6, Pbmiw6, Wbmiw6, Dcmiw6, Kcmiw6, Rcmiw6, Ycmiw6, Fdmiw6, Mdmiw6;
wire Tdmiw6, Aemiw6, Hemiw6, Oemiw6, Vemiw6, Cfmiw6, Jfmiw6, Qfmiw6, Xfmiw6, Egmiw6;
wire Lgmiw6, Sgmiw6, Zgmiw6, Ghmiw6, Nhmiw6, Uhmiw6, Bimiw6, Iimiw6, Pimiw6, Wimiw6;
wire Djmiw6, Kjmiw6, Rjmiw6, Yjmiw6, Fkmiw6, Mkmiw6, Tkmiw6, Almiw6, Hlmiw6, Olmiw6;
wire Vlmiw6, Cmmiw6, Jmmiw6, Qmmiw6, Xmmiw6, Enmiw6, Lnmiw6, Snmiw6, Znmiw6, Gomiw6;
wire Nomiw6, Uomiw6, Bpmiw6, Ipmiw6, Ppmiw6, Wpmiw6, Dqmiw6, Kqmiw6, Rqmiw6, Yqmiw6;
wire Frmiw6, Mrmiw6, Trmiw6, Asmiw6, Hsmiw6, Osmiw6, Vsmiw6, Ctmiw6, Jtmiw6, Qtmiw6;
wire Xtmiw6, Eumiw6, Lumiw6, Sumiw6, Zumiw6, Gvmiw6, Nvmiw6, Uvmiw6, Bwmiw6, Iwmiw6;
wire Pwmiw6, Wwmiw6, Dxmiw6, Kxmiw6, Rxmiw6, Yxmiw6, Fymiw6, Mymiw6, Tymiw6, Azmiw6;
wire Hzmiw6, Ozmiw6, Vzmiw6, C0niw6, J0niw6, Q0niw6, X0niw6, E1niw6, L1niw6, S1niw6;
wire Z1niw6, G2niw6, N2niw6, U2niw6, B3niw6, I3niw6, P3niw6, W3niw6, D4niw6, K4niw6;
wire R4niw6, Y4niw6, F5niw6, M5niw6, T5niw6, A6niw6, H6niw6, O6niw6, V6niw6, C7niw6;
wire J7niw6, Q7niw6, X7niw6, E8niw6, L8niw6, S8niw6, Z8niw6, G9niw6, N9niw6, U9niw6;
wire Baniw6, Ianiw6, Paniw6, Waniw6, Dbniw6, Kbniw6, Rbniw6, Ybniw6, Fcniw6, Mcniw6;
wire Tcniw6, Adniw6, Hdniw6, Odniw6, Vdniw6, Ceniw6, Jeniw6, Qeniw6, Xeniw6, Efniw6;
wire Lfniw6, Sfniw6, Zfniw6, Ggniw6, Ngniw6, Ugniw6, Bhniw6, Ihniw6, Phniw6, Whniw6;
wire Diniw6, Kiniw6, Riniw6, Yiniw6, Fjniw6, Mjniw6, Tjniw6, Akniw6, Hkniw6, Okniw6;
wire Vkniw6, Clniw6, Jlniw6, Qlniw6, Xlniw6, Emniw6, Lmniw6, Smniw6, Zmniw6, Gnniw6;
wire Nnniw6, Unniw6, Boniw6, Ioniw6, Poniw6, Woniw6, Dpniw6, Kpniw6, Rpniw6, Ypniw6;
wire Fqniw6, Mqniw6, Tqniw6, Arniw6, Hrniw6, Orniw6, Vrniw6, Csniw6, Jsniw6, Qsniw6;
wire Xsniw6, Etniw6, Ltniw6, Stniw6, Ztniw6, Guniw6, Nuniw6, Uuniw6, Bvniw6, Ivniw6;
wire Pvniw6, Wvniw6, Dwniw6, Kwniw6, Rwniw6, Ywniw6, Fxniw6, Mxniw6, Txniw6, Ayniw6;
wire Hyniw6, Oyniw6, Vyniw6, Czniw6, Jzniw6, Qzniw6, Xzniw6, E0oiw6, L0oiw6, S0oiw6;
wire Z0oiw6, G1oiw6, N1oiw6, U1oiw6, B2oiw6, I2oiw6, P2oiw6, W2oiw6, D3oiw6, K3oiw6;
wire R3oiw6, Y3oiw6, F4oiw6, M4oiw6, T4oiw6, A5oiw6, H5oiw6, O5oiw6, V5oiw6, C6oiw6;
wire J6oiw6, Q6oiw6, X6oiw6, E7oiw6, L7oiw6, S7oiw6, Z7oiw6, G8oiw6, N8oiw6, U8oiw6;
wire B9oiw6, I9oiw6, P9oiw6, W9oiw6, Daoiw6, Kaoiw6, Raoiw6, Yaoiw6, Fboiw6, Mboiw6;
wire Tboiw6, Acoiw6, Hcoiw6, Ocoiw6, Vcoiw6, Cdoiw6, Jdoiw6, Qdoiw6, Xdoiw6, Eeoiw6;
wire Leoiw6, Seoiw6, Zeoiw6, Gfoiw6, Nfoiw6, Ufoiw6, Bgoiw6, Igoiw6, Pgoiw6, Wgoiw6;
wire Dhoiw6, Khoiw6, Rhoiw6, Yhoiw6, Fioiw6, Mioiw6, Tioiw6, Ajoiw6, Hjoiw6, Ojoiw6;
wire Vjoiw6, Ckoiw6, Jkoiw6, Qkoiw6, Xkoiw6, Eloiw6, Lloiw6, Sloiw6, Zloiw6, Gmoiw6;
wire Nmoiw6, Umoiw6, Bnoiw6, Inoiw6, Pnoiw6, Wnoiw6, Dooiw6, Kooiw6, Rooiw6, Yooiw6;
wire Fpoiw6, Mpoiw6, Tpoiw6, Aqoiw6, Hqoiw6, Oqoiw6, Vqoiw6, Croiw6, Jroiw6, Qroiw6;
wire Xroiw6, Esoiw6, Lsoiw6, Ssoiw6, Zsoiw6, Gtoiw6, Ntoiw6, Utoiw6, Buoiw6, Iuoiw6;
wire Puoiw6, Wuoiw6, Dvoiw6, Kvoiw6, Rvoiw6, Yvoiw6, Fwoiw6, Mwoiw6, Twoiw6, Axoiw6;
wire Hxoiw6, Oxoiw6, Vxoiw6, Cyoiw6, Jyoiw6, Qyoiw6, Xyoiw6, Ezoiw6, Lzoiw6, Szoiw6;
wire Zzoiw6, G0piw6, N0piw6, U0piw6, B1piw6, I1piw6, P1piw6, W1piw6, D2piw6, K2piw6;
wire R2piw6, Y2piw6, F3piw6, M3piw6, T3piw6, A4piw6, H4piw6, O4piw6, V4piw6, C5piw6;
wire J5piw6, Q5piw6, X5piw6, E6piw6, L6piw6, S6piw6, Z6piw6, G7piw6, N7piw6, U7piw6;
wire B8piw6, I8piw6, P8piw6, W8piw6, D9piw6, K9piw6, R9piw6, Y9piw6, Fapiw6, Mapiw6;
wire Tapiw6, Abpiw6, Hbpiw6, Obpiw6, Vbpiw6, Ccpiw6, Jcpiw6, Qcpiw6, Xcpiw6, Edpiw6;
wire Ldpiw6, Sdpiw6, Zdpiw6, Gepiw6, Nepiw6, Uepiw6, Bfpiw6, Ifpiw6, Pfpiw6, Wfpiw6;
wire Dgpiw6, Kgpiw6, Rgpiw6, Ygpiw6, Fhpiw6, Mhpiw6, Thpiw6, Aipiw6, Hipiw6, Oipiw6;
wire Vipiw6, Cjpiw6, Jjpiw6, Qjpiw6, Xjpiw6, Ekpiw6, Lkpiw6, Skpiw6, Zkpiw6, Glpiw6;
wire Nlpiw6, Ulpiw6, Bmpiw6, Impiw6, Pmpiw6, Wmpiw6, Dnpiw6, Knpiw6, Rnpiw6, Ynpiw6;
wire Fopiw6, Mopiw6, Topiw6, Appiw6, Hppiw6, Oppiw6, Vppiw6, Cqpiw6, Jqpiw6, Qqpiw6;
wire Xqpiw6, Erpiw6, Lrpiw6, Srpiw6, Zrpiw6, Gspiw6, Nspiw6, Uspiw6, Btpiw6, Itpiw6;
wire Ptpiw6, Wtpiw6, Dupiw6, Kupiw6, Rupiw6, Yupiw6, Fvpiw6, Mvpiw6, Tvpiw6, Awpiw6;
wire Hwpiw6, Owpiw6, Vwpiw6, Cxpiw6, Jxpiw6, Qxpiw6, Xxpiw6, Eypiw6, Lypiw6, Sypiw6;
wire Zypiw6, Gzpiw6, Nzpiw6, Uzpiw6, B0qiw6, I0qiw6, P0qiw6, W0qiw6, D1qiw6, K1qiw6;
wire R1qiw6, Y1qiw6, F2qiw6, M2qiw6, T2qiw6, A3qiw6, H3qiw6, O3qiw6, V3qiw6, C4qiw6;
wire J4qiw6, Q4qiw6, X4qiw6, E5qiw6, L5qiw6, S5qiw6, Z5qiw6, G6qiw6, N6qiw6, U6qiw6;
wire B7qiw6, I7qiw6, P7qiw6, W7qiw6, D8qiw6, K8qiw6, R8qiw6, Y8qiw6, F9qiw6, M9qiw6;
wire T9qiw6, Aaqiw6, Haqiw6, Oaqiw6, Vaqiw6, Cbqiw6, Jbqiw6, Qbqiw6, Xbqiw6, Ecqiw6;
wire Lcqiw6, Scqiw6, Zcqiw6, Gdqiw6, Ndqiw6, Udqiw6, Beqiw6, Ieqiw6, Peqiw6, Weqiw6;
wire Dfqiw6, Kfqiw6, Rfqiw6, Yfqiw6, Fgqiw6, Mgqiw6, Tgqiw6, Ahqiw6, Hhqiw6, Ohqiw6;
wire Vhqiw6, Ciqiw6, Jiqiw6, Qiqiw6, Xiqiw6, Ejqiw6, Ljqiw6, Sjqiw6, Zjqiw6, Gkqiw6;
wire Nkqiw6, Ukqiw6, Blqiw6, Ilqiw6, Plqiw6, Wlqiw6, Dmqiw6, Kmqiw6, Rmqiw6, Ymqiw6;
wire Fnqiw6, Mnqiw6, Tnqiw6, Aoqiw6, Hoqiw6, Ooqiw6, Voqiw6, Cpqiw6, Jpqiw6, Qpqiw6;
wire Xpqiw6, Eqqiw6, Lqqiw6, Sqqiw6, Zqqiw6, Grqiw6, Nrqiw6, Urqiw6, Bsqiw6, Isqiw6;
wire Psqiw6, Wsqiw6, Dtqiw6, Ktqiw6, Rtqiw6, Ytqiw6, Fuqiw6, Muqiw6, Tuqiw6, Avqiw6;
wire Hvqiw6, Ovqiw6, Vvqiw6, Cwqiw6, Jwqiw6, Qwqiw6, Xwqiw6, Exqiw6, Lxqiw6, Sxqiw6;
wire Zxqiw6, Gyqiw6, Nyqiw6, Uyqiw6, Bzqiw6, Izqiw6, Pzqiw6, Wzqiw6, D0riw6, K0riw6;
wire R0riw6, Y0riw6, F1riw6, M1riw6, T1riw6, A2riw6, H2riw6, O2riw6, V2riw6, C3riw6;
wire J3riw6, Q3riw6, X3riw6, E4riw6, L4riw6, S4riw6, Z4riw6, G5riw6, N5riw6, U5riw6;
wire B6riw6, I6riw6, P6riw6, W6riw6, D7riw6, K7riw6, R7riw6, Y7riw6, F8riw6, M8riw6;
wire T8riw6, A9riw6, H9riw6, O9riw6, V9riw6, Cariw6, Jariw6, Qariw6, Xariw6, Ebriw6;
wire Lbriw6, Sbriw6, Zbriw6, Gcriw6, Ncriw6, Ucriw6, Bdriw6, Idriw6, Pdriw6, Wdriw6;
wire Deriw6, Keriw6, Reriw6, Yeriw6, Ffriw6, Mfriw6, Tfriw6, Agriw6, Hgriw6, Ogriw6;
wire Vgriw6, Chriw6, Jhriw6, Qhriw6, Xhriw6, Eiriw6, Liriw6, Siriw6, Ziriw6, Gjriw6;
wire Njriw6, Ujriw6, Bkriw6, Ikriw6, Pkriw6, Wkriw6, Dlriw6, Klriw6, Rlriw6, Ylriw6;
wire Fmriw6, Mmriw6, Tmriw6, Anriw6, Hnriw6, Onriw6, Vnriw6, Coriw6, Joriw6, Qoriw6;
wire Xoriw6, Epriw6, Lpriw6, Spriw6, Zpriw6, Gqriw6, Nqriw6, Uqriw6, Brriw6, Irriw6;
wire Prriw6, Wrriw6, Dsriw6, Ksriw6, Rsriw6, Ysriw6, Ftriw6, Mtriw6, Ttriw6, Auriw6;
wire Huriw6, Ouriw6, Vuriw6, Cvriw6, Jvriw6, Qvriw6, Xvriw6, Ewriw6, Lwriw6, Swriw6;
wire Zwriw6, Gxriw6, Nxriw6, Uxriw6, Byriw6, Iyriw6, Pyriw6, Wyriw6, Dzriw6, Kzriw6;
wire Rzriw6, Yzriw6, F0siw6, M0siw6, T0siw6, A1siw6, H1siw6, O1siw6, V1siw6, C2siw6;
wire J2siw6, Q2siw6, X2siw6, E3siw6, L3siw6, S3siw6, Z3siw6, G4siw6, N4siw6, U4siw6;
wire B5siw6, I5siw6, P5siw6, W5siw6, D6siw6, K6siw6, R6siw6, Y6siw6, F7siw6, M7siw6;
wire T7siw6, A8siw6, H8siw6, O8siw6, V8siw6, C9siw6, J9siw6, Q9siw6, X9siw6, Easiw6;
wire Lasiw6, Sasiw6, Zasiw6, Gbsiw6, Nbsiw6, Ubsiw6, Bcsiw6, Icsiw6, Pcsiw6, Wcsiw6;
wire Ddsiw6, Kdsiw6, Rdsiw6, Ydsiw6, Fesiw6, Mesiw6, Tesiw6, Afsiw6, Hfsiw6, Ofsiw6;
wire Vfsiw6, Cgsiw6, Jgsiw6, Qgsiw6, Xgsiw6, Ehsiw6, Lhsiw6, Shsiw6, Zhsiw6, Gisiw6;
wire Nisiw6, Uisiw6, Bjsiw6, Ijsiw6, Pjsiw6, Wjsiw6, Dksiw6, Kksiw6, Rksiw6, Yksiw6;
wire Flsiw6, Mlsiw6, Tlsiw6, Amsiw6, Hmsiw6, Omsiw6, Vmsiw6, Cnsiw6, Jnsiw6, Qnsiw6;
wire Xnsiw6, Eosiw6, Losiw6, Sosiw6, Zosiw6, Gpsiw6, Npsiw6, Upsiw6, Bqsiw6, Iqsiw6;
wire Pqsiw6, Wqsiw6, Drsiw6, Krsiw6, Rrsiw6, Yrsiw6, Fssiw6, Mssiw6, Tssiw6, Atsiw6;
wire Htsiw6, Otsiw6, Vtsiw6, Cusiw6, Jusiw6, Qusiw6, Xusiw6, Evsiw6, Lvsiw6, Svsiw6;
wire Zvsiw6, Gwsiw6, Nwsiw6, Uwsiw6, Bxsiw6, Ixsiw6, Pxsiw6, Wxsiw6, Dysiw6, Kysiw6;
wire Rysiw6, Yysiw6, Fzsiw6, Mzsiw6, Tzsiw6, A0tiw6, H0tiw6, O0tiw6, V0tiw6, C1tiw6;
wire J1tiw6, Q1tiw6, X1tiw6, E2tiw6, L2tiw6, S2tiw6, Z2tiw6, G3tiw6, N3tiw6, U3tiw6;
wire B4tiw6, I4tiw6, P4tiw6, W4tiw6, D5tiw6, K5tiw6, R5tiw6, Y5tiw6, F6tiw6, M6tiw6;
wire T6tiw6, A7tiw6, H7tiw6, O7tiw6, V7tiw6, C8tiw6, J8tiw6, Q8tiw6, X8tiw6, E9tiw6;
wire L9tiw6, S9tiw6, Z9tiw6, Gatiw6, Natiw6, Uatiw6, Bbtiw6, Ibtiw6, Pbtiw6, Wbtiw6;
wire Dctiw6, Kctiw6, Rctiw6, Yctiw6, Fdtiw6, Mdtiw6, Tdtiw6, Aetiw6, Hetiw6, Oetiw6;
wire Vetiw6, Cftiw6, Jftiw6, Qftiw6, Xftiw6, Egtiw6, Lgtiw6, Sgtiw6, Zgtiw6, Ghtiw6;
wire Nhtiw6, Uhtiw6, Bitiw6, Iitiw6, Pitiw6, Witiw6, Djtiw6, Kjtiw6, Rjtiw6, Yjtiw6;
wire Fktiw6, Mktiw6, Tktiw6, Altiw6, Hltiw6, Oltiw6, Vltiw6, Cmtiw6, Jmtiw6, Qmtiw6;
wire Xmtiw6, Entiw6, Lntiw6, Sntiw6, Zntiw6, Gotiw6, Notiw6, Uotiw6, Bptiw6, Iptiw6;
wire Pptiw6, Wptiw6, Dqtiw6, Kqtiw6, Rqtiw6, Yqtiw6, Frtiw6, Mrtiw6, Trtiw6, Astiw6;
wire Hstiw6, Ostiw6, Vstiw6, Cttiw6, Jttiw6, Qttiw6, Xttiw6, Eutiw6, Lutiw6, Sutiw6;
wire Zutiw6, Gvtiw6, Nvtiw6, Uvtiw6, Bwtiw6, Iwtiw6, Pwtiw6, Wwtiw6, Dxtiw6, Kxtiw6;
wire Rxtiw6, Yxtiw6, Fytiw6, Mytiw6, Tytiw6, Aztiw6, Hztiw6, Oztiw6, Vztiw6, C0uiw6;
wire J0uiw6, Q0uiw6, X0uiw6, E1uiw6, L1uiw6, S1uiw6, Z1uiw6, G2uiw6, N2uiw6, U2uiw6;
wire B3uiw6, I3uiw6, P3uiw6, W3uiw6, D4uiw6, K4uiw6, R4uiw6, Y4uiw6, F5uiw6, M5uiw6;
wire T5uiw6, A6uiw6, H6uiw6, O6uiw6, V6uiw6, C7uiw6, J7uiw6, Q7uiw6, X7uiw6, E8uiw6;
wire L8uiw6, S8uiw6, Z8uiw6, G9uiw6, N9uiw6, U9uiw6, Bauiw6, Iauiw6, Pauiw6, Wauiw6;
wire Dbuiw6, Kbuiw6, Rbuiw6, Ybuiw6, Fcuiw6, Mcuiw6, Tcuiw6, Aduiw6, Hduiw6, Oduiw6;
wire Vduiw6, Ceuiw6, Jeuiw6, Qeuiw6, Xeuiw6, Efuiw6, Lfuiw6, Sfuiw6, Zfuiw6, Gguiw6;
wire Nguiw6, Uguiw6, Bhuiw6, Ihuiw6, Phuiw6, Whuiw6, Diuiw6, Kiuiw6, Riuiw6, Yiuiw6;
wire Fjuiw6, Mjuiw6, Tjuiw6, Akuiw6, Hkuiw6, Okuiw6, Vkuiw6, Cluiw6, Jluiw6, Qluiw6;
wire Xluiw6, Emuiw6, Lmuiw6, Smuiw6, Zmuiw6, Gnuiw6, Nnuiw6, Unuiw6, Bouiw6, Iouiw6;
wire Pouiw6, Wouiw6, Dpuiw6, Kpuiw6, Rpuiw6, Ypuiw6, Fquiw6, Mquiw6, Tquiw6, Aruiw6;
wire Hruiw6, Oruiw6, Vruiw6, Csuiw6, Jsuiw6, Qsuiw6, Xsuiw6, Etuiw6, Ltuiw6, Stuiw6;
wire Ztuiw6, Guuiw6, Nuuiw6, Uuuiw6, Bvuiw6, Ivuiw6, Pvuiw6, Wvuiw6, Dwuiw6, Kwuiw6;
wire Rwuiw6, Ywuiw6, Fxuiw6, Mxuiw6, Txuiw6, Ayuiw6, Hyuiw6, Oyuiw6, Vyuiw6, Czuiw6;
wire Jzuiw6, Qzuiw6, Xzuiw6, E0viw6, L0viw6, S0viw6, Z0viw6, G1viw6, N1viw6, U1viw6;
wire B2viw6, I2viw6, P2viw6, W2viw6, D3viw6, K3viw6, R3viw6, Y3viw6, F4viw6, M4viw6;
wire T4viw6, A5viw6, H5viw6, O5viw6, V5viw6, C6viw6, J6viw6, Q6viw6, X6viw6, E7viw6;
wire L7viw6, S7viw6, Z7viw6, G8viw6, N8viw6, U8viw6, B9viw6, I9viw6, P9viw6, W9viw6;
wire Daviw6, Kaviw6, Raviw6, Yaviw6, Fbviw6, Mbviw6, Tbviw6, Acviw6, Hcviw6, Ocviw6;
wire Vcviw6, Cdviw6, Jdviw6, Qdviw6, Xdviw6, Eeviw6, Leviw6, Seviw6, Zeviw6, Gfviw6;
wire Nfviw6, Ufviw6, Bgviw6, Igviw6, Pgviw6, Wgviw6, Dhviw6, Khviw6, Rhviw6, Yhviw6;
wire Fiviw6, Miviw6, Tiviw6, Ajviw6, Hjviw6, Ojviw6, Vjviw6, Ckviw6, Jkviw6, Qkviw6;
wire Xkviw6, Elviw6, Llviw6, Slviw6, Zlviw6, Gmviw6, Nmviw6, Umviw6, Bnviw6, Inviw6;
wire Pnviw6, Wnviw6, Doviw6, Koviw6, Roviw6, Yoviw6, Fpviw6, Mpviw6, Tpviw6, Aqviw6;
wire Hqviw6, Oqviw6, Vqviw6, Crviw6, Jrviw6, Qrviw6, Xrviw6, Esviw6, Lsviw6, Ssviw6;
wire Zsviw6, Gtviw6, Ntviw6, Utviw6, Buviw6, Iuviw6, Puviw6, Wuviw6, Dvviw6, Kvviw6;
wire Rvviw6, Yvviw6, Fwviw6, Mwviw6, Twviw6, Axviw6, Hxviw6, Oxviw6, Vxviw6, Cyviw6;
wire Jyviw6, Qyviw6, Xyviw6, Ezviw6, Lzviw6, Szviw6, Zzviw6, G0wiw6, N0wiw6, U0wiw6;
wire B1wiw6, I1wiw6, P1wiw6, W1wiw6, D2wiw6, K2wiw6, R2wiw6, Y2wiw6, F3wiw6, M3wiw6;
wire T3wiw6, A4wiw6, H4wiw6, O4wiw6, V4wiw6, C5wiw6, J5wiw6, Q5wiw6, X5wiw6, E6wiw6;
wire L6wiw6, S6wiw6, Z6wiw6, G7wiw6, N7wiw6, U7wiw6, B8wiw6, I8wiw6, P8wiw6, W8wiw6;
wire D9wiw6, K9wiw6, R9wiw6, Y9wiw6, Fawiw6, Mawiw6, Tawiw6, Abwiw6, Hbwiw6, Obwiw6;
wire Vbwiw6, Ccwiw6, Jcwiw6, Qcwiw6, Xcwiw6, Edwiw6, Ldwiw6, Sdwiw6, Zdwiw6, Gewiw6;
wire Newiw6, Uewiw6, Bfwiw6, Ifwiw6, Pfwiw6, Wfwiw6, Dgwiw6, Kgwiw6, Rgwiw6, Ygwiw6;
wire Fhwiw6, Mhwiw6, Thwiw6, Aiwiw6, Hiwiw6, Oiwiw6, Viwiw6, Cjwiw6, Jjwiw6, Qjwiw6;
wire Xjwiw6, Ekwiw6, Lkwiw6, Skwiw6, Zkwiw6, Glwiw6, Nlwiw6, Ulwiw6, Bmwiw6, Imwiw6;
wire Pmwiw6, Wmwiw6, Dnwiw6, Knwiw6, Rnwiw6, Ynwiw6, Fowiw6, Mowiw6, Towiw6, Apwiw6;
wire Hpwiw6, Opwiw6, Vpwiw6, Cqwiw6, Jqwiw6, Qqwiw6, Xqwiw6, Erwiw6, Lrwiw6, Srwiw6;
wire Zrwiw6, Gswiw6, Nswiw6, Uswiw6, Btwiw6, Itwiw6, Ptwiw6, Wtwiw6, Duwiw6, Kuwiw6;
wire Ruwiw6, Yuwiw6, Fvwiw6, Mvwiw6, Tvwiw6, Awwiw6, Hwwiw6, Owwiw6, Vwwiw6, Cxwiw6;
wire Jxwiw6, Qxwiw6, Xxwiw6, Eywiw6, Lywiw6, Sywiw6, Zywiw6, Gzwiw6, Nzwiw6, Uzwiw6;
wire B0xiw6, I0xiw6, P0xiw6, W0xiw6, D1xiw6, K1xiw6, R1xiw6, Y1xiw6, F2xiw6, M2xiw6;
wire T2xiw6, A3xiw6, H3xiw6, O3xiw6, V3xiw6, C4xiw6, J4xiw6, Q4xiw6, X4xiw6, E5xiw6;
wire L5xiw6, S5xiw6, Z5xiw6, G6xiw6, N6xiw6, U6xiw6, B7xiw6, I7xiw6, P7xiw6, W7xiw6;
wire D8xiw6, K8xiw6, R8xiw6, Y8xiw6, F9xiw6, M9xiw6, T9xiw6, Aaxiw6, Haxiw6, Oaxiw6;
wire Vaxiw6, Cbxiw6, Jbxiw6, Qbxiw6, Xbxiw6, Ecxiw6, Lcxiw6, Scxiw6, Zcxiw6, Gdxiw6;
wire Ndxiw6, Udxiw6, Bexiw6, Iexiw6, Pexiw6, Wexiw6, Dfxiw6, Kfxiw6, Rfxiw6, Yfxiw6;
wire Fgxiw6, Mgxiw6, Tgxiw6, Ahxiw6, Hhxiw6, Ohxiw6, Vhxiw6, Cixiw6, Jixiw6, Qixiw6;
wire Xixiw6, Ejxiw6, Ljxiw6, Sjxiw6, Zjxiw6, Gkxiw6, Nkxiw6, Ukxiw6, Blxiw6, Ilxiw6;
wire Plxiw6, Wlxiw6, Dmxiw6, Kmxiw6, Rmxiw6, Ymxiw6, Fnxiw6, Mnxiw6, Tnxiw6, Aoxiw6;
wire Hoxiw6, Ooxiw6, Voxiw6, Cpxiw6, Jpxiw6, Qpxiw6, Xpxiw6, Eqxiw6, Lqxiw6, Sqxiw6;
wire Zqxiw6, Grxiw6, Nrxiw6, Urxiw6, Bsxiw6, Isxiw6, Psxiw6, Wsxiw6, Dtxiw6, Ktxiw6;
wire Rtxiw6, Ytxiw6, Fuxiw6, Muxiw6, Tuxiw6, Avxiw6, Hvxiw6, Ovxiw6, Vvxiw6, Cwxiw6;
wire Jwxiw6, Qwxiw6, Xwxiw6, Exxiw6, Lxxiw6, Sxxiw6, Zxxiw6, Gyxiw6, Nyxiw6, Uyxiw6;
wire Bzxiw6, Izxiw6, Pzxiw6, Wzxiw6, D0yiw6, K0yiw6, R0yiw6, Y0yiw6, F1yiw6, M1yiw6;
wire T1yiw6, A2yiw6, H2yiw6, O2yiw6, V2yiw6, C3yiw6, J3yiw6, Q3yiw6, X3yiw6, E4yiw6;
wire L4yiw6, S4yiw6, Z4yiw6, G5yiw6, N5yiw6, U5yiw6, B6yiw6, I6yiw6, P6yiw6, W6yiw6;
wire D7yiw6, K7yiw6, R7yiw6, Y7yiw6, F8yiw6, M8yiw6, T8yiw6, A9yiw6, H9yiw6, O9yiw6;
wire V9yiw6, Cayiw6, Jayiw6, Qayiw6, Xayiw6, Ebyiw6, Lbyiw6, Sbyiw6, Zbyiw6, Gcyiw6;
wire Ncyiw6, Ucyiw6, Bdyiw6, Idyiw6, Pdyiw6, Wdyiw6, Deyiw6, Keyiw6, Reyiw6, Yeyiw6;
wire Ffyiw6, Mfyiw6, Tfyiw6, Agyiw6, Hgyiw6, Ogyiw6, Vgyiw6, Chyiw6, Jhyiw6, Qhyiw6;
wire Xhyiw6, Eiyiw6, Liyiw6, Siyiw6, Ziyiw6, Gjyiw6, Njyiw6, Ujyiw6, Bkyiw6, Ikyiw6;
wire Pkyiw6, Wkyiw6, Dlyiw6, Klyiw6, Rlyiw6, Ylyiw6, Fmyiw6, Mmyiw6, Tmyiw6, Anyiw6;
wire Hnyiw6, Onyiw6, Vnyiw6, Coyiw6, Joyiw6, Qoyiw6, Xoyiw6, Epyiw6, Lpyiw6, Spyiw6;
wire Zpyiw6, Gqyiw6, Nqyiw6, Uqyiw6, Bryiw6, Iryiw6, Pryiw6, Wryiw6, Dsyiw6, Ksyiw6;
wire Rsyiw6, Ysyiw6, Ftyiw6, Mtyiw6, Ttyiw6, Auyiw6, Huyiw6, Ouyiw6, Vuyiw6, Cvyiw6;
wire Jvyiw6, Qvyiw6, Xvyiw6, Ewyiw6, Lwyiw6, Swyiw6, Zwyiw6, Gxyiw6, Nxyiw6, Uxyiw6;
wire Byyiw6, Iyyiw6, Pyyiw6, Wyyiw6, Dzyiw6, Kzyiw6, Rzyiw6, Yzyiw6, F0ziw6, M0ziw6;
wire T0ziw6, A1ziw6, H1ziw6, O1ziw6, V1ziw6, C2ziw6, J2ziw6, Q2ziw6, X2ziw6, E3ziw6;
wire L3ziw6, S3ziw6, Z3ziw6, G4ziw6, N4ziw6, U4ziw6, B5ziw6, I5ziw6, P5ziw6, W5ziw6;
wire D6ziw6, K6ziw6, R6ziw6, Y6ziw6, F7ziw6, M7ziw6, T7ziw6, A8ziw6, H8ziw6, O8ziw6;
wire V8ziw6, C9ziw6, J9ziw6, Q9ziw6, X9ziw6, Eaziw6, Laziw6, Saziw6, Zaziw6, Gbziw6;
wire Nbziw6, Ubziw6, Bcziw6, Icziw6, Pcziw6, Wcziw6, Ddziw6, Kdziw6, Rdziw6, Ydziw6;
wire Feziw6, Meziw6, Teziw6, Afziw6, Hfziw6, Ofziw6, Vfziw6, Cgziw6, Jgziw6, Qgziw6;
wire Xgziw6, Ehziw6, Lhziw6, Shziw6, Zhziw6, Giziw6, Niziw6, Uiziw6, Bjziw6, Ijziw6;
wire Pjziw6, Wjziw6, Dkziw6, Kkziw6, Rkziw6, Ykziw6, Flziw6, Mlziw6, Tlziw6, Amziw6;
wire Hmziw6, Omziw6, Vmziw6, Cnziw6, Jnziw6, Qnziw6, Xnziw6, Eoziw6, Loziw6, Soziw6;
wire Zoziw6, Gpziw6, Npziw6, Upziw6, Bqziw6, Iqziw6, Pqziw6, Wqziw6, Drziw6, Krziw6;
wire Rrziw6, Yrziw6, Fsziw6, Msziw6, Tsziw6, Atziw6, Htziw6, Otziw6, Vtziw6, Cuziw6;
wire Juziw6, Quziw6, Xuziw6, Evziw6, Lvziw6, Svziw6, Zvziw6, Gwziw6, Nwziw6, Uwziw6;
wire Bxziw6, Ixziw6, Pxziw6, Wxziw6, Dyziw6, Kyziw6, Ryziw6, Yyziw6, Fzziw6, Mzziw6;
wire Tzziw6, A00jw6, H00jw6, O00jw6, V00jw6, C10jw6, J10jw6, Q10jw6, X10jw6, E20jw6;
wire L20jw6, S20jw6, Z20jw6, G30jw6, N30jw6, U30jw6, B40jw6, I40jw6, P40jw6, W40jw6;
wire D50jw6, K50jw6, R50jw6, Y50jw6, F60jw6, M60jw6, T60jw6, A70jw6, H70jw6, O70jw6;
wire V70jw6, C80jw6, J80jw6, Q80jw6, X80jw6, E90jw6, L90jw6, S90jw6, Z90jw6, Ga0jw6;
wire Na0jw6, Ua0jw6, Bb0jw6, Ib0jw6, Pb0jw6, Wb0jw6, Dc0jw6, Kc0jw6, Rc0jw6, Yc0jw6;
wire Fd0jw6, Md0jw6, Td0jw6, Ae0jw6, He0jw6, Oe0jw6, Ve0jw6, Cf0jw6, Jf0jw6, Qf0jw6;
wire Xf0jw6, Eg0jw6, Lg0jw6, Sg0jw6, Zg0jw6, Gh0jw6, Nh0jw6, Uh0jw6, Bi0jw6, Ii0jw6;
wire Pi0jw6, Wi0jw6, Dj0jw6, Kj0jw6, Rj0jw6, Yj0jw6, Fk0jw6, Mk0jw6, Tk0jw6, Al0jw6;
wire Hl0jw6, Ol0jw6, Vl0jw6, Cm0jw6, Jm0jw6, Qm0jw6, Xm0jw6, En0jw6, Ln0jw6, Sn0jw6;
wire Zn0jw6, Go0jw6, No0jw6, Uo0jw6, Bp0jw6, Ip0jw6, Pp0jw6, Wp0jw6, Dq0jw6, Kq0jw6;
wire Rq0jw6, Yq0jw6, Fr0jw6, Mr0jw6, Tr0jw6, As0jw6, Hs0jw6, Os0jw6, Vs0jw6, Ct0jw6;
wire Jt0jw6, Qt0jw6, Xt0jw6, Eu0jw6, Lu0jw6, Su0jw6, Zu0jw6, Gv0jw6, Nv0jw6, Uv0jw6;
wire Bw0jw6, Iw0jw6, Pw0jw6, Ww0jw6, Dx0jw6, Kx0jw6, Rx0jw6, Yx0jw6, Fy0jw6, My0jw6;
wire Ty0jw6, Az0jw6, Hz0jw6, Oz0jw6, Vz0jw6, C01jw6, J01jw6, Q01jw6, X01jw6, E11jw6;
wire L11jw6, S11jw6, Z11jw6, G21jw6, N21jw6, U21jw6, B31jw6, I31jw6, P31jw6, W31jw6;
wire D41jw6, K41jw6, R41jw6, Y41jw6, F51jw6, M51jw6, T51jw6, A61jw6, H61jw6, O61jw6;
wire V61jw6, C71jw6, J71jw6, Q71jw6, X71jw6, E81jw6, L81jw6, S81jw6, Z81jw6, G91jw6;
wire N91jw6, U91jw6, Ba1jw6, Ia1jw6, Pa1jw6, Wa1jw6, Db1jw6, Kb1jw6, Rb1jw6, Yb1jw6;
wire Fc1jw6, Mc1jw6, Tc1jw6, Ad1jw6, Hd1jw6, Od1jw6, Vd1jw6, Ce1jw6, Je1jw6, Qe1jw6;
wire Xe1jw6, Ef1jw6, Lf1jw6, Sf1jw6, Zf1jw6, Gg1jw6, Ng1jw6, Ug1jw6, Bh1jw6, Ih1jw6;
wire Ph1jw6, Wh1jw6, Di1jw6, Ki1jw6, Ri1jw6, Yi1jw6, Fj1jw6, Mj1jw6, Tj1jw6, Ak1jw6;
wire Hk1jw6, Ok1jw6, Vk1jw6, Cl1jw6, Jl1jw6, Ql1jw6, Xl1jw6, Em1jw6, Lm1jw6, Sm1jw6;
wire Zm1jw6, Gn1jw6, Nn1jw6, Un1jw6, Bo1jw6, Io1jw6, Po1jw6, Wo1jw6, Dp1jw6, Kp1jw6;
wire Rp1jw6, Yp1jw6, Fq1jw6, Mq1jw6, Tq1jw6, Ar1jw6, Hr1jw6, Or1jw6, Vr1jw6, Cs1jw6;
wire Js1jw6, Qs1jw6, Xs1jw6, Et1jw6, Lt1jw6, St1jw6, Zt1jw6, Gu1jw6, Nu1jw6, Uu1jw6;
wire Bv1jw6, Iv1jw6, Pv1jw6, Wv1jw6, Dw1jw6, Kw1jw6, Rw1jw6, Yw1jw6, Fx1jw6, Mx1jw6;
wire Tx1jw6, Ay1jw6, Hy1jw6, Oy1jw6, Vy1jw6, Cz1jw6, Jz1jw6, Qz1jw6, Xz1jw6, E02jw6;
wire L02jw6, S02jw6, Z02jw6, G12jw6, N12jw6, U12jw6, B22jw6, I22jw6, P22jw6, W22jw6;
wire D32jw6, K32jw6, R32jw6, Y32jw6, F42jw6, M42jw6, T42jw6, A52jw6, H52jw6, O52jw6;
wire V52jw6, C62jw6, J62jw6, Q62jw6, X62jw6, E72jw6, L72jw6, S72jw6, Z72jw6, G82jw6;
wire N82jw6, U82jw6, B92jw6, I92jw6, P92jw6, W92jw6, Da2jw6, Ka2jw6, Ra2jw6, Ya2jw6;
wire Fb2jw6, Mb2jw6, Tb2jw6, Ac2jw6, Hc2jw6, Oc2jw6, Vc2jw6, Cd2jw6, Jd2jw6, Qd2jw6;
wire Xd2jw6, Ee2jw6, Le2jw6, Se2jw6, Ze2jw6, Gf2jw6, Nf2jw6, Uf2jw6, Bg2jw6, Ig2jw6;
wire Pg2jw6, Wg2jw6, Dh2jw6, Kh2jw6, Rh2jw6, Yh2jw6, Fi2jw6, Mi2jw6, Ti2jw6, Aj2jw6;
wire Hj2jw6, Oj2jw6, Vj2jw6, Ck2jw6, Jk2jw6, Qk2jw6, Xk2jw6, El2jw6, Ll2jw6, Sl2jw6;
wire Zl2jw6, Gm2jw6, Nm2jw6, Um2jw6, Bn2jw6, In2jw6, Pn2jw6, Wn2jw6, Do2jw6, Ko2jw6;
wire Ro2jw6, Yo2jw6, Fp2jw6, Mp2jw6, Tp2jw6, Aq2jw6, Hq2jw6, Oq2jw6, Vq2jw6, Cr2jw6;
wire Jr2jw6, Qr2jw6, Xr2jw6, Es2jw6, Ls2jw6, Ss2jw6, Zs2jw6, Gt2jw6, Nt2jw6, Ut2jw6;
wire Bu2jw6, Iu2jw6, Pu2jw6, Wu2jw6, Dv2jw6, Kv2jw6, Rv2jw6, Yv2jw6, Fw2jw6, Mw2jw6;
wire Tw2jw6, Ax2jw6, Hx2jw6, Ox2jw6, Vx2jw6, Cy2jw6, Jy2jw6, Qy2jw6, Xy2jw6, Ez2jw6;
wire Lz2jw6, Sz2jw6, Zz2jw6, G03jw6, N03jw6, U03jw6, B13jw6, I13jw6, P13jw6, W13jw6;
wire D23jw6, K23jw6, R23jw6, Y23jw6, F33jw6, M33jw6, T33jw6, A43jw6, H43jw6, O43jw6;
wire V43jw6, C53jw6, J53jw6, Q53jw6, X53jw6, E63jw6, L63jw6, S63jw6, Z63jw6, G73jw6;
wire N73jw6, U73jw6, B83jw6, I83jw6, P83jw6, W83jw6, D93jw6, K93jw6, R93jw6, Y93jw6;
wire Fa3jw6, Ma3jw6, Ta3jw6, Ab3jw6, Hb3jw6, Ob3jw6, Vb3jw6, Cc3jw6, Jc3jw6, Qc3jw6;
wire Xc3jw6, Ed3jw6, Ld3jw6, Sd3jw6, Zd3jw6, Ge3jw6, Ne3jw6, Ue3jw6, Bf3jw6, If3jw6;
wire Pf3jw6, Wf3jw6, Dg3jw6, Kg3jw6, Rg3jw6, Yg3jw6, Fh3jw6, Mh3jw6, Th3jw6, Ai3jw6;
wire Hi3jw6, Oi3jw6, Vi3jw6, Cj3jw6, Jj3jw6, Qj3jw6, Xj3jw6, Ek3jw6, Lk3jw6, Sk3jw6;
wire Zk3jw6, Gl3jw6, Nl3jw6, Ul3jw6, Bm3jw6, Im3jw6, Pm3jw6, Wm3jw6, Dn3jw6, Kn3jw6;
wire Rn3jw6, Yn3jw6, Fo3jw6, Mo3jw6, To3jw6, Ap3jw6, Hp3jw6, Op3jw6, Vp3jw6, Cq3jw6;
wire Jq3jw6, Qq3jw6, Xq3jw6, Er3jw6, Lr3jw6, Sr3jw6, Zr3jw6, Gs3jw6, Ns3jw6, Us3jw6;
wire Bt3jw6, It3jw6, Pt3jw6, Wt3jw6, Du3jw6, Ku3jw6, Ru3jw6, Yu3jw6, Fv3jw6, Mv3jw6;
wire Tv3jw6, Aw3jw6, Hw3jw6, Ow3jw6, Vw3jw6, Cx3jw6, Jx3jw6, Qx3jw6, Xx3jw6, Ey3jw6;
wire Ly3jw6, Sy3jw6, Zy3jw6, Gz3jw6, Nz3jw6, Uz3jw6, B04jw6, I04jw6, P04jw6, W04jw6;
wire D14jw6, K14jw6, R14jw6, Y14jw6, F24jw6, M24jw6, T24jw6, A34jw6, H34jw6, O34jw6;
wire V34jw6, C44jw6, J44jw6, Q44jw6, X44jw6, E54jw6, L54jw6, S54jw6, Z54jw6, G64jw6;
wire N64jw6, U64jw6, B74jw6, I74jw6, P74jw6, W74jw6, D84jw6, K84jw6, R84jw6, Y84jw6;
wire F94jw6, M94jw6, T94jw6, Aa4jw6, Ha4jw6, Oa4jw6, Va4jw6, Cb4jw6, Jb4jw6, Qb4jw6;
wire Xb4jw6, Ec4jw6, Lc4jw6, Sc4jw6, Zc4jw6, Gd4jw6, Nd4jw6, Ud4jw6, Be4jw6, Ie4jw6;
wire Pe4jw6, We4jw6, Df4jw6, Kf4jw6, Rf4jw6, Yf4jw6, Fg4jw6, Mg4jw6, Tg4jw6, Ah4jw6;
wire Hh4jw6, Oh4jw6, Vh4jw6, Ci4jw6, Ji4jw6, Qi4jw6, Xi4jw6, Ej4jw6, Lj4jw6, Sj4jw6;
wire Zj4jw6, Gk4jw6, Nk4jw6, Uk4jw6, Bl4jw6, Il4jw6, Pl4jw6, Wl4jw6, Dm4jw6, Km4jw6;
wire Rm4jw6, Ym4jw6, Fn4jw6, Mn4jw6, Tn4jw6, Ao4jw6, Ho4jw6, Oo4jw6, Vo4jw6, Cp4jw6;
wire Jp4jw6, Qp4jw6, Xp4jw6, Eq4jw6, Lq4jw6, Sq4jw6, Zq4jw6, Gr4jw6, Nr4jw6, Ur4jw6;
wire Bs4jw6, Is4jw6, Ps4jw6, Ws4jw6, Dt4jw6, Kt4jw6, Rt4jw6, Yt4jw6, Fu4jw6, Mu4jw6;
wire Tu4jw6, Av4jw6, Hv4jw6, Ov4jw6, Vv4jw6, Cw4jw6, Jw4jw6, Qw4jw6, Xw4jw6, Ex4jw6;
wire Lx4jw6, Sx4jw6, Zx4jw6, Gy4jw6, Ny4jw6, Uy4jw6, Bz4jw6, Iz4jw6, Pz4jw6, Wz4jw6;
wire D05jw6, K05jw6, R05jw6, Y05jw6, F15jw6, M15jw6, T15jw6, A25jw6, H25jw6, O25jw6;
wire V25jw6, C35jw6, J35jw6, Q35jw6, X35jw6, E45jw6, L45jw6, S45jw6, Z45jw6, G55jw6;
wire N55jw6, U55jw6, B65jw6, I65jw6, P65jw6, W65jw6, D75jw6, K75jw6, R75jw6, Y75jw6;
wire F85jw6, M85jw6, T85jw6, A95jw6, H95jw6, O95jw6, V95jw6, Ca5jw6, Ja5jw6, Qa5jw6;
wire Xa5jw6, Eb5jw6, Lb5jw6, Sb5jw6, Zb5jw6, Gc5jw6, Nc5jw6, Uc5jw6, Bd5jw6, Id5jw6;
wire Pd5jw6, Wd5jw6, De5jw6, Ke5jw6, Re5jw6, Ye5jw6, Ff5jw6, Mf5jw6, Tf5jw6, Ag5jw6;
wire Hg5jw6, Og5jw6, Vg5jw6, Ch5jw6, Jh5jw6, Qh5jw6, Xh5jw6, Ei5jw6, Li5jw6, Si5jw6;
wire Zi5jw6, Gj5jw6, Nj5jw6, Uj5jw6, Bk5jw6, Ik5jw6, Pk5jw6, Wk5jw6, Dl5jw6, Kl5jw6;
wire Rl5jw6, Yl5jw6, Fm5jw6, Mm5jw6, Tm5jw6, An5jw6, Hn5jw6, On5jw6, Vn5jw6, Co5jw6;
wire Jo5jw6, Qo5jw6, Xo5jw6, Ep5jw6, Lp5jw6, Sp5jw6, Zp5jw6, Gq5jw6, Nq5jw6, Uq5jw6;
wire Br5jw6, Ir5jw6, Pr5jw6, Wr5jw6, Ds5jw6, Ks5jw6, Rs5jw6, Ys5jw6, Ft5jw6, Mt5jw6;
wire Tt5jw6, Au5jw6, Hu5jw6, Ou5jw6, Vu5jw6, Cv5jw6, Jv5jw6, Qv5jw6, Xv5jw6, Ew5jw6;
wire Lw5jw6, Sw5jw6, Zw5jw6, Gx5jw6, Nx5jw6, Ux5jw6, By5jw6, Iy5jw6, Py5jw6, Wy5jw6;
wire Dz5jw6, Kz5jw6, Rz5jw6, Yz5jw6, F06jw6, M06jw6, T06jw6, A16jw6, H16jw6, O16jw6;
wire V16jw6, C26jw6, J26jw6, Q26jw6, X26jw6, E36jw6, L36jw6, S36jw6, Z36jw6, G46jw6;
wire N46jw6, U46jw6, B56jw6, I56jw6, P56jw6, W56jw6, D66jw6, K66jw6, R66jw6, Y66jw6;
wire F76jw6, M76jw6, T76jw6, A86jw6, H86jw6, O86jw6, V86jw6, C96jw6, J96jw6, Q96jw6;
wire X96jw6, Ea6jw6, La6jw6, Sa6jw6, Za6jw6, Gb6jw6, Nb6jw6, Ub6jw6, Bc6jw6, Ic6jw6;
wire Pc6jw6, Wc6jw6, Dd6jw6, Kd6jw6, Rd6jw6, Yd6jw6, Fe6jw6, Me6jw6, Te6jw6, Af6jw6;
wire Hf6jw6, Of6jw6, Vf6jw6, Cg6jw6, Jg6jw6, Qg6jw6, Xg6jw6, Eh6jw6, Lh6jw6, Sh6jw6;
wire Zh6jw6, Gi6jw6, Ni6jw6, Ui6jw6, Bj6jw6, Ij6jw6, Pj6jw6, Wj6jw6, Dk6jw6, Kk6jw6;
wire Rk6jw6, Yk6jw6, Fl6jw6, Ml6jw6, Tl6jw6, Am6jw6, Hm6jw6, Om6jw6, Vm6jw6, Cn6jw6;
wire Jn6jw6, Qn6jw6, Xn6jw6, Eo6jw6, Lo6jw6, So6jw6, Zo6jw6, Gp6jw6, Np6jw6, Up6jw6;
wire Bq6jw6, Iq6jw6, Pq6jw6, Wq6jw6, Dr6jw6, Kr6jw6, Rr6jw6, Yr6jw6, Fs6jw6, Ms6jw6;
wire Ts6jw6, At6jw6, Ht6jw6, Ot6jw6, Vt6jw6, Cu6jw6, Ju6jw6, Qu6jw6, Xu6jw6, Ev6jw6;
wire Lv6jw6, Sv6jw6, Zv6jw6, Gw6jw6, Nw6jw6, Uw6jw6, Bx6jw6, Ix6jw6, Px6jw6, Wx6jw6;
wire Dy6jw6, Ky6jw6, Ry6jw6, Yy6jw6, Fz6jw6, Mz6jw6, Tz6jw6, A07jw6, H07jw6, O07jw6;
wire V07jw6, C17jw6, J17jw6, Q17jw6, X17jw6, E27jw6, L27jw6, S27jw6, Z27jw6, G37jw6;
wire N37jw6, U37jw6, B47jw6, I47jw6, P47jw6, W47jw6, D57jw6, K57jw6, R57jw6, Y57jw6;
wire F67jw6, M67jw6, T67jw6, A77jw6, H77jw6, O77jw6, V77jw6, C87jw6, J87jw6, Q87jw6;
wire X87jw6, E97jw6, L97jw6, S97jw6, Z97jw6, Ga7jw6, Na7jw6, Ua7jw6, Bb7jw6, Ib7jw6;
wire Pb7jw6, Wb7jw6, Dc7jw6, Kc7jw6, Rc7jw6, Yc7jw6, Fd7jw6, Md7jw6, Td7jw6, Ae7jw6;
wire He7jw6, Oe7jw6, Ve7jw6, Cf7jw6, Jf7jw6, Qf7jw6, Xf7jw6, Eg7jw6, Lg7jw6, Sg7jw6;
wire Zg7jw6, Gh7jw6, Nh7jw6, Uh7jw6, Bi7jw6, Ii7jw6, Pi7jw6, Wi7jw6, Dj7jw6, Kj7jw6;
wire Rj7jw6, Yj7jw6, Fk7jw6, Mk7jw6, Tk7jw6, Al7jw6, Hl7jw6, Ol7jw6, Vl7jw6, Cm7jw6;
wire Jm7jw6, Qm7jw6, Xm7jw6, En7jw6, Ln7jw6, Sn7jw6, Zn7jw6, Go7jw6, No7jw6, Uo7jw6;
wire Bp7jw6, Ip7jw6, Pp7jw6, Wp7jw6, Dq7jw6, Kq7jw6, Rq7jw6, Yq7jw6, Fr7jw6, Mr7jw6;
wire Tr7jw6, As7jw6, Hs7jw6, Os7jw6, Vs7jw6, Ct7jw6, Jt7jw6, Qt7jw6, Xt7jw6, Eu7jw6;
wire Lu7jw6, Su7jw6, Zu7jw6, Gv7jw6, Nv7jw6, Uv7jw6, Bw7jw6, Iw7jw6, Pw7jw6, Ww7jw6;
wire Dx7jw6, Kx7jw6, Rx7jw6, Yx7jw6, Fy7jw6, My7jw6, Ty7jw6, Az7jw6, Hz7jw6, Oz7jw6;
wire Vz7jw6, C08jw6, J08jw6, Q08jw6, X08jw6, E18jw6, L18jw6, S18jw6, Z18jw6, G28jw6;
wire N28jw6, U28jw6, B38jw6, I38jw6, P38jw6, W38jw6, D48jw6, K48jw6, R48jw6, Y48jw6;
wire F58jw6, M58jw6, T58jw6, A68jw6, H68jw6, O68jw6, V68jw6, C78jw6, J78jw6, Q78jw6;
wire X78jw6, E88jw6, L88jw6, S88jw6, Z88jw6, G98jw6, N98jw6, U98jw6, Ba8jw6, Ia8jw6;
wire Pa8jw6, Wa8jw6, Db8jw6, Kb8jw6, Rb8jw6, Yb8jw6, Fc8jw6, Mc8jw6, Tc8jw6, Ad8jw6;
wire Hd8jw6, Od8jw6, Vd8jw6, Ce8jw6, Je8jw6, Qe8jw6, Xe8jw6, Ef8jw6, Lf8jw6, Sf8jw6;
wire Zf8jw6, Gg8jw6, Ng8jw6, Ug8jw6, Bh8jw6, Ih8jw6, Ph8jw6, Wh8jw6, Di8jw6, Ki8jw6;
wire Ri8jw6, Yi8jw6, Fj8jw6, Mj8jw6, Tj8jw6, Ak8jw6, Hk8jw6, Ok8jw6, Vk8jw6, Cl8jw6;
wire Jl8jw6, Ql8jw6, Xl8jw6, Em8jw6, Lm8jw6, Sm8jw6, Zm8jw6, Gn8jw6, Nn8jw6, Un8jw6;
wire Bo8jw6, Io8jw6, Po8jw6, Wo8jw6, Dp8jw6, Kp8jw6, Rp8jw6, Yp8jw6, Fq8jw6, Mq8jw6;
wire Tq8jw6, Ar8jw6, Hr8jw6, Or8jw6, Vr8jw6, Cs8jw6, Js8jw6, Qs8jw6, Xs8jw6, Et8jw6;
wire Lt8jw6, St8jw6, Zt8jw6, Gu8jw6, Nu8jw6, Uu8jw6, Bv8jw6, Iv8jw6, Pv8jw6, Wv8jw6;
wire Dw8jw6, Kw8jw6, Rw8jw6, Yw8jw6, Fx8jw6, Mx8jw6, Tx8jw6, Ay8jw6, Hy8jw6, Oy8jw6;
wire Vy8jw6, Cz8jw6, Jz8jw6, Qz8jw6, Xz8jw6, E09jw6, L09jw6, S09jw6, Z09jw6, G19jw6;
wire N19jw6, U19jw6, B29jw6, I29jw6, P29jw6, W29jw6, D39jw6, K39jw6, R39jw6, Y39jw6;
wire F49jw6, M49jw6, T49jw6, A59jw6, H59jw6, O59jw6, V59jw6, C69jw6, J69jw6, Q69jw6;
wire X69jw6, E79jw6, L79jw6, S79jw6, Z79jw6, G89jw6, N89jw6, U89jw6, B99jw6, I99jw6;
wire P99jw6, W99jw6, Da9jw6, Ka9jw6, Ra9jw6, Ya9jw6, Fb9jw6, Mb9jw6, Tb9jw6, Ac9jw6;
wire Hc9jw6, Oc9jw6, Vc9jw6, Cd9jw6, Jd9jw6, Qd9jw6, Xd9jw6, Ee9jw6, Le9jw6, Se9jw6;
wire Ze9jw6, Gf9jw6, Nf9jw6, Uf9jw6, Bg9jw6, Ig9jw6, Pg9jw6, Wg9jw6, Dh9jw6, Kh9jw6;
wire Rh9jw6, Yh9jw6, Fi9jw6, Mi9jw6, Ti9jw6, Aj9jw6, Hj9jw6, Oj9jw6, Vj9jw6, Ck9jw6;
wire Jk9jw6, Qk9jw6, Xk9jw6, El9jw6, Ll9jw6, Sl9jw6, Zl9jw6, Gm9jw6, Nm9jw6, Um9jw6;
wire Bn9jw6, In9jw6, Pn9jw6, Wn9jw6, Do9jw6, Ko9jw6, Ro9jw6, Yo9jw6, Fp9jw6, Mp9jw6;
wire Tp9jw6, Aq9jw6, Hq9jw6, Oq9jw6, Vq9jw6, Cr9jw6, Jr9jw6, Qr9jw6, Xr9jw6, Es9jw6;
wire Ls9jw6, Ss9jw6, Zs9jw6, Gt9jw6, Nt9jw6, Ut9jw6, Bu9jw6, Iu9jw6, Pu9jw6, Wu9jw6;
wire Dv9jw6, Kv9jw6, Rv9jw6, Yv9jw6, Fw9jw6, Mw9jw6, Tw9jw6, Ax9jw6, Hx9jw6, Ox9jw6;
wire Vx9jw6, Cy9jw6, Jy9jw6, Qy9jw6, Xy9jw6, Ez9jw6, Lz9jw6, Sz9jw6, Zz9jw6, G0ajw6;
wire N0ajw6, U0ajw6, B1ajw6, I1ajw6, P1ajw6, W1ajw6, D2ajw6, K2ajw6, R2ajw6, Y2ajw6;
wire F3ajw6, M3ajw6, T3ajw6, A4ajw6, H4ajw6, O4ajw6, V4ajw6, C5ajw6, J5ajw6, Q5ajw6;
wire X5ajw6, E6ajw6, L6ajw6, S6ajw6, Z6ajw6, G7ajw6, N7ajw6, U7ajw6, B8ajw6, I8ajw6;
wire P8ajw6, W8ajw6, D9ajw6, K9ajw6, R9ajw6, Y9ajw6, Faajw6, Maajw6, Taajw6, Abajw6;
wire Hbajw6, Obajw6, Vbajw6, Ccajw6, Jcajw6, Qcajw6, Xcajw6, Edajw6, Ldajw6, Sdajw6;
wire Zdajw6, Geajw6, Neajw6, Ueajw6, Bfajw6, Ifajw6, Pfajw6, Wfajw6, Dgajw6, Kgajw6;
wire Rgajw6, Ygajw6, Fhajw6, Mhajw6, Thajw6, Aiajw6, Hiajw6, Oiajw6, Viajw6, Cjajw6;
wire Jjajw6, Qjajw6, Xjajw6, Ekajw6, Lkajw6, Skajw6, Zkajw6, Glajw6, Nlajw6, Ulajw6;
wire Bmajw6, Imajw6, Pmajw6, Wmajw6, Dnajw6, Knajw6, Rnajw6, Ynajw6, Foajw6, Moajw6;
wire Toajw6, Apajw6, Hpajw6, Opajw6, Vpajw6, Cqajw6, Jqajw6, Qqajw6, Xqajw6, Erajw6;
wire Lrajw6, Srajw6, Zrajw6, Gsajw6, Nsajw6, Usajw6, Btajw6, Itajw6, Ptajw6, Wtajw6;
wire Duajw6, Kuajw6, Ruajw6, Yuajw6, Fvajw6, Mvajw6, Tvajw6, Awajw6, Hwajw6, Owajw6;
wire Vwajw6, Cxajw6, Jxajw6, Qxajw6, Xxajw6, Eyajw6, Lyajw6, Syajw6, Zyajw6, Gzajw6;
wire Nzajw6, Uzajw6, B0bjw6, I0bjw6, P0bjw6, W0bjw6, D1bjw6, K1bjw6, R1bjw6, Y1bjw6;
wire F2bjw6, M2bjw6, T2bjw6, A3bjw6, H3bjw6, O3bjw6, V3bjw6, C4bjw6, J4bjw6, Q4bjw6;
wire X4bjw6, E5bjw6, L5bjw6, S5bjw6, Z5bjw6, G6bjw6, N6bjw6, U6bjw6, B7bjw6, I7bjw6;
wire P7bjw6, W7bjw6, D8bjw6, K8bjw6, R8bjw6, Y8bjw6, F9bjw6, M9bjw6, T9bjw6, Aabjw6;
wire Habjw6, Oabjw6, Vabjw6, Cbbjw6, Jbbjw6, Qbbjw6, Xbbjw6, Ecbjw6, Lcbjw6, Scbjw6;
wire Zcbjw6, Gdbjw6, Ndbjw6, Udbjw6, Bebjw6, Iebjw6, Pebjw6, Webjw6, Dfbjw6, Kfbjw6;
wire Rfbjw6, Yfbjw6, Fgbjw6, Mgbjw6, Tgbjw6, Ahbjw6, Hhbjw6, Ohbjw6, Vhbjw6, Cibjw6;
wire Jibjw6, Qibjw6, Xibjw6, Ejbjw6, Ljbjw6, Sjbjw6, Zjbjw6, Gkbjw6, Nkbjw6, Ukbjw6;
wire Blbjw6, Ilbjw6, Plbjw6, Wlbjw6, Dmbjw6, Kmbjw6, Rmbjw6, Ymbjw6, Fnbjw6, Mnbjw6;
wire Tnbjw6, Aobjw6, Hobjw6, Oobjw6, Vobjw6, Cpbjw6, Jpbjw6, Qpbjw6, Xpbjw6, Eqbjw6;
wire Lqbjw6, Sqbjw6, Zqbjw6, Grbjw6, Nrbjw6, Urbjw6, Bsbjw6, Isbjw6, Psbjw6, Wsbjw6;
wire Dtbjw6, Ktbjw6, Rtbjw6, Ytbjw6, Fubjw6, Mubjw6, Tubjw6, Avbjw6, Hvbjw6, Ovbjw6;
wire Vvbjw6, Cwbjw6, Jwbjw6, Qwbjw6, Xwbjw6, Exbjw6, Lxbjw6, Sxbjw6, Zxbjw6, Gybjw6;
wire Nybjw6, Uybjw6, Bzbjw6, Izbjw6, Pzbjw6, Wzbjw6, D0cjw6, K0cjw6, R0cjw6, Y0cjw6;
wire F1cjw6, M1cjw6, T1cjw6, A2cjw6, H2cjw6, O2cjw6, V2cjw6, C3cjw6, J3cjw6, Q3cjw6;
wire X3cjw6, E4cjw6, L4cjw6, S4cjw6, Z4cjw6, G5cjw6, N5cjw6, U5cjw6, B6cjw6, I6cjw6;
wire P6cjw6, W6cjw6, D7cjw6, K7cjw6, R7cjw6, Y7cjw6, F8cjw6, M8cjw6, T8cjw6, A9cjw6;
wire H9cjw6, O9cjw6, V9cjw6, Cacjw6, Jacjw6, Qacjw6, Xacjw6, Ebcjw6, Lbcjw6, Sbcjw6;
wire Zbcjw6, Gccjw6, Nccjw6, Uccjw6, Bdcjw6, Idcjw6, Pdcjw6, Wdcjw6, Decjw6, Kecjw6;
wire Recjw6, Yecjw6, Ffcjw6, Mfcjw6, Tfcjw6, Agcjw6, Hgcjw6, Ogcjw6, Vgcjw6, Chcjw6;
wire Jhcjw6, Qhcjw6, Xhcjw6, Eicjw6, Licjw6, Sicjw6, Zicjw6, Gjcjw6, Njcjw6, Ujcjw6;
wire Bkcjw6, Ikcjw6, Pkcjw6, Wkcjw6, Dlcjw6, Klcjw6, Rlcjw6, Ylcjw6, Fmcjw6, Mmcjw6;
wire Tmcjw6, Ikg6x6, Pkg6x6, Wkg6x6, Dlg6x6, Klg6x6, Rlg6x6, Ylg6x6, Fmg6x6, Mmg6x6;
wire Tmg6x6, Ang6x6, Hng6x6, Ong6x6, Vng6x6, Cog6x6, Jog6x6, Qog6x6, Xog6x6, Epg6x6;
wire Lpg6x6, Spg6x6, Zpg6x6, Gqg6x6, Nqg6x6, Uqg6x6, Brg6x6, Irg6x6, Prg6x6, Wrg6x6;
wire Dsg6x6, Ksg6x6, Rsg6x6, Ysg6x6, Ftg6x6, Mtg6x6, Ttg6x6, Aug6x6, Hug6x6, Oug6x6;
wire Vug6x6, Cvg6x6, Jvg6x6, Qvg6x6, Xvg6x6, Ewg6x6, Lwg6x6, Swg6x6, Zwg6x6, Gxg6x6;
wire Nxg6x6, Uxg6x6, Byg6x6, Iyg6x6, Pyg6x6, Wyg6x6, Dzg6x6, Kzg6x6, Rzg6x6, Yzg6x6;
wire F0h6x6, M0h6x6, T0h6x6, A1h6x6, H1h6x6, O1h6x6, V1h6x6, C2h6x6, J2h6x6, Q2h6x6;
wire X2h6x6, E3h6x6, L3h6x6, S3h6x6, Z3h6x6, G4h6x6, N4h6x6, U4h6x6, B5h6x6, I5h6x6;
wire P5h6x6, W5h6x6, D6h6x6, K6h6x6, R6h6x6, Y6h6x6, F7h6x6, M7h6x6, T7h6x6, A8h6x6;
wire H8h6x6, O8h6x6, V8h6x6, C9h6x6, J9h6x6, Q9h6x6, X9h6x6, Eah6x6, Lah6x6, Sah6x6;
wire Zah6x6, Gbh6x6, Nbh6x6, Ubh6x6, Bch6x6, Ich6x6, Pch6x6, Wch6x6, Ddh6x6, Kdh6x6;
wire Rdh6x6, Ydh6x6, Feh6x6, Meh6x6, Teh6x6, Afh6x6, Hfh6x6, Ofh6x6, Vfh6x6, Cgh6x6;
wire Jgh6x6, Qgh6x6, Xgh6x6, Ehh6x6, Lhh6x6, Shh6x6, Zhh6x6, Gih6x6, Nih6x6, Uih6x6;
wire Bjh6x6, Ijh6x6, Pjh6x6, Wjh6x6, Dkh6x6, Kkh6x6, Rkh6x6, Ykh6x6, Flh6x6, Mlh6x6;
wire Tlh6x6, Amh6x6, Hmh6x6, Omh6x6, Vmh6x6, Cnh6x6, Jnh6x6, Qnh6x6, Xnh6x6, Eoh6x6;
wire Loh6x6, Soh6x6, Zoh6x6, Gph6x6, Nph6x6, Uph6x6, Bqh6x6, Iqh6x6, Pqh6x6, Wqh6x6;
wire Drh6x6, Krh6x6, Rrh6x6, Yrh6x6, Fsh6x6, Msh6x6, Tsh6x6, Ath6x6, Hth6x6, Oth6x6;
wire Vth6x6, Cuh6x6, Juh6x6, Quh6x6, Xuh6x6, Evh6x6, Lvh6x6, Svh6x6, Zvh6x6, Gwh6x6;
wire Nwh6x6, Uwh6x6, Bxh6x6, Ixh6x6, Pxh6x6, Wxh6x6, Dyh6x6, Kyh6x6, Ryh6x6, Yyh6x6;
wire Fzh6x6, Mzh6x6, Tzh6x6, A0i6x6, H0i6x6, O0i6x6, V0i6x6, C1i6x6, J1i6x6, Q1i6x6;
wire X1i6x6, E2i6x6, L2i6x6, S2i6x6, Z2i6x6, G3i6x6, N3i6x6, U3i6x6, B4i6x6, I4i6x6;
wire P4i6x6, W4i6x6, D5i6x6, K5i6x6, R5i6x6, Y5i6x6, F6i6x6, M6i6x6, T6i6x6, A7i6x6;
wire H7i6x6, O7i6x6, V7i6x6, C8i6x6, J8i6x6, Q8i6x6, X8i6x6, E9i6x6, L9i6x6, S9i6x6;
wire Z9i6x6, Gai6x6, Nai6x6, Uai6x6, Bbi6x6, Ibi6x6, Pbi6x6, Wbi6x6, Dci6x6, Kci6x6;
wire Rci6x6, Yci6x6, Fdi6x6, Mdi6x6, Tdi6x6, Aei6x6, Hei6x6, Oei6x6, Vei6x6, Cfi6x6;
wire Jfi6x6, Qfi6x6, Xfi6x6, Egi6x6, Lgi6x6, Sgi6x6, Zgi6x6, Ghi6x6, Nhi6x6, Uhi6x6;
wire Bii6x6, Iii6x6, Pii6x6, Wii6x6, Dji6x6, Kji6x6, Rji6x6, Yji6x6, Fki6x6, Mki6x6;
wire Tki6x6, Ali6x6, Hli6x6, Oli6x6, Vli6x6, Cmi6x6, Jmi6x6, Qmi6x6, Xmi6x6, Eni6x6;
wire Lni6x6, Sni6x6, Zni6x6, Goi6x6, Noi6x6, Uoi6x6, Bpi6x6, Ipi6x6, Ppi6x6, Wpi6x6;
wire Dqi6x6, Kqi6x6, Rqi6x6, Yqi6x6, Fri6x6, Mri6x6, Tri6x6, Asi6x6, Hsi6x6, Osi6x6;
wire Vsi6x6, Cti6x6, Jti6x6, Qti6x6, Xti6x6, Eui6x6, Lui6x6, Sui6x6, Zui6x6, Gvi6x6;
wire Nvi6x6, Uvi6x6, Bwi6x6, Iwi6x6, Pwi6x6, Wwi6x6, Dxi6x6, Kxi6x6, Rxi6x6, Yxi6x6;
wire Fyi6x6, Myi6x6, Tyi6x6, Azi6x6, Hzi6x6, Ozi6x6, Vzi6x6, C0j6x6, J0j6x6, Q0j6x6;
wire X0j6x6, E1j6x6, L1j6x6, S1j6x6, Z1j6x6, G2j6x6, N2j6x6, U2j6x6, B3j6x6, I3j6x6;
wire P3j6x6, W3j6x6, D4j6x6, K4j6x6, R4j6x6, Y4j6x6, F5j6x6, M5j6x6, T5j6x6, A6j6x6;
wire H6j6x6, O6j6x6, V6j6x6, C7j6x6, J7j6x6, Q7j6x6, X7j6x6, E8j6x6, L8j6x6, S8j6x6;
wire Z8j6x6, G9j6x6, N9j6x6, U9j6x6, Baj6x6, Iaj6x6, Paj6x6, Waj6x6, Dbj6x6, Kbj6x6;
wire Rbj6x6, Ybj6x6, Fcj6x6, Mcj6x6, Tcj6x6, Adj6x6, Hdj6x6, Odj6x6, Vdj6x6, Cej6x6;
wire Jej6x6, Qej6x6, Xej6x6, Efj6x6, Lfj6x6, Sfj6x6, Zfj6x6, Ggj6x6, Ngj6x6, Ugj6x6;
wire Bhj6x6, Ihj6x6, Phj6x6, Whj6x6, Dij6x6, Kij6x6, Rij6x6, Yij6x6, Fjj6x6, Mjj6x6;
wire Tjj6x6, Akj6x6, Hkj6x6, Okj6x6, Vkj6x6, Clj6x6, Jlj6x6, Qlj6x6, Xlj6x6, Emj6x6;
wire Lmj6x6, Smj6x6, Zmj6x6, Gnj6x6, Nnj6x6, Unj6x6, Boj6x6, Ioj6x6, Poj6x6, Woj6x6;
wire Dpj6x6, Kpj6x6, Rpj6x6, Ypj6x6, Fqj6x6, Mqj6x6, Tqj6x6, Arj6x6, Hrj6x6, Orj6x6;
wire Vrj6x6, Csj6x6, Jsj6x6, Qsj6x6, Xsj6x6, Etj6x6, Ltj6x6, Stj6x6, Ztj6x6, Guj6x6;
wire Nuj6x6, Uuj6x6, Bvj6x6, Ivj6x6, Pvj6x6, Wvj6x6, Dwj6x6, Kwj6x6, Rwj6x6, Ywj6x6;
wire Fxj6x6, Mxj6x6, Txj6x6, Ayj6x6, Hyj6x6, Oyj6x6, Vyj6x6, Czj6x6, Jzj6x6, Qzj6x6;
wire Xzj6x6, E0k6x6, L0k6x6, S0k6x6, Z0k6x6, G1k6x6, N1k6x6, U1k6x6, B2k6x6, I2k6x6;
wire P2k6x6, W2k6x6, D3k6x6, K3k6x6, R3k6x6, Y3k6x6, F4k6x6, M4k6x6, T4k6x6, A5k6x6;
wire H5k6x6, O5k6x6, V5k6x6, C6k6x6, J6k6x6, Q6k6x6, X6k6x6, E7k6x6, L7k6x6, S7k6x6;
wire Z7k6x6, G8k6x6, N8k6x6, U8k6x6, B9k6x6, I9k6x6, P9k6x6, W9k6x6, Dak6x6, Kak6x6;
wire Rak6x6, Yak6x6, Fbk6x6, Mbk6x6, Tbk6x6, Ack6x6, Hck6x6, Ock6x6, Vck6x6, Cdk6x6;
wire Jdk6x6, Qdk6x6, Xdk6x6, Eek6x6, Lek6x6, Sek6x6, Zek6x6, Gfk6x6, Nfk6x6, Ufk6x6;
wire Bgk6x6, Igk6x6, Pgk6x6, Wgk6x6, Dhk6x6, Khk6x6, Rhk6x6, Yhk6x6, Fik6x6, Mik6x6;
wire Tik6x6, Ajk6x6, Hjk6x6, Ojk6x6, Vjk6x6, Ckk6x6, Jkk6x6, Qkk6x6, Xkk6x6, Elk6x6;
wire Llk6x6, Slk6x6, Zlk6x6, Gmk6x6, Nmk6x6, Umk6x6, Bnk6x6, Ink6x6, Pnk6x6, Wnk6x6;
wire Dok6x6, Kok6x6, Rok6x6, Yok6x6, Fpk6x6, Mpk6x6, Tpk6x6, Aqk6x6, Hqk6x6, Oqk6x6;
wire Vqk6x6, Crk6x6, Jrk6x6, Qrk6x6, Xrk6x6, Esk6x6, Lsk6x6, Ssk6x6, Zsk6x6, Gtk6x6;
wire Ntk6x6, Utk6x6, Buk6x6, Iuk6x6, Puk6x6, Wuk6x6, Dvk6x6, Kvk6x6, Rvk6x6, Yvk6x6;
wire Fwk6x6, Mwk6x6, Twk6x6, Axk6x6, Hxk6x6, Oxk6x6, Vxk6x6, Cyk6x6, Jyk6x6, Qyk6x6;
wire Xyk6x6, Ezk6x6, Lzk6x6, Szk6x6, Zzk6x6, G0l6x6, N0l6x6, U0l6x6, B1l6x6, I1l6x6;
wire P1l6x6, W1l6x6, D2l6x6, K2l6x6, R2l6x6, Y2l6x6, F3l6x6, M3l6x6, T3l6x6, A4l6x6;
wire H4l6x6, O4l6x6, V4l6x6, C5l6x6, J5l6x6, Q5l6x6, X5l6x6, E6l6x6, L6l6x6, S6l6x6;
wire Z6l6x6, G7l6x6, N7l6x6, U7l6x6, B8l6x6, I8l6x6, P8l6x6, W8l6x6, D9l6x6, K9l6x6;
wire R9l6x6, Y9l6x6, Fal6x6, Mal6x6, Tal6x6, Abl6x6, Hbl6x6, Obl6x6, Vbl6x6, Ccl6x6;
wire Jcl6x6, Qcl6x6, Xcl6x6, Edl6x6, Ldl6x6, Sdl6x6, Zdl6x6, Gel6x6, Nel6x6, Uel6x6;
wire Bfl6x6, Ifl6x6, Pfl6x6, Wfl6x6, Dgl6x6, Kgl6x6, Rgl6x6, Ygl6x6, Fhl6x6, Mhl6x6;
wire Thl6x6, Ail6x6, Hil6x6, Oil6x6, Vil6x6, Cjl6x6, Jjl6x6, Qjl6x6, Xjl6x6, Ekl6x6;
wire Lkl6x6, Skl6x6, Zkl6x6, Gll6x6, Nll6x6, Ull6x6, Bml6x6, Iml6x6, Pml6x6, Wml6x6;
wire Dnl6x6, Knl6x6, Rnl6x6, Ynl6x6, Fol6x6, Mol6x6, Tol6x6, Apl6x6, Hpl6x6, Opl6x6;
wire Vpl6x6, Cql6x6, Jql6x6, Qql6x6, Xql6x6, Erl6x6, Lrl6x6, Srl6x6, Zrl6x6, Gsl6x6;
wire Nsl6x6, Usl6x6, Btl6x6, Itl6x6, Ptl6x6, Wtl6x6, Dul6x6, Kul6x6, Rul6x6, Yul6x6;
wire Fvl6x6, Mvl6x6, Tvl6x6, Awl6x6, Hwl6x6, Owl6x6, Vwl6x6, Cxl6x6, Jxl6x6, Qxl6x6;
wire Xxl6x6, Eyl6x6, Lyl6x6, Syl6x6, Zyl6x6, Gzl6x6, Nzl6x6, Uzl6x6, B0m6x6, I0m6x6;
wire P0m6x6, W0m6x6, D1m6x6, K1m6x6, R1m6x6, Y1m6x6, F2m6x6, M2m6x6, T2m6x6, A3m6x6;
wire H3m6x6, O3m6x6, V3m6x6, C4m6x6, J4m6x6, Q4m6x6, X4m6x6, E5m6x6, L5m6x6, S5m6x6;
wire Z5m6x6, G6m6x6, N6m6x6, U6m6x6, B7m6x6, I7m6x6, P7m6x6, W7m6x6, D8m6x6, K8m6x6;
wire R8m6x6, Y8m6x6, F9m6x6, M9m6x6, T9m6x6, Aam6x6, Ham6x6, Oam6x6, Vam6x6, Cbm6x6;
wire Jbm6x6, Qbm6x6, Xbm6x6, Ecm6x6, Lcm6x6, Scm6x6, Zcm6x6, Gdm6x6, Ndm6x6, Udm6x6;
wire Bem6x6, Iem6x6, Pem6x6, Wem6x6, Dfm6x6, Kfm6x6, Rfm6x6, Yfm6x6, Fgm6x6, Mgm6x6;
wire Tgm6x6, Ahm6x6, Hhm6x6, Ohm6x6, Vhm6x6, Cim6x6, Jim6x6, Qim6x6, Xim6x6, Ejm6x6;
wire Ljm6x6, Sjm6x6, Zjm6x6, Gkm6x6, Nkm6x6, Ukm6x6, Blm6x6, Ilm6x6, Plm6x6, Wlm6x6;
wire Dmm6x6, Kmm6x6, Rmm6x6, Ymm6x6, Fnm6x6, Mnm6x6, Tnm6x6, Aom6x6, Hom6x6, Oom6x6;
wire Vom6x6, Cpm6x6, Jpm6x6, Qpm6x6, Xpm6x6, Eqm6x6, Lqm6x6, Sqm6x6, Zqm6x6, Grm6x6;
wire Nrm6x6, Urm6x6, Bsm6x6, Ism6x6, Psm6x6, Wsm6x6, Dtm6x6, Ktm6x6, Rtm6x6, Ytm6x6;
wire Fum6x6, Mum6x6, Tum6x6, Avm6x6, Hvm6x6, Ovm6x6, Vvm6x6, Cwm6x6, Jwm6x6, Qwm6x6;
wire Xwm6x6, Exm6x6, Lxm6x6, Sxm6x6, Zxm6x6, Gym6x6, Nym6x6, Uym6x6, Bzm6x6, Izm6x6;
wire Pzm6x6, Wzm6x6, D0n6x6, K0n6x6, R0n6x6, Y0n6x6, F1n6x6, M1n6x6, T1n6x6, A2n6x6;
wire H2n6x6, O2n6x6, V2n6x6, C3n6x6, J3n6x6, Q3n6x6, X3n6x6, E4n6x6, L4n6x6, S4n6x6;
wire Z4n6x6, G5n6x6, N5n6x6, U5n6x6, B6n6x6, I6n6x6, P6n6x6, W6n6x6, D7n6x6, K7n6x6;
wire R7n6x6, Y7n6x6, F8n6x6, M8n6x6, T8n6x6, A9n6x6, H9n6x6, O9n6x6, V9n6x6, Can6x6;
wire Jan6x6, Qan6x6, Xan6x6, Ebn6x6, Lbn6x6, Sbn6x6, Zbn6x6, Gcn6x6, Ncn6x6, Ucn6x6;
wire Bdn6x6, Idn6x6, Pdn6x6, Wdn6x6, Den6x6, Ken6x6, Ren6x6, Yen6x6, Ffn6x6, Mfn6x6;
wire Tfn6x6, Agn6x6, Hgn6x6, Ogn6x6, Vgn6x6, Chn6x6, Jhn6x6, Qhn6x6, Xhn6x6, Ein6x6;
wire Lin6x6, Sin6x6, Zin6x6, Gjn6x6, Njn6x6, Ujn6x6, Bkn6x6, Ikn6x6, Pkn6x6, Wkn6x6;
wire Dln6x6, Kln6x6, Rln6x6, Yln6x6, Fmn6x6, Mmn6x6, Tmn6x6, Ann6x6, Hnn6x6, Onn6x6;
wire Vnn6x6, Con6x6, Jon6x6, Qon6x6, Xon6x6, Epn6x6, Lpn6x6, Spn6x6, Zpn6x6, Gqn6x6;
wire Nqn6x6, Uqn6x6, Brn6x6, Irn6x6, Prn6x6, Wrn6x6, Dsn6x6, Ksn6x6, Rsn6x6, Ysn6x6;
wire Ftn6x6, Mtn6x6, Ttn6x6, Aun6x6, Hun6x6, Oun6x6, Vun6x6, Cvn6x6, Jvn6x6, Qvn6x6;
wire Xvn6x6, Ewn6x6, Lwn6x6, Swn6x6, Zwn6x6, Gxn6x6, Nxn6x6, Uxn6x6, Byn6x6, Iyn6x6;
wire Pyn6x6, Wyn6x6, Dzn6x6, Kzn6x6, Rzn6x6, Yzn6x6, F0o6x6, M0o6x6, T0o6x6, A1o6x6;
wire H1o6x6, O1o6x6, V1o6x6, C2o6x6, J2o6x6, Q2o6x6, X2o6x6, E3o6x6, L3o6x6, S3o6x6;
wire Z3o6x6, G4o6x6, N4o6x6, U4o6x6, B5o6x6, I5o6x6, P5o6x6, W5o6x6, D6o6x6, K6o6x6;
wire R6o6x6, Y6o6x6, F7o6x6, M7o6x6, T7o6x6, A8o6x6, H8o6x6, O8o6x6, V8o6x6, C9o6x6;
wire J9o6x6, Q9o6x6, X9o6x6, Eao6x6, Lao6x6, Sao6x6, Zao6x6, Gbo6x6, Nbo6x6, Ubo6x6;
wire Bco6x6, Ico6x6, Pco6x6, Wco6x6, Ddo6x6, Kdo6x6, Rdo6x6, Ydo6x6, Feo6x6, Meo6x6;
wire Teo6x6, Afo6x6, Hfo6x6, Ofo6x6, Vfo6x6, Cgo6x6, Jgo6x6, Qgo6x6, Xgo6x6, Eho6x6;
wire Lho6x6, Sho6x6, Zho6x6, Gio6x6, Nio6x6, Uio6x6, Bjo6x6, Ijo6x6, Pjo6x6, Wjo6x6;
wire Dko6x6, Kko6x6, Rko6x6, Yko6x6, Flo6x6, Mlo6x6, Tlo6x6, Amo6x6, Hmo6x6, Omo6x6;
wire Vmo6x6, Cno6x6, Jno6x6, Qno6x6, Xno6x6, Eoo6x6, Loo6x6, Soo6x6, Zoo6x6, Gpo6x6;
wire Npo6x6, Upo6x6, Bqo6x6, Iqo6x6, Pqo6x6, Wqo6x6, Dro6x6, Kro6x6, Rro6x6, Yro6x6;
wire Fso6x6, Mso6x6, Tso6x6, Ato6x6, Hto6x6, Oto6x6, Vto6x6, Cuo6x6, Juo6x6, Quo6x6;
wire Xuo6x6, Evo6x6, Lvo6x6, Svo6x6, Zvo6x6, Gwo6x6, Nwo6x6, Uwo6x6, Bxo6x6, Ixo6x6;
wire Pxo6x6, Wxo6x6, Dyo6x6, Kyo6x6, Ryo6x6, Yyo6x6, Fzo6x6, Mzo6x6, Tzo6x6, A0p6x6;
wire H0p6x6, O0p6x6, V0p6x6, C1p6x6, J1p6x6, Q1p6x6, X1p6x6, E2p6x6, L2p6x6, S2p6x6;
wire Z2p6x6, G3p6x6, N3p6x6, U3p6x6, B4p6x6, I4p6x6, P4p6x6, W4p6x6, D5p6x6, K5p6x6;
wire R5p6x6, Y5p6x6, F6p6x6, M6p6x6, T6p6x6, A7p6x6, H7p6x6, O7p6x6, V7p6x6, C8p6x6;
wire J8p6x6, Q8p6x6, X8p6x6, E9p6x6, L9p6x6, S9p6x6, Z9p6x6, Gap6x6, Nap6x6, Uap6x6;
wire Bbp6x6, Ibp6x6, Pbp6x6, Wbp6x6, Dcp6x6, Kcp6x6, Rcp6x6, Ycp6x6, Fdp6x6, Mdp6x6;
wire Tdp6x6, Aep6x6, Hep6x6, Oep6x6, Vep6x6, Cfp6x6, Jfp6x6, Qfp6x6, Xfp6x6, Egp6x6;
wire Lgp6x6, Sgp6x6, Zgp6x6, Ghp6x6, Nhp6x6, Uhp6x6, Bip6x6, Iip6x6, Pip6x6, Wip6x6;
wire Djp6x6, Kjp6x6, Rjp6x6, Yjp6x6, Fkp6x6, Mkp6x6, Tkp6x6, Alp6x6, Hlp6x6, Olp6x6;
wire Vlp6x6, Cmp6x6, Jmp6x6, Qmp6x6, Xmp6x6, Enp6x6, Lnp6x6, Snp6x6, Znp6x6, Gop6x6;
wire Nop6x6, Uop6x6, Bpp6x6, Ipp6x6, Ppp6x6, Wpp6x6, Dqp6x6, Kqp6x6, Rqp6x6, Yqp6x6;
wire Frp6x6, Mrp6x6, Trp6x6, Asp6x6, Hsp6x6, Osp6x6, Vsp6x6, Ctp6x6, Jtp6x6, Qtp6x6;
wire Xtp6x6, Eup6x6, Lup6x6, Sup6x6, Zup6x6, Gvp6x6, Nvp6x6, Uvp6x6, Bwp6x6, Iwp6x6;
wire Pwp6x6, Wwp6x6, Dxp6x6, Kxp6x6, Rxp6x6, Yxp6x6, Fyp6x6, Myp6x6, Typ6x6, Azp6x6;
wire Hzp6x6, Ozp6x6, Vzp6x6, C0q6x6, J0q6x6, Q0q6x6, X0q6x6, E1q6x6, L1q6x6, S1q6x6;
wire Z1q6x6, G2q6x6, N2q6x6, U2q6x6, B3q6x6, I3q6x6, P3q6x6, W3q6x6, D4q6x6, K4q6x6;
wire R4q6x6, Y4q6x6, F5q6x6, M5q6x6, T5q6x6, A6q6x6, H6q6x6, O6q6x6, V6q6x6, C7q6x6;
wire J7q6x6, Q7q6x6, X7q6x6, E8q6x6, L8q6x6, S8q6x6, Z8q6x6, G9q6x6, N9q6x6, U9q6x6;
wire Baq6x6, Iaq6x6, Paq6x6, Waq6x6, Dbq6x6, Kbq6x6, Rbq6x6, Ybq6x6, Fcq6x6, Mcq6x6;
wire Tcq6x6, Adq6x6, Hdq6x6, Odq6x6, Vdq6x6, Ceq6x6, Jeq6x6, Qeq6x6, Xeq6x6, Efq6x6;
wire Lfq6x6, Sfq6x6, Zfq6x6, Ggq6x6, Ngq6x6, Ugq6x6, Bhq6x6, Ihq6x6, Phq6x6, Whq6x6;
wire Diq6x6, Kiq6x6, Riq6x6, Yiq6x6, Fjq6x6, Mjq6x6, Tjq6x6, Akq6x6, Hkq6x6, Okq6x6;
wire Vkq6x6, Clq6x6, Jlq6x6, Qlq6x6, Xlq6x6, Emq6x6, Lmq6x6, Smq6x6, Zmq6x6, Gnq6x6;
wire Nnq6x6, Unq6x6, Boq6x6, Ioq6x6, Poq6x6, Woq6x6, Dpq6x6, Kpq6x6, Rpq6x6, Ypq6x6;
wire Fqq6x6, Mqq6x6, Tqq6x6, Arq6x6, Hrq6x6, Orq6x6, Vrq6x6, Csq6x6, Jsq6x6, Qsq6x6;
wire Xsq6x6, Etq6x6, Ltq6x6, Stq6x6, Ztq6x6, Guq6x6, Nuq6x6, Uuq6x6, Bvq6x6, Ivq6x6;
wire Pvq6x6, Wvq6x6, Dwq6x6, Kwq6x6, Rwq6x6, Ywq6x6, Fxq6x6, Mxq6x6, Txq6x6, Ayq6x6;
wire Hyq6x6, Oyq6x6, Vyq6x6, Czq6x6, Jzq6x6, Qzq6x6, Xzq6x6, E0r6x6, L0r6x6, S0r6x6;
wire Z0r6x6, G1r6x6, N1r6x6, U1r6x6, B2r6x6, I2r6x6, P2r6x6, W2r6x6, D3r6x6, K3r6x6;
wire R3r6x6, Y3r6x6, F4r6x6, M4r6x6, T4r6x6, A5r6x6, H5r6x6, O5r6x6, V5r6x6, C6r6x6;
wire J6r6x6, Q6r6x6, X6r6x6, E7r6x6, L7r6x6, S7r6x6, Z7r6x6, G8r6x6, N8r6x6, U8r6x6;
wire B9r6x6, I9r6x6, P9r6x6, W9r6x6, Dar6x6, Kar6x6, Rar6x6, Yar6x6, Fbr6x6, Mbr6x6;
wire Tbr6x6, Acr6x6, Hcr6x6, Ocr6x6, Vcr6x6, Cdr6x6, Jdr6x6, Qdr6x6, Xdr6x6, Eer6x6;
wire Ler6x6, Ser6x6, Zer6x6, Gfr6x6, Nfr6x6, Ufr6x6, Bgr6x6, Igr6x6, Pgr6x6, Wgr6x6;
wire Dhr6x6, Khr6x6, Rhr6x6, Yhr6x6, Fir6x6, Mir6x6, Tir6x6, Ajr6x6, Hjr6x6, Ojr6x6;
wire Vjr6x6, Ckr6x6, Jkr6x6, Qkr6x6, Xkr6x6, Elr6x6, Llr6x6, Slr6x6, Zlr6x6, Gmr6x6;
wire Nmr6x6, Umr6x6, Bnr6x6, Inr6x6, Pnr6x6, Wnr6x6, Dor6x6, Kor6x6, Ror6x6, Yor6x6;
wire Fpr6x6, Mpr6x6, Tpr6x6, Aqr6x6, Hqr6x6, Oqr6x6, Vqr6x6, Crr6x6, Jrr6x6, Qrr6x6;
wire Xrr6x6, Esr6x6, Lsr6x6, Ssr6x6, Zsr6x6, Gtr6x6, Ntr6x6, Utr6x6, Bur6x6, Iur6x6;
wire Pur6x6, Wur6x6, Dvr6x6, Kvr6x6, Rvr6x6, Yvr6x6, Fwr6x6, Mwr6x6, Twr6x6, Axr6x6;
wire Hxr6x6, Oxr6x6, Vxr6x6, Cyr6x6, Jyr6x6, Qyr6x6, Xyr6x6, Ezr6x6, Lzr6x6, Szr6x6;
wire Zzr6x6, G0s6x6, N0s6x6, U0s6x6, B1s6x6, I1s6x6, P1s6x6, W1s6x6, D2s6x6, K2s6x6;
wire R2s6x6, Y2s6x6, F3s6x6, M3s6x6, T3s6x6, A4s6x6, H4s6x6, O4s6x6, V4s6x6, C5s6x6;
wire J5s6x6, Q5s6x6, X5s6x6, E6s6x6, L6s6x6, S6s6x6, Z6s6x6, G7s6x6, N7s6x6, U7s6x6;
wire B8s6x6, I8s6x6, P8s6x6, W8s6x6, D9s6x6, K9s6x6, R9s6x6, Y9s6x6, Fas6x6, Mas6x6;
wire Tas6x6, Abs6x6, Hbs6x6, Obs6x6, Vbs6x6, Ccs6x6, Jcs6x6, Qcs6x6, Xcs6x6, Eds6x6;
wire Lds6x6, Sds6x6, Zds6x6, Ges6x6, Nes6x6, Ues6x6, Bfs6x6, Ifs6x6, Pfs6x6, Wfs6x6;
wire Dgs6x6, Kgs6x6, Rgs6x6, Ygs6x6, Fhs6x6, Mhs6x6, Ths6x6, Ais6x6, His6x6, Ois6x6;
wire Vis6x6, Cjs6x6, Jjs6x6, Qjs6x6, Xjs6x6, Eks6x6, Lks6x6, Sks6x6, Zks6x6, Gls6x6;
wire Nls6x6, Uls6x6, Bms6x6, Ims6x6, Pms6x6, Wms6x6, Dns6x6, Kns6x6, Rns6x6, Yns6x6;
wire Fos6x6, Mos6x6, Tos6x6, Aps6x6, Hps6x6, Ops6x6, Vps6x6, Cqs6x6, Jqs6x6, Qqs6x6;
wire Xqs6x6, Ers6x6, Lrs6x6, Srs6x6, Zrs6x6, Gss6x6, Nss6x6, Uss6x6, Bts6x6, Its6x6;
wire Pts6x6, Wts6x6, Dus6x6, Kus6x6, Rus6x6, Yus6x6, Fvs6x6, Mvs6x6, Tvs6x6, Aws6x6;
wire Hws6x6, Ows6x6, Vws6x6, Cxs6x6, Jxs6x6, Qxs6x6, Xxs6x6, Eys6x6, Lys6x6, Sys6x6;
wire Zys6x6, Gzs6x6, Nzs6x6, Uzs6x6, B0t6x6, I0t6x6, P0t6x6, W0t6x6, D1t6x6, K1t6x6;
wire R1t6x6, Y1t6x6, F2t6x6, M2t6x6, T2t6x6, A3t6x6, H3t6x6, O3t6x6, V3t6x6, C4t6x6;
wire J4t6x6, Q4t6x6, X4t6x6, E5t6x6, L5t6x6, S5t6x6, Z5t6x6, G6t6x6, N6t6x6, U6t6x6;
wire B7t6x6, I7t6x6, P7t6x6, W7t6x6, D8t6x6, K8t6x6, R8t6x6, Y8t6x6, F9t6x6, M9t6x6;
wire T9t6x6, Aat6x6, Hat6x6, Oat6x6, Vat6x6, Cbt6x6, Jbt6x6, Qbt6x6, Xbt6x6, Ect6x6;
wire Lct6x6, Sct6x6, Zct6x6, Gdt6x6, Ndt6x6, Udt6x6, Bet6x6, Iet6x6, Pet6x6, Wet6x6;
wire Dft6x6, Kft6x6, Rft6x6, Yft6x6, Fgt6x6, Mgt6x6, Tgt6x6, Aht6x6, Hht6x6, Oht6x6;
wire Vht6x6, Cit6x6, Jit6x6, Qit6x6, Xit6x6, Ejt6x6, Ljt6x6, Sjt6x6, Zjt6x6, Gkt6x6;
wire Nkt6x6, Ukt6x6, Blt6x6, Ilt6x6, Plt6x6, Wlt6x6, Dmt6x6, Kmt6x6, Rmt6x6, Ymt6x6;
wire Fnt6x6, Mnt6x6, Tnt6x6, Aot6x6, Hot6x6, Oot6x6, Vot6x6, Cpt6x6, Jpt6x6, Qpt6x6;
wire Xpt6x6, Eqt6x6, Lqt6x6, Sqt6x6, Zqt6x6, Grt6x6, Nrt6x6, Urt6x6, Bst6x6, Ist6x6;
wire Pst6x6, Wst6x6, Dtt6x6, Ktt6x6, Rtt6x6, Ytt6x6, Fut6x6, Mut6x6, Tut6x6, Avt6x6;
wire Hvt6x6, Ovt6x6, Vvt6x6, Cwt6x6, Jwt6x6, Qwt6x6, Xwt6x6, Ext6x6, Lxt6x6, Sxt6x6;
wire Zxt6x6, Gyt6x6, Nyt6x6, Uyt6x6, Bzt6x6, Izt6x6, Pzt6x6, Wzt6x6, D0u6x6, K0u6x6;
wire R0u6x6, Y0u6x6, F1u6x6, M1u6x6, T1u6x6, A2u6x6, H2u6x6, O2u6x6, V2u6x6, C3u6x6;
wire J3u6x6, Q3u6x6, X3u6x6, E4u6x6, L4u6x6, S4u6x6, Z4u6x6, G5u6x6, N5u6x6, U5u6x6;
wire B6u6x6, I6u6x6, P6u6x6, W6u6x6, D7u6x6, K7u6x6, R7u6x6, Y7u6x6, F8u6x6, M8u6x6;
wire T8u6x6, A9u6x6, H9u6x6, O9u6x6, V9u6x6, Cau6x6, Jau6x6, Qau6x6, Xau6x6, Ebu6x6;
wire Lbu6x6, Sbu6x6, Zbu6x6, Gcu6x6, Ncu6x6, Ucu6x6, Bdu6x6, Idu6x6, Pdu6x6, Wdu6x6;
wire Deu6x6, Keu6x6, Reu6x6, Yeu6x6, Ffu6x6, Mfu6x6, Tfu6x6, Agu6x6, Hgu6x6, Ogu6x6;
wire Vgu6x6, Chu6x6, Jhu6x6, Qhu6x6, Xhu6x6, Eiu6x6, Liu6x6, Siu6x6, Ziu6x6, Gju6x6;
wire Nju6x6, Uju6x6, Bku6x6, Iku6x6, Pku6x6, Wku6x6, Dlu6x6, Klu6x6, Rlu6x6, Ylu6x6;
wire Fmu6x6, Mmu6x6, Tmu6x6, Anu6x6, Hnu6x6, Onu6x6, Vnu6x6, Cou6x6, Jou6x6, Qou6x6;
wire Xou6x6, Epu6x6, Lpu6x6, Spu6x6, Zpu6x6, Gqu6x6, Nqu6x6, Uqu6x6, Bru6x6, Iru6x6;
wire Pru6x6, Wru6x6, Dsu6x6, Ksu6x6, Rsu6x6, Ysu6x6, Ftu6x6, Mtu6x6, Ttu6x6, Auu6x6;
wire Huu6x6, Ouu6x6, Vuu6x6, Cvu6x6, Jvu6x6, Qvu6x6, Xvu6x6, Ewu6x6, Lwu6x6, Swu6x6;
wire Zwu6x6, Gxu6x6, Nxu6x6, Uxu6x6, Byu6x6, Iyu6x6, Pyu6x6, Wyu6x6, Dzu6x6, Kzu6x6;
wire Rzu6x6, Yzu6x6, F0v6x6, M0v6x6, T0v6x6, A1v6x6, H1v6x6, O1v6x6, V1v6x6, C2v6x6;
wire J2v6x6, Q2v6x6, X2v6x6, E3v6x6, L3v6x6, S3v6x6, Z3v6x6, G4v6x6, N4v6x6, U4v6x6;
wire B5v6x6, I5v6x6, P5v6x6, W5v6x6, D6v6x6, K6v6x6, R6v6x6, Y6v6x6, F7v6x6, M7v6x6;
wire T7v6x6, A8v6x6, H8v6x6, O8v6x6, V8v6x6, C9v6x6, J9v6x6, Q9v6x6, X9v6x6, Eav6x6;
wire Lav6x6, Sav6x6, Zav6x6, Gbv6x6, Nbv6x6, Ubv6x6, Bcv6x6, Icv6x6, Pcv6x6, Wcv6x6;
wire Ddv6x6, Kdv6x6, Rdv6x6, Ydv6x6, Fev6x6, Mev6x6, Tev6x6, Afv6x6, Hfv6x6, Ofv6x6;
wire Vfv6x6, Cgv6x6, Jgv6x6, Qgv6x6, Xgv6x6, Ehv6x6, Lhv6x6, Shv6x6, Zhv6x6, Giv6x6;
wire Niv6x6, Uiv6x6, Bjv6x6, Ijv6x6, Pjv6x6, Wjv6x6, Dkv6x6, Kkv6x6, Rkv6x6, Ykv6x6;
wire Flv6x6, Mlv6x6, Tlv6x6, Amv6x6, Hmv6x6, Omv6x6, Vmv6x6, Cnv6x6, Jnv6x6, Qnv6x6;
wire Xnv6x6, Eov6x6, Lov6x6, Sov6x6, Zov6x6, Gpv6x6, Npv6x6, Upv6x6, Bqv6x6, Iqv6x6;
wire Pqv6x6, Wqv6x6, Drv6x6, Krv6x6, Rrv6x6, Yrv6x6, Fsv6x6, Msv6x6, Tsv6x6, Atv6x6;
wire Htv6x6, Otv6x6, Vtv6x6, Cuv6x6, Juv6x6, Quv6x6, Xuv6x6, Evv6x6, Lvv6x6, Svv6x6;
wire Zvv6x6, Gwv6x6, Nwv6x6, Uwv6x6, Bxv6x6, Ixv6x6, Pxv6x6, Wxv6x6, Dyv6x6, Kyv6x6;
wire Ryv6x6, Yyv6x6, Fzv6x6, Mzv6x6, Tzv6x6, A0w6x6, H0w6x6, O0w6x6, V0w6x6, C1w6x6;
wire J1w6x6, Q1w6x6, X1w6x6, E2w6x6, L2w6x6, S2w6x6, Z2w6x6, G3w6x6, N3w6x6, U3w6x6;
wire B4w6x6, I4w6x6, P4w6x6, W4w6x6, D5w6x6, K5w6x6, R5w6x6, Y5w6x6, F6w6x6, M6w6x6;
wire T6w6x6, A7w6x6, H7w6x6, O7w6x6, V7w6x6, C8w6x6, J8w6x6, Q8w6x6, X8w6x6, E9w6x6;
wire L9w6x6, S9w6x6, Z9w6x6, Gaw6x6, Naw6x6, Uaw6x6, Bbw6x6, Ibw6x6, Pbw6x6, Wbw6x6;
wire Dcw6x6, Kcw6x6, Rcw6x6, Ycw6x6, Fdw6x6, Mdw6x6, Tdw6x6, Aew6x6, Hew6x6, Oew6x6;
wire Vew6x6, Cfw6x6, Jfw6x6, Qfw6x6, Xfw6x6, Egw6x6, Lgw6x6, Sgw6x6, Zgw6x6, Ghw6x6;
wire Nhw6x6, Uhw6x6, Biw6x6, Iiw6x6, Piw6x6, Wiw6x6, Djw6x6, Kjw6x6, Rjw6x6, Yjw6x6;
wire Fkw6x6, Mkw6x6, Tkw6x6, Alw6x6, Hlw6x6, Olw6x6, Vlw6x6, Cmw6x6, Jmw6x6, Qmw6x6;
wire Xmw6x6, Enw6x6, Lnw6x6, Snw6x6, Znw6x6, Gow6x6, Now6x6, Uow6x6, Bpw6x6, Ipw6x6;
wire Ppw6x6, Wpw6x6, Dqw6x6, Kqw6x6, Rqw6x6, Yqw6x6, Frw6x6, Mrw6x6, Trw6x6, Asw6x6;
wire Hsw6x6, Osw6x6, Vsw6x6, Ctw6x6, Jtw6x6, Qtw6x6, Xtw6x6, Euw6x6, Luw6x6, Suw6x6;
wire Zuw6x6, Gvw6x6, Nvw6x6, Uvw6x6, Bww6x6, Iww6x6, Pww6x6, Www6x6, Dxw6x6, Kxw6x6;
wire Rxw6x6, Yxw6x6, Fyw6x6, Myw6x6, Tyw6x6, Azw6x6, Hzw6x6, Ozw6x6, Vzw6x6, C0x6x6;
wire J0x6x6, Q0x6x6, X0x6x6, E1x6x6, L1x6x6, S1x6x6, Z1x6x6, G2x6x6, N2x6x6, U2x6x6;
wire B3x6x6, I3x6x6, P3x6x6, W3x6x6, D4x6x6, K4x6x6, R4x6x6, Y4x6x6, F5x6x6, M5x6x6;
wire T5x6x6, A6x6x6, H6x6x6, O6x6x6, V6x6x6, C7x6x6, J7x6x6, Q7x6x6, X7x6x6, E8x6x6;
wire L8x6x6, S8x6x6, Z8x6x6, G9x6x6, N9x6x6, U9x6x6, Bax6x6, Iax6x6, Pax6x6, Wax6x6;
wire Dbx6x6, Kbx6x6, Rbx6x6, Ybx6x6, Fcx6x6, Mcx6x6, Tcx6x6, Adx6x6, Hdx6x6, Odx6x6;
wire Vdx6x6, Cex6x6, Jex6x6, Qex6x6, Xex6x6, Efx6x6, Lfx6x6, Sfx6x6, Zfx6x6, Ggx6x6;
wire Ngx6x6, Ugx6x6, Bhx6x6, Ihx6x6, Phx6x6, Whx6x6, Dix6x6, Kix6x6, Rix6x6, Yix6x6;
wire Fjx6x6, Mjx6x6, Tjx6x6, Akx6x6, Hkx6x6, Okx6x6, Vkx6x6, Clx6x6, Jlx6x6, Qlx6x6;
wire Xlx6x6, Emx6x6, Lmx6x6, Smx6x6, Zmx6x6, Gnx6x6, Nnx6x6, Unx6x6, Box6x6, Iox6x6;
wire Pox6x6, Wox6x6, Dpx6x6, Kpx6x6, Rpx6x6, Ypx6x6, Fqx6x6, Mqx6x6, Tqx6x6, Arx6x6;
wire Hrx6x6, Orx6x6, Vrx6x6, Csx6x6, Jsx6x6, Qsx6x6, Xsx6x6, Etx6x6, Ltx6x6, Stx6x6;
wire Ztx6x6, Gux6x6, Nux6x6, Uux6x6, Bvx6x6, Ivx6x6, Pvx6x6, Wvx6x6, Dwx6x6, Kwx6x6;
wire Rwx6x6, Ywx6x6, Fxx6x6, Mxx6x6, Txx6x6, Ayx6x6, Hyx6x6, Oyx6x6, Vyx6x6, Czx6x6;
wire Jzx6x6, Qzx6x6, Xzx6x6, E0y6x6, L0y6x6, S0y6x6, Z0y6x6, G1y6x6, N1y6x6, U1y6x6;
wire B2y6x6, I2y6x6, P2y6x6, W2y6x6, D3y6x6, K3y6x6, R3y6x6, Y3y6x6, F4y6x6, M4y6x6;
wire T4y6x6, A5y6x6, H5y6x6, O5y6x6, V5y6x6, C6y6x6, J6y6x6, Q6y6x6, X6y6x6, E7y6x6;
wire L7y6x6, S7y6x6, Z7y6x6, G8y6x6, N8y6x6, U8y6x6, B9y6x6, I9y6x6, P9y6x6, W9y6x6;
wire Day6x6, Kay6x6, Ray6x6, Yay6x6, Fby6x6, Mby6x6, Tby6x6, Acy6x6, Hcy6x6, Ocy6x6;
wire Vcy6x6, Cdy6x6, Jdy6x6, Qdy6x6, Xdy6x6, Eey6x6, Ley6x6, Sey6x6, Zey6x6, Gfy6x6;
wire Nfy6x6, Ufy6x6, Bgy6x6, Igy6x6, Pgy6x6, Wgy6x6, Dhy6x6, Khy6x6, Rhy6x6, Yhy6x6;
wire Fiy6x6, Miy6x6, Tiy6x6, Ajy6x6, Hjy6x6, Ojy6x6, Vjy6x6, Cky6x6, Jky6x6, Qky6x6;
wire Xky6x6, Ely6x6, Lly6x6, Sly6x6, Zly6x6, Gmy6x6, Nmy6x6, Umy6x6, Bny6x6, Iny6x6;
wire Pny6x6, Wny6x6, Doy6x6, Koy6x6, Roy6x6, Yoy6x6, Fpy6x6, Mpy6x6, Tpy6x6, Aqy6x6;
wire Hqy6x6, Oqy6x6, Vqy6x6, Cry6x6, Jry6x6, Qry6x6, Xry6x6, Esy6x6, Lsy6x6, Ssy6x6;
wire Zsy6x6, Gty6x6, Nty6x6, Uty6x6, Buy6x6, Iuy6x6, Puy6x6, Wuy6x6, Dvy6x6, Kvy6x6;
wire Rvy6x6, Yvy6x6, Fwy6x6, Mwy6x6, Twy6x6, Axy6x6, Hxy6x6, Oxy6x6, Vxy6x6, Cyy6x6;
wire Jyy6x6, Qyy6x6, Xyy6x6, Ezy6x6, Lzy6x6, Szy6x6, Zzy6x6, G0z6x6, N0z6x6, U0z6x6;
wire B1z6x6, I1z6x6, P1z6x6, W1z6x6, D2z6x6, K2z6x6, R2z6x6, Y2z6x6, F3z6x6, M3z6x6;
wire T3z6x6, A4z6x6, H4z6x6, O4z6x6, V4z6x6, C5z6x6, J5z6x6, Q5z6x6, X5z6x6, E6z6x6;
wire L6z6x6, S6z6x6, Z6z6x6, G7z6x6, N7z6x6, U7z6x6, B8z6x6, I8z6x6, P8z6x6, W8z6x6;
wire D9z6x6, K9z6x6, R9z6x6, Y9z6x6, Faz6x6, Maz6x6, Taz6x6, Abz6x6, Hbz6x6, Obz6x6;
wire Vbz6x6, Ccz6x6, Jcz6x6, Qcz6x6, Xcz6x6, Edz6x6, Ldz6x6, Sdz6x6, Zdz6x6, Gez6x6;
wire Nez6x6, Uez6x6, Bfz6x6, Ifz6x6, Pfz6x6, Wfz6x6, Dgz6x6, Kgz6x6, Rgz6x6, Ygz6x6;
wire Fhz6x6, Mhz6x6, Thz6x6, Aiz6x6, Hiz6x6, Oiz6x6, Viz6x6, Cjz6x6, Jjz6x6, Qjz6x6;
wire Xjz6x6, Ekz6x6, Lkz6x6, Skz6x6, Zkz6x6, Glz6x6, Nlz6x6, Ulz6x6, Bmz6x6, Imz6x6;
wire Pmz6x6, Wmz6x6, Dnz6x6, Knz6x6, Rnz6x6, Ynz6x6, Foz6x6, Moz6x6, Toz6x6, Apz6x6;
wire Hpz6x6, Opz6x6, Vpz6x6, Cqz6x6, Jqz6x6, Qqz6x6, Xqz6x6, Erz6x6, Lrz6x6, Srz6x6;
wire Zrz6x6, Gsz6x6, Nsz6x6, Usz6x6, Btz6x6, Itz6x6, Ptz6x6, Wtz6x6, Duz6x6, Kuz6x6;
wire Ruz6x6, Yuz6x6, Fvz6x6, Mvz6x6, Tvz6x6, Awz6x6, Hwz6x6, Owz6x6, Vwz6x6, Cxz6x6;
wire Jxz6x6, Qxz6x6, Xxz6x6, Eyz6x6, Lyz6x6, Syz6x6, Zyz6x6, Gzz6x6, Nzz6x6, Uzz6x6;
wire B007x6, I007x6, P007x6, W007x6, D107x6, K107x6, R107x6, Y107x6, F207x6, M207x6;
wire T207x6, A307x6, H307x6, O307x6, V307x6, C407x6, J407x6, Q407x6, X407x6, E507x6;
wire L507x6, S507x6, Z507x6, G607x6, N607x6, U607x6, B707x6, I707x6, P707x6, W707x6;
wire D807x6, K807x6, R807x6, Y807x6, F907x6, M907x6, T907x6, Aa07x6, Ha07x6, Oa07x6;
wire Va07x6, Cb07x6, Jb07x6, Qb07x6, Xb07x6, Ec07x6, Lc07x6, Sc07x6, Zc07x6, Gd07x6;
wire Nd07x6, Ud07x6, Be07x6, Ie07x6, Pe07x6, We07x6, Df07x6, Kf07x6, Rf07x6, Yf07x6;
wire Fg07x6, Mg07x6, Tg07x6, Ah07x6, Hh07x6, Oh07x6, Vh07x6, Ci07x6, Ji07x6, Qi07x6;
wire Xi07x6, Ej07x6, Lj07x6, Sj07x6, Zj07x6, Gk07x6, Nk07x6, Uk07x6, Bl07x6, Il07x6;
wire Pl07x6, Wl07x6, Dm07x6, Km07x6, Rm07x6, Ym07x6, Fn07x6, Mn07x6, Tn07x6, Ao07x6;
wire Ho07x6, Oo07x6, Vo07x6, Cp07x6, Jp07x6, Qp07x6, Xp07x6, Eq07x6, Lq07x6, Sq07x6;
wire Zq07x6, Gr07x6, Nr07x6, Ur07x6, Bs07x6, Is07x6, Ps07x6, Ws07x6, Dt07x6, Kt07x6;
wire Rt07x6, Yt07x6, Fu07x6, Mu07x6, Tu07x6, Av07x6, Hv07x6, Ov07x6, Vv07x6, Cw07x6;
wire Jw07x6, Qw07x6, Xw07x6, Ex07x6, Lx07x6, Sx07x6, Zx07x6, Gy07x6, Ny07x6, Uy07x6;
wire Bz07x6, Iz07x6, Pz07x6, Wz07x6, D017x6, K017x6, R017x6, Y017x6, F117x6, M117x6;
wire T117x6, A217x6, H217x6, O217x6, V217x6, C317x6, J317x6, Q317x6, X317x6, E417x6;
wire L417x6, S417x6, Z417x6, G517x6, N517x6, U517x6, B617x6, I617x6, P617x6, W617x6;
wire D717x6, K717x6, R717x6, Y717x6, F817x6, M817x6, T817x6, A917x6, H917x6, O917x6;
wire V917x6, Ca17x6, Ja17x6, Qa17x6, Xa17x6, Eb17x6, Lb17x6, Sb17x6, Zb17x6, Gc17x6;
wire Nc17x6, Uc17x6, Bd17x6, Id17x6, Pd17x6, Wd17x6, De17x6, Ke17x6, Re17x6, Ye17x6;
wire Ff17x6, Mf17x6, Tf17x6, Ag17x6, Hg17x6, Og17x6, Vg17x6, Ch17x6, Jh17x6, Qh17x6;
wire Xh17x6, Ei17x6, Li17x6, Si17x6, Zi17x6, Gj17x6, Nj17x6, Uj17x6, Bk17x6, Ik17x6;
wire Pk17x6, Wk17x6, Dl17x6, Kl17x6, Rl17x6, Yl17x6, Fm17x6, Mm17x6, Tm17x6, An17x6;
wire Hn17x6, On17x6, Vn17x6, Co17x6, Jo17x6, Qo17x6, Xo17x6, Ep17x6, Lp17x6, Sp17x6;
wire Zp17x6, Gq17x6, Nq17x6, Uq17x6, Br17x6, Ir17x6, Pr17x6, Wr17x6, Ds17x6, Ks17x6;
wire Rs17x6, Ys17x6, Ft17x6, Mt17x6, Tt17x6, Au17x6, Hu17x6, Ou17x6, Vu17x6, Cv17x6;
wire Jv17x6, Qv17x6, Xv17x6, Ew17x6, Lw17x6, Sw17x6, Zw17x6, Gx17x6, Nx17x6, Ux17x6;
wire By17x6, Iy17x6, Py17x6, Wy17x6, Dz17x6, Kz17x6, Rz17x6, Yz17x6, F027x6, M027x6;
wire T027x6, A127x6, H127x6, O127x6, V127x6, C227x6, J227x6, Q227x6, X227x6, E327x6;
wire L327x6, S327x6, Z327x6, G427x6, N427x6, U427x6, B527x6, I527x6, P527x6, W527x6;
wire D627x6, K627x6, R627x6, Y627x6, F727x6, M727x6, T727x6, A827x6, H827x6, O827x6;
wire V827x6, C927x6, J927x6, Q927x6, X927x6, Ea27x6, La27x6, Sa27x6, Za27x6, Gb27x6;
wire Nb27x6, Ub27x6, Bc27x6, Ic27x6, Pc27x6, Wc27x6, Dd27x6, Kd27x6, Rd27x6, Yd27x6;
wire Fe27x6, Me27x6, Te27x6, Af27x6, Hf27x6, Of27x6, Vf27x6, Cg27x6, Jg27x6, Qg27x6;
wire Xg27x6, Eh27x6, Lh27x6, Sh27x6, Zh27x6, Gi27x6, Ni27x6, Ui27x6, Bj27x6, Ij27x6;
wire Pj27x6, Wj27x6, Dk27x6, Kk27x6, Rk27x6, Yk27x6, Fl27x6, Ml27x6, Tl27x6, Am27x6;
wire Hm27x6, Om27x6, Vm27x6, Cn27x6, Jn27x6, Qn27x6, Xn27x6, Eo27x6, Lo27x6, So27x6;
wire Zo27x6, Gp27x6, Np27x6, Up27x6, Bq27x6, Iq27x6, Pq27x6, Wq27x6, Dr27x6, Kr27x6;
wire Rr27x6, Yr27x6, Fs27x6, Ms27x6, Ts27x6, At27x6, Ht27x6, Ot27x6, Vt27x6, Cu27x6;
wire Ju27x6, Qu27x6, Xu27x6, Ev27x6, Lv27x6, Sv27x6, Zv27x6, Gw27x6, Nw27x6, Uw27x6;
wire Bx27x6, Ix27x6, Px27x6, Wx27x6, Dy27x6, Ky27x6, Ry27x6, Yy27x6, Fz27x6, Mz27x6;
wire Tz27x6, A037x6, H037x6, O037x6, V037x6, C137x6, J137x6, Q137x6, X137x6, E237x6;
wire L237x6, S237x6, Z237x6, G337x6, N337x6, U337x6, B437x6, I437x6, P437x6, W437x6;
wire D537x6, K537x6, R537x6, Y537x6, F637x6, M637x6, T637x6, A737x6, H737x6, O737x6;
wire V737x6, C837x6, J837x6, Q837x6, X837x6, E937x6, L937x6, S937x6, Z937x6, Ga37x6;
wire Na37x6, Ua37x6, Bb37x6, Ib37x6, Pb37x6, Wb37x6, Dc37x6, Kc37x6, Rc37x6, Yc37x6;
wire Fd37x6, Md37x6, Td37x6, Ae37x6, He37x6, Oe37x6, Ve37x6, Cf37x6, Jf37x6, Qf37x6;
wire Xf37x6, Eg37x6, Lg37x6, Sg37x6, Zg37x6, Gh37x6, Nh37x6, Uh37x6, Bi37x6, Ii37x6;
wire Pi37x6, Wi37x6, Dj37x6, Kj37x6, Rj37x6, Yj37x6, Fk37x6, Mk37x6, Tk37x6, Al37x6;
wire Hl37x6, Ol37x6, Vl37x6, Cm37x6, Jm37x6, Qm37x6, Xm37x6, En37x6, Ln37x6, Sn37x6;
wire Zn37x6, Go37x6, No37x6, Uo37x6, Bp37x6, Ip37x6, Pp37x6, Wp37x6, Dq37x6, Kq37x6;
wire Rq37x6, Yq37x6, Fr37x6, Mr37x6, Tr37x6, As37x6, Hs37x6, Os37x6, Vs37x6, Ct37x6;
wire Jt37x6, Qt37x6, Xt37x6, Eu37x6, Lu37x6, Su37x6, Zu37x6, Gv37x6, Nv37x6, Uv37x6;
wire Bw37x6, Iw37x6, Pw37x6, Ww37x6, Dx37x6, Kx37x6, Rx37x6, Yx37x6, Fy37x6, My37x6;
wire Ty37x6, Az37x6, Hz37x6, Oz37x6, Vz37x6, C047x6, J047x6, Q047x6, X047x6, E147x6;
wire L147x6, S147x6, Z147x6, G247x6, N247x6, U247x6, B347x6, I347x6, P347x6, W347x6;
wire D447x6, K447x6, R447x6, Y447x6, F547x6, M547x6, T547x6, A647x6, H647x6, O647x6;
wire V647x6, C747x6, J747x6, Q747x6, X747x6, E847x6, L847x6, S847x6, Z847x6, G947x6;
wire N947x6, U947x6, Ba47x6, Ia47x6, Pa47x6, Wa47x6, Db47x6, Kb47x6, Rb47x6, Yb47x6;
wire Fc47x6, Mc47x6, Tc47x6, Ad47x6, Hd47x6, Od47x6, Vd47x6, Ce47x6, Je47x6, Qe47x6;
wire Xe47x6, Ef47x6, Lf47x6, Sf47x6, Zf47x6, Gg47x6, Ng47x6, Ug47x6, Bh47x6, Ih47x6;
wire Ph47x6, Wh47x6, Di47x6, Ki47x6, Ri47x6, Yi47x6, Fj47x6, Mj47x6, Tj47x6, Ak47x6;
wire Hk47x6, Ok47x6, Vk47x6, Cl47x6, Jl47x6, Ql47x6, Xl47x6, Em47x6, Lm47x6, Sm47x6;
wire Zm47x6, Gn47x6, Nn47x6, Un47x6, Bo47x6, Io47x6, Po47x6, Wo47x6, Dp47x6, Kp47x6;
wire Rp47x6, Yp47x6, Fq47x6, Mq47x6, Tq47x6, Ar47x6, Hr47x6, Or47x6, Vr47x6, Cs47x6;
wire Js47x6, Qs47x6, Xs47x6, Et47x6, Lt47x6, St47x6, Zt47x6, Gu47x6, Nu47x6, Uu47x6;
wire Bv47x6, Iv47x6, Pv47x6, Wv47x6, Dw47x6, Kw47x6, Rw47x6, Yw47x6, Fx47x6, Mx47x6;
wire Tx47x6, Ay47x6, Hy47x6, Oy47x6, Vy47x6, Cz47x6, Jz47x6, Qz47x6, Xz47x6, E057x6;
wire L057x6, S057x6, Z057x6, G157x6, N157x6, U157x6, B257x6, I257x6, P257x6, W257x6;
wire D357x6, K357x6, R357x6, Y357x6, F457x6, M457x6, T457x6, A557x6, H557x6, O557x6;
wire V557x6, C657x6, J657x6, Q657x6, X657x6, E757x6, L757x6, S757x6, Z757x6, G857x6;
wire N857x6, U857x6, B957x6, I957x6, P957x6, W957x6, Da57x6, Ka57x6, Ra57x6, Ya57x6;
wire Fb57x6, Mb57x6, Tb57x6, Ac57x6, Hc57x6, Oc57x6, Vc57x6, Cd57x6, Jd57x6, Qd57x6;
wire Xd57x6, Ee57x6, Le57x6, Se57x6, Ze57x6, Gf57x6, Nf57x6, Uf57x6, Bg57x6, Ig57x6;
wire Pg57x6, Wg57x6, Dh57x6, Kh57x6, Rh57x6, Yh57x6, Fi57x6, Mi57x6, Ti57x6, Aj57x6;
wire Hj57x6, Oj57x6, Vj57x6, Ck57x6, Jk57x6, Qk57x6, Xk57x6, El57x6, Ll57x6, Sl57x6;
wire Zl57x6, Gm57x6, Nm57x6, Um57x6, Bn57x6, In57x6, Pn57x6, Wn57x6, Do57x6, Ko57x6;
wire Ro57x6, Yo57x6, Fp57x6, Mp57x6, Tp57x6, Aq57x6, Hq57x6, Oq57x6, Vq57x6, Cr57x6;
wire Jr57x6, Qr57x6, Xr57x6, Es57x6, Ls57x6, Ss57x6, Zs57x6, Gt57x6, Nt57x6, Ut57x6;
wire Bu57x6, Iu57x6, Pu57x6, Wu57x6, Dv57x6, Kv57x6, Rv57x6, Yv57x6, Fw57x6, Mw57x6;
wire Tw57x6, Ax57x6, Hx57x6, Ox57x6, Vx57x6, Cy57x6, Jy57x6, Qy57x6, Xy57x6, Ez57x6;
wire Lz57x6, Sz57x6, Zz57x6, G067x6, N067x6, U067x6, B167x6, I167x6, P167x6, W167x6;
wire D267x6, K267x6, R267x6, Y267x6, F367x6, M367x6, T367x6, A467x6, H467x6, O467x6;
wire V467x6, C567x6, J567x6, Q567x6, X567x6, E667x6, L667x6, S667x6, Z667x6, G767x6;
wire N767x6, U767x6, B867x6, I867x6, P867x6, W867x6, D967x6, K967x6, R967x6, Y967x6;
wire Fa67x6, Ma67x6, Ta67x6, Ab67x6, Hb67x6, Ob67x6, Vb67x6, Cc67x6, Jc67x6, Qc67x6;
wire Xc67x6, Ed67x6, Ld67x6, Sd67x6, Zd67x6, Ge67x6, Ne67x6, Ue67x6, Bf67x6, If67x6;
wire Pf67x6, Wf67x6, Dg67x6, Kg67x6, Rg67x6, Yg67x6, Fh67x6, Mh67x6, Th67x6, Ai67x6;
wire Hi67x6, Oi67x6, Vi67x6, Cj67x6, Jj67x6, Qj67x6, Xj67x6, Ek67x6, Lk67x6, Sk67x6;
wire Zk67x6, Gl67x6, Nl67x6, Ul67x6, Bm67x6, Im67x6, Pm67x6, Wm67x6, Dn67x6, Kn67x6;
wire Rn67x6, Yn67x6, Fo67x6, Mo67x6, To67x6, Ap67x6, Hp67x6, Op67x6, Vp67x6, Cq67x6;
wire Jq67x6, Qq67x6, Xq67x6, Er67x6, Lr67x6, Sr67x6, Zr67x6, Gs67x6, Ns67x6, Us67x6;
wire Bt67x6, It67x6, Pt67x6, Wt67x6, Du67x6, Ku67x6, Ru67x6, Yu67x6, Fv67x6, Mv67x6;
wire Tv67x6, Aw67x6, Hw67x6, Ow67x6, Vw67x6, Cx67x6, Jx67x6, Qx67x6, Xx67x6, Ey67x6;
wire Ly67x6, Sy67x6, Zy67x6, Gz67x6, Nz67x6, Uz67x6, B077x6, I077x6, P077x6, W077x6;
wire D177x6, K177x6, R177x6, Y177x6, F277x6, M277x6, T277x6, A377x6, H377x6, O377x6;
wire V377x6, C477x6, J477x6, Q477x6, X477x6, E577x6, L577x6, S577x6, Z577x6, G677x6;
wire N677x6, U677x6, B777x6, I777x6, P777x6, W777x6, D877x6, K877x6, R877x6, Y877x6;
wire F977x6, M977x6, T977x6, Aa77x6, Ha77x6, Oa77x6, Va77x6, Cb77x6, Jb77x6, Qb77x6;
wire Xb77x6, Ec77x6, Lc77x6, Sc77x6, Zc77x6, Gd77x6, Nd77x6, Ud77x6, Be77x6, Ie77x6;
wire Pe77x6, We77x6, Df77x6, Kf77x6, Rf77x6, Yf77x6, Fg77x6, Mg77x6, Tg77x6, Ah77x6;
wire Hh77x6, Oh77x6, Vh77x6, Ci77x6, Ji77x6, Qi77x6, Xi77x6, Ej77x6, Lj77x6, Sj77x6;
wire Zj77x6, Gk77x6, Nk77x6, Uk77x6, Bl77x6, Il77x6, Pl77x6, Wl77x6, Dm77x6, Km77x6;
wire Rm77x6, Ym77x6, Fn77x6, Mn77x6, Tn77x6, Ao77x6, Ho77x6, Oo77x6, Vo77x6, Cp77x6;
wire Jp77x6, Qp77x6, Xp77x6, Eq77x6, Lq77x6, Sq77x6, Zq77x6, Gr77x6, Nr77x6, Ur77x6;
wire Bs77x6, Is77x6, Ps77x6, Ws77x6, Dt77x6, Kt77x6, Rt77x6, Yt77x6, Fu77x6, Mu77x6;
wire Tu77x6, Av77x6, Hv77x6, Ov77x6, Vv77x6, Cw77x6, Jw77x6, Qw77x6, Xw77x6, Ex77x6;
wire Lx77x6, Sx77x6, Zx77x6, Gy77x6, Ny77x6, Uy77x6, Bz77x6, Iz77x6, Pz77x6, Wz77x6;
wire D087x6, K087x6, R087x6, Y087x6, F187x6, M187x6, T187x6, A287x6, H287x6, O287x6;
wire V287x6, C387x6, J387x6, Q387x6, X387x6, E487x6, L487x6, S487x6, Z487x6, G587x6;
wire N587x6, U587x6, B687x6, I687x6, P687x6, W687x6, D787x6, K787x6, R787x6, Y787x6;
wire F887x6, M887x6, T887x6, A987x6, H987x6, O987x6, V987x6, Ca87x6, Ja87x6, Qa87x6;
wire Xa87x6, Eb87x6, Lb87x6, Sb87x6, Zb87x6, Gc87x6, Nc87x6, Uc87x6, Bd87x6, Id87x6;
wire Pd87x6, Wd87x6, De87x6, Ke87x6, Re87x6, Ye87x6, Ff87x6, Mf87x6, Tf87x6, Ag87x6;
wire Hg87x6, Og87x6, Vg87x6, Ch87x6, Jh87x6, Qh87x6, Xh87x6, Ei87x6, Li87x6, Si87x6;
wire Zi87x6, Gj87x6, Nj87x6, Uj87x6, Bk87x6, Ik87x6, Pk87x6, Wk87x6, Dl87x6, Kl87x6;
wire Rl87x6, Yl87x6, Fm87x6, Mm87x6, Tm87x6, An87x6, Hn87x6, On87x6, Vn87x6, Co87x6;
wire Jo87x6, Qo87x6, Xo87x6, Ep87x6, Lp87x6, Sp87x6, Zp87x6, Gq87x6, Nq87x6, Uq87x6;
wire Br87x6, Ir87x6, Pr87x6, Wr87x6, Ds87x6, Ks87x6, Rs87x6, Ys87x6, Ft87x6, Mt87x6;
wire Tt87x6, Au87x6, Hu87x6, Ou87x6, Vu87x6, Cv87x6, Jv87x6, Qv87x6, Xv87x6, Ew87x6;
wire Lw87x6, Sw87x6, Zw87x6, Gx87x6, Nx87x6, Ux87x6, By87x6, Iy87x6, Py87x6, Wy87x6;
wire Dz87x6, Kz87x6, Rz87x6, Yz87x6, F097x6, M097x6, T097x6, A197x6, H197x6, O197x6;
wire V197x6, C297x6, J297x6, Q297x6, X297x6, E397x6, L397x6, S397x6, Z397x6, G497x6;
wire N497x6, U497x6, B597x6, I597x6, P597x6, W597x6, D697x6, K697x6, R697x6, Y697x6;
wire F797x6, M797x6, T797x6, A897x6, H897x6, O897x6, V897x6, C997x6, J997x6, Q997x6;
wire X997x6, Ea97x6, La97x6, Sa97x6, Za97x6, Gb97x6, Nb97x6, Ub97x6, Bc97x6, Ic97x6;
wire Pc97x6, Wc97x6, Dd97x6, Kd97x6, Rd97x6, Yd97x6, Fe97x6, Me97x6, Te97x6, Af97x6;
wire Hf97x6, Of97x6, Vf97x6, Cg97x6, Jg97x6, Qg97x6, Xg97x6, Eh97x6, Lh97x6, Sh97x6;
wire Zh97x6, Gi97x6, Ni97x6, Ui97x6, Bj97x6, Ij97x6, Pj97x6, Wj97x6, Dk97x6, Kk97x6;
wire Rk97x6, Yk97x6, Fl97x6, Ml97x6, Tl97x6, Am97x6, Hm97x6, Om97x6, Vm97x6, Cn97x6;
wire Jn97x6, Qn97x6, Xn97x6, Eo97x6, Lo97x6, So97x6, Zo97x6, Gp97x6, Np97x6, Up97x6;
wire Bq97x6, Iq97x6, Pq97x6, Wq97x6, Dr97x6, Kr97x6, Rr97x6, Yr97x6, Fs97x6, Ms97x6;
wire Ts97x6, At97x6, Ht97x6, Ot97x6, Vt97x6, Cu97x6, Ju97x6, Qu97x6, Xu97x6, Ev97x6;
wire Lv97x6, Sv97x6, Zv97x6, Gw97x6, Nw97x6, Uw97x6, Bx97x6, Ix97x6, Px97x6, Wx97x6;
wire Dy97x6, Ky97x6, Ry97x6, Yy97x6, Fz97x6, Mz97x6, Tz97x6, A0a7x6, H0a7x6, O0a7x6;
wire V0a7x6, C1a7x6, J1a7x6, Q1a7x6, X1a7x6, E2a7x6, L2a7x6, S2a7x6, Z2a7x6, G3a7x6;
wire N3a7x6, U3a7x6, B4a7x6, I4a7x6, P4a7x6, W4a7x6, D5a7x6, K5a7x6, R5a7x6, Y5a7x6;
wire F6a7x6, M6a7x6, T6a7x6, A7a7x6, H7a7x6, O7a7x6, V7a7x6, C8a7x6, J8a7x6, Q8a7x6;
wire X8a7x6, E9a7x6, L9a7x6, S9a7x6, Z9a7x6, Gaa7x6, Naa7x6, Uaa7x6, Bba7x6, Iba7x6;
wire Pba7x6, Wba7x6, Dca7x6, Kca7x6, Rca7x6, Yca7x6, Fda7x6, Mda7x6, Tda7x6, Aea7x6;
wire Hea7x6, Oea7x6, Vea7x6, Cfa7x6, Jfa7x6, Qfa7x6, Xfa7x6, Ega7x6, Lga7x6, Sga7x6;
wire Zga7x6, Gha7x6, Nha7x6, Uha7x6, Bia7x6, Iia7x6, Pia7x6, Wia7x6, Dja7x6, Kja7x6;
wire Rja7x6, Yja7x6, Fka7x6, Mka7x6, Tka7x6, Ala7x6, Hla7x6, Ola7x6, Vla7x6, Cma7x6;
wire Jma7x6, Qma7x6, Xma7x6, Ena7x6, Lna7x6, Sna7x6, Zna7x6, Goa7x6, Noa7x6, Uoa7x6;
wire Bpa7x6, Ipa7x6, Ppa7x6, Wpa7x6, Dqa7x6, Kqa7x6, Rqa7x6, Yqa7x6, Fra7x6, Mra7x6;
wire Tra7x6, Asa7x6, Hsa7x6, Osa7x6, Vsa7x6, Cta7x6, Jta7x6, Qta7x6, Xta7x6, Eua7x6;
wire Lua7x6, Sua7x6, Zua7x6, Gva7x6, Nva7x6, Uva7x6, Bwa7x6, Iwa7x6, Pwa7x6, Wwa7x6;
wire Dxa7x6, Kxa7x6, Rxa7x6, Yxa7x6, Fya7x6, Mya7x6, Tya7x6, Aza7x6, Hza7x6, Oza7x6;
wire Vza7x6, C0b7x6, J0b7x6, Q0b7x6, X0b7x6, E1b7x6, L1b7x6, S1b7x6, Z1b7x6, G2b7x6;
wire N2b7x6, U2b7x6, B3b7x6, I3b7x6, P3b7x6, W3b7x6, D4b7x6, K4b7x6, R4b7x6, Y4b7x6;
wire F5b7x6, M5b7x6, T5b7x6, A6b7x6, H6b7x6, O6b7x6, V6b7x6, C7b7x6, J7b7x6, Q7b7x6;
wire X7b7x6, E8b7x6, L8b7x6, S8b7x6, Z8b7x6, G9b7x6, N9b7x6, U9b7x6, Bab7x6, Iab7x6;
wire Pab7x6, Wab7x6, Dbb7x6, Kbb7x6, Rbb7x6, Ybb7x6, Fcb7x6, Mcb7x6, Tcb7x6, Adb7x6;
wire Hdb7x6, Odb7x6, Vdb7x6, Ceb7x6, Jeb7x6, Qeb7x6, Xeb7x6, Efb7x6, Lfb7x6, Sfb7x6;
wire Zfb7x6, Ggb7x6, Ngb7x6, Ugb7x6, Bhb7x6, Ihb7x6, Phb7x6, Whb7x6, Dib7x6, Kib7x6;
wire Rib7x6, Yib7x6, Fjb7x6, Mjb7x6, Tjb7x6, Akb7x6, Hkb7x6, Okb7x6, Vkb7x6, Clb7x6;
wire Jlb7x6, Qlb7x6, Xlb7x6, Emb7x6, Lmb7x6, Smb7x6, Zmb7x6, Gnb7x6, Nnb7x6, Unb7x6;
wire Bob7x6, Iob7x6, Pob7x6, Wob7x6, Dpb7x6, Kpb7x6, Rpb7x6, Ypb7x6, Fqb7x6, Mqb7x6;
wire Tqb7x6, Arb7x6, Hrb7x6, Orb7x6, Vrb7x6, Csb7x6, Jsb7x6, Qsb7x6, Xsb7x6, Etb7x6;
wire Ltb7x6, Stb7x6, Ztb7x6, Gub7x6, Nub7x6, Uub7x6, Bvb7x6, Ivb7x6, Pvb7x6, Wvb7x6;
wire Dwb7x6, Kwb7x6, Rwb7x6, Ywb7x6, Fxb7x6, Mxb7x6, Txb7x6, Ayb7x6, Hyb7x6, Oyb7x6;
wire Vyb7x6, Czb7x6, Jzb7x6, Qzb7x6, Xzb7x6, E0c7x6, L0c7x6, S0c7x6, Z0c7x6, G1c7x6;
wire N1c7x6, U1c7x6, B2c7x6, I2c7x6, P2c7x6, W2c7x6, D3c7x6, K3c7x6, R3c7x6, Y3c7x6;
wire F4c7x6, M4c7x6, T4c7x6, A5c7x6, H5c7x6, O5c7x6, V5c7x6, C6c7x6, J6c7x6, Q6c7x6;
wire X6c7x6, E7c7x6, L7c7x6, S7c7x6, Z7c7x6, G8c7x6, N8c7x6, U8c7x6, B9c7x6, I9c7x6;
wire P9c7x6, W9c7x6, Dac7x6, Kac7x6, Rac7x6, Yac7x6, Fbc7x6, Mbc7x6, Tbc7x6, Acc7x6;
wire Hcc7x6, Occ7x6, Vcc7x6, Cdc7x6, Jdc7x6, Qdc7x6, Xdc7x6, Eec7x6, Lec7x6, Sec7x6;
wire Zec7x6, Gfc7x6, Nfc7x6, Ufc7x6, Bgc7x6, Igc7x6, Pgc7x6, Wgc7x6, Dhc7x6, Khc7x6;
wire Rhc7x6, Yhc7x6, Fic7x6, Mic7x6, Tic7x6, Ajc7x6, Hjc7x6, Ojc7x6, Vjc7x6, Ckc7x6;
wire Jkc7x6, Qkc7x6, Xkc7x6, Elc7x6, Llc7x6, Slc7x6, Zlc7x6, Gmc7x6, Nmc7x6, Umc7x6;
wire Bnc7x6, Inc7x6, Pnc7x6, Wnc7x6, Doc7x6, Koc7x6, Roc7x6, Yoc7x6, Fpc7x6, Mpc7x6;
wire Tpc7x6, Aqc7x6, Hqc7x6, Oqc7x6, Vqc7x6, Crc7x6, Jrc7x6, Qrc7x6, Xrc7x6, Esc7x6;
wire Lsc7x6, Ssc7x6, Zsc7x6, Gtc7x6, Ntc7x6, Utc7x6, Buc7x6, Iuc7x6, Puc7x6, Wuc7x6;
wire Dvc7x6, Kvc7x6, Rvc7x6, Yvc7x6, Fwc7x6, Mwc7x6, Twc7x6, Axc7x6, Hxc7x6, Oxc7x6;
wire Vxc7x6, Cyc7x6, Jyc7x6, Qyc7x6, Xyc7x6, Ezc7x6, Lzc7x6, Szc7x6, Zzc7x6, G0d7x6;
wire N0d7x6, U0d7x6, B1d7x6, I1d7x6, P1d7x6, W1d7x6, D2d7x6, K2d7x6, R2d7x6, Y2d7x6;
wire F3d7x6, M3d7x6, T3d7x6, A4d7x6, H4d7x6, O4d7x6, V4d7x6, C5d7x6, J5d7x6, Q5d7x6;
wire X5d7x6, E6d7x6, L6d7x6, S6d7x6, Z6d7x6, G7d7x6, N7d7x6, U7d7x6, B8d7x6, I8d7x6;
wire P8d7x6, W8d7x6, D9d7x6, K9d7x6, R9d7x6, Y9d7x6, Fad7x6, Mad7x6, Tad7x6, Abd7x6;
wire Hbd7x6, Obd7x6, Vbd7x6, Ccd7x6, Jcd7x6, Qcd7x6, Xcd7x6, Edd7x6, Ldd7x6, Sdd7x6;
wire Zdd7x6, Ged7x6, Ned7x6, Ued7x6, Bfd7x6, Ifd7x6, Pfd7x6, Wfd7x6, Dgd7x6, Kgd7x6;
wire Rgd7x6, Ygd7x6, Fhd7x6, Mhd7x6, Thd7x6, Aid7x6, Hid7x6, Oid7x6, Vid7x6, Cjd7x6;
wire Jjd7x6, Qjd7x6, Xjd7x6, Ekd7x6, Lkd7x6, Skd7x6, Zkd7x6, Gld7x6, Nld7x6, Uld7x6;
wire Bmd7x6, Imd7x6, Pmd7x6, Wmd7x6, Dnd7x6, Knd7x6, Rnd7x6, Ynd7x6, Fod7x6, Mod7x6;
wire Tod7x6, Apd7x6, Hpd7x6, Opd7x6, Vpd7x6, Cqd7x6, Jqd7x6, Qqd7x6, Xqd7x6, Erd7x6;
wire Lrd7x6, Srd7x6, Zrd7x6, Gsd7x6, Nsd7x6, Usd7x6, Btd7x6, Itd7x6, Ptd7x6, Wtd7x6;
wire Dud7x6, Kud7x6, Rud7x6, Yud7x6, Fvd7x6, Mvd7x6, Tvd7x6, Awd7x6, Hwd7x6, Owd7x6;
wire Vwd7x6, Cxd7x6, Jxd7x6, Qxd7x6, Xxd7x6, Eyd7x6, Lyd7x6, Syd7x6, Zyd7x6, Gzd7x6;
wire Nzd7x6, Uzd7x6, B0e7x6, I0e7x6, P0e7x6, W0e7x6, D1e7x6, K1e7x6, R1e7x6, Y1e7x6;
wire F2e7x6, M2e7x6, T2e7x6, A3e7x6, H3e7x6, O3e7x6, V3e7x6, C4e7x6, J4e7x6, Q4e7x6;
wire X4e7x6, E5e7x6, L5e7x6, S5e7x6, Z5e7x6, G6e7x6, N6e7x6, U6e7x6, B7e7x6, I7e7x6;
wire P7e7x6, W7e7x6, D8e7x6, K8e7x6, R8e7x6, Y8e7x6, F9e7x6, M9e7x6, T9e7x6, Aae7x6;
wire Hae7x6, Oae7x6, Vae7x6, Cbe7x6, Jbe7x6, Qbe7x6, Xbe7x6, Ece7x6, Lce7x6, Sce7x6;
wire Zce7x6, Gde7x6, Nde7x6, Ude7x6, Bee7x6, Iee7x6, Pee7x6, Wee7x6, Dfe7x6, Kfe7x6;
wire Rfe7x6, Yfe7x6, Fge7x6, Mge7x6, Tge7x6, Ahe7x6, Hhe7x6, Ohe7x6, Vhe7x6, Cie7x6;
wire Jie7x6, Qie7x6, Xie7x6, Eje7x6, Lje7x6, Sje7x6, Zje7x6, Gke7x6, Nke7x6, Uke7x6;
wire Ble7x6, Ile7x6, Ple7x6, Wle7x6, Dme7x6, Kme7x6, Rme7x6, Yme7x6, Fne7x6, Mne7x6;
wire Tne7x6, Aoe7x6, Hoe7x6, Ooe7x6, Voe7x6, Cpe7x6, Jpe7x6, Qpe7x6, Xpe7x6, Eqe7x6;
wire Lqe7x6, Sqe7x6, Zqe7x6, Gre7x6, Nre7x6, Ure7x6, Bse7x6, Ise7x6, Pse7x6, Wse7x6;
wire Dte7x6, Kte7x6, Rte7x6, Yte7x6, Fue7x6, Mue7x6, Tue7x6, Ave7x6, Hve7x6, Ove7x6;
wire Vve7x6, Cwe7x6, Jwe7x6, Qwe7x6, Xwe7x6, Exe7x6, Lxe7x6, Sxe7x6, Zxe7x6, Gye7x6;
wire Nye7x6, Uye7x6, Bze7x6, Ize7x6, Pze7x6, Wze7x6, D0f7x6, K0f7x6, R0f7x6, Y0f7x6;
wire F1f7x6, M1f7x6, T1f7x6, A2f7x6, H2f7x6, O2f7x6, V2f7x6, C3f7x6, J3f7x6, Q3f7x6;
wire X3f7x6, E4f7x6, L4f7x6, S4f7x6, Z4f7x6, G5f7x6, N5f7x6, U5f7x6, B6f7x6, I6f7x6;
wire P6f7x6, W6f7x6, D7f7x6, K7f7x6, R7f7x6, Y7f7x6, F8f7x6, M8f7x6, T8f7x6, A9f7x6;
wire H9f7x6, O9f7x6, V9f7x6, Caf7x6, Jaf7x6, Qaf7x6, Xaf7x6, Ebf7x6, Lbf7x6, Sbf7x6;
wire Zbf7x6, Gcf7x6, Ncf7x6, Ucf7x6, Bdf7x6, Idf7x6, Pdf7x6, Wdf7x6, Def7x6, Kef7x6;
wire Ref7x6, Yef7x6, Fff7x6, Mff7x6, Tff7x6, Agf7x6, Hgf7x6, Ogf7x6, Vgf7x6, Chf7x6;
wire Jhf7x6, Qhf7x6, Xhf7x6, Eif7x6, Lif7x6, Sif7x6, Zif7x6, Gjf7x6, Njf7x6, Ujf7x6;
wire Bkf7x6, Ikf7x6, Pkf7x6, Wkf7x6, Dlf7x6, Klf7x6, Rlf7x6, Ylf7x6, Fmf7x6, Mmf7x6;
wire Tmf7x6, Anf7x6, Hnf7x6, Onf7x6, Vnf7x6, Cof7x6, Jof7x6, Qof7x6, Xof7x6, Epf7x6;
wire Lpf7x6, Spf7x6, Zpf7x6, Gqf7x6, Nqf7x6, Uqf7x6, Brf7x6, Irf7x6, Prf7x6, Wrf7x6;
wire Dsf7x6, Ksf7x6, Rsf7x6, Ysf7x6, Ftf7x6, Mtf7x6, Ttf7x6, Auf7x6, Huf7x6, Ouf7x6;
wire Vuf7x6, Cvf7x6, Jvf7x6, Qvf7x6, Xvf7x6, Ewf7x6, Lwf7x6, Swf7x6, Zwf7x6, Gxf7x6;
wire Nxf7x6, Uxf7x6, Byf7x6, Iyf7x6, Pyf7x6, Wyf7x6, Dzf7x6, Kzf7x6, Rzf7x6, Yzf7x6;
wire F0g7x6, M0g7x6, T0g7x6, A1g7x6, H1g7x6, O1g7x6, V1g7x6, C2g7x6, J2g7x6, Q2g7x6;
wire X2g7x6, E3g7x6, L3g7x6, S3g7x6, Z3g7x6, G4g7x6, N4g7x6, U4g7x6, B5g7x6, I5g7x6;
wire P5g7x6, W5g7x6, D6g7x6, K6g7x6, R6g7x6, Y6g7x6, F7g7x6, M7g7x6, T7g7x6, A8g7x6;
wire H8g7x6, O8g7x6, V8g7x6, C9g7x6, J9g7x6, Q9g7x6, X9g7x6, Eag7x6, Lag7x6, Sag7x6;
wire Zag7x6, Gbg7x6, Nbg7x6, Ubg7x6, Bcg7x6, Icg7x6, Pcg7x6, Wcg7x6, Ddg7x6, Kdg7x6;
wire Rdg7x6, Ydg7x6, Feg7x6, Meg7x6, Teg7x6, Afg7x6, Hfg7x6, Ofg7x6, Vfg7x6, Cgg7x6;
wire Jgg7x6, Qgg7x6, Xgg7x6, Ehg7x6, Lhg7x6, Shg7x6, Zhg7x6, Gig7x6, Nig7x6, Uig7x6;
wire Bjg7x6, Ijg7x6, Pjg7x6, Wjg7x6, Dkg7x6, Kkg7x6, Rkg7x6, Ykg7x6, Flg7x6, Mlg7x6;
wire Tlg7x6, Amg7x6, Hmg7x6, Omg7x6, Vmg7x6, Cng7x6, Jng7x6, Qng7x6, Xng7x6, Eog7x6;
wire Log7x6, Sog7x6, Zog7x6, Gpg7x6, Npg7x6, Upg7x6, Bqg7x6, Iqg7x6, Pqg7x6, Wqg7x6;
wire Drg7x6, Krg7x6, Rrg7x6, Yrg7x6, Fsg7x6, Msg7x6, Tsg7x6, Atg7x6, Htg7x6, Otg7x6;
wire Vtg7x6, Cug7x6, Jug7x6, Qug7x6, Xug7x6, Evg7x6, Lvg7x6, Svg7x6, Zvg7x6, Gwg7x6;
wire Nwg7x6, Uwg7x6, Bxg7x6, Ixg7x6, Pxg7x6, Wxg7x6, Dyg7x6, Kyg7x6, Ryg7x6, Yyg7x6;
wire Fzg7x6, Mzg7x6, Tzg7x6, A0h7x6, H0h7x6, O0h7x6, V0h7x6, C1h7x6, J1h7x6, Q1h7x6;
wire X1h7x6, E2h7x6, L2h7x6, S2h7x6, Z2h7x6, G3h7x6, N3h7x6, U3h7x6, B4h7x6, I4h7x6;
wire P4h7x6, W4h7x6, D5h7x6, K5h7x6, R5h7x6, Y5h7x6, F6h7x6, M6h7x6, T6h7x6, A7h7x6;
wire H7h7x6, O7h7x6, V7h7x6, C8h7x6, J8h7x6, Q8h7x6, X8h7x6, E9h7x6, L9h7x6, S9h7x6;
wire Z9h7x6, Gah7x6, Nah7x6, Uah7x6, Bbh7x6, Ibh7x6, Pbh7x6, Wbh7x6, Dch7x6, Kch7x6;
wire Rch7x6, Ych7x6, Fdh7x6, Mdh7x6, Tdh7x6, Aeh7x6, Heh7x6, Oeh7x6, Veh7x6, Cfh7x6;
wire Jfh7x6, Qfh7x6, Xfh7x6, Egh7x6, Lgh7x6, Sgh7x6, Zgh7x6, Ghh7x6, Nhh7x6, Uhh7x6;
wire Bih7x6, Iih7x6, Pih7x6, Wih7x6, Djh7x6, Kjh7x6, Rjh7x6, Yjh7x6, Fkh7x6, Mkh7x6;
wire Tkh7x6, Alh7x6, Hlh7x6, Olh7x6, Vlh7x6, Cmh7x6, Jmh7x6, Qmh7x6, Xmh7x6, Enh7x6;
wire Lnh7x6, Snh7x6, Znh7x6, Goh7x6, Noh7x6, Uoh7x6, Bph7x6, Iph7x6, Pph7x6, Wph7x6;
wire Dqh7x6, Kqh7x6, Rqh7x6, Yqh7x6, Frh7x6, Mrh7x6, Trh7x6, Ash7x6, Hsh7x6, Osh7x6;
wire Vsh7x6, Cth7x6, Jth7x6, Qth7x6, Xth7x6, Euh7x6, Luh7x6, Suh7x6, Zuh7x6, Gvh7x6;
wire Nvh7x6, Uvh7x6, Bwh7x6, Iwh7x6, Pwh7x6, Wwh7x6, Dxh7x6, Kxh7x6, Rxh7x6, Yxh7x6;
wire Fyh7x6, Myh7x6, Tyh7x6, Azh7x6, Hzh7x6, Ozh7x6, Vzh7x6, C0i7x6, J0i7x6, Q0i7x6;
wire X0i7x6, E1i7x6, L1i7x6, S1i7x6, Z1i7x6, G2i7x6, N2i7x6, U2i7x6, B3i7x6, I3i7x6;
wire P3i7x6, W3i7x6, D4i7x6, K4i7x6, R4i7x6, Y4i7x6, F5i7x6, M5i7x6, T5i7x6, A6i7x6;
wire H6i7x6, O6i7x6, V6i7x6, C7i7x6, J7i7x6, Q7i7x6, X7i7x6, E8i7x6, L8i7x6, S8i7x6;
wire Z8i7x6, G9i7x6, N9i7x6, U9i7x6, Bai7x6, Iai7x6, Pai7x6, Wai7x6, Dbi7x6, Kbi7x6;
wire Rbi7x6, Ybi7x6, Fci7x6, Mci7x6, Tci7x6, Adi7x6, Hdi7x6, Odi7x6, Vdi7x6, Cei7x6;
wire Jei7x6, Qei7x6, Xei7x6, Efi7x6, Lfi7x6, Sfi7x6, Zfi7x6, Ggi7x6, Ngi7x6, Ugi7x6;
wire Bhi7x6, Ihi7x6, Phi7x6, Whi7x6, Dii7x6, Kii7x6, Rii7x6, Yii7x6, Fji7x6, Mji7x6;
wire Tji7x6, Aki7x6, Hki7x6, Oki7x6, Vki7x6, Cli7x6, Jli7x6, Qli7x6, Xli7x6, Emi7x6;
wire Lmi7x6, Smi7x6, Zmi7x6, Gni7x6, Nni7x6, Uni7x6, Boi7x6, Ioi7x6, Poi7x6, Woi7x6;
wire Dpi7x6, Kpi7x6, Rpi7x6, Ypi7x6, Fqi7x6, Mqi7x6, Tqi7x6, Ari7x6, Hri7x6, Ori7x6;
wire Vri7x6, Csi7x6, Jsi7x6, Qsi7x6, Xsi7x6, Eti7x6, Lti7x6, Sti7x6, Zti7x6, Gui7x6;
wire Nui7x6, Uui7x6, Bvi7x6, Ivi7x6, Pvi7x6, Wvi7x6, Dwi7x6, Kwi7x6, Rwi7x6, Ywi7x6;
wire Fxi7x6, Mxi7x6, Txi7x6, Ayi7x6, Hyi7x6, Oyi7x6, Vyi7x6, Czi7x6, Jzi7x6, Qzi7x6;
wire Xzi7x6, E0j7x6, L0j7x6, S0j7x6, Z0j7x6, G1j7x6, N1j7x6, U1j7x6, B2j7x6, I2j7x6;
wire P2j7x6, W2j7x6, D3j7x6, K3j7x6, R3j7x6, Y3j7x6, F4j7x6, M4j7x6, T4j7x6, A5j7x6;
wire H5j7x6, O5j7x6, V5j7x6, C6j7x6, J6j7x6, Q6j7x6, X6j7x6, E7j7x6, L7j7x6, S7j7x6;
wire Z7j7x6, G8j7x6, N8j7x6, U8j7x6, B9j7x6, I9j7x6, P9j7x6, W9j7x6, Daj7x6, Kaj7x6;
wire Raj7x6, Yaj7x6, Fbj7x6, Mbj7x6, Tbj7x6, Acj7x6, Hcj7x6, Ocj7x6, Vcj7x6, Cdj7x6;
wire Jdj7x6, Qdj7x6, Xdj7x6, Eej7x6, Lej7x6, Sej7x6, Zej7x6, Gfj7x6, Nfj7x6, Ufj7x6;
wire Bgj7x6, Igj7x6, Pgj7x6, Wgj7x6, Dhj7x6, Khj7x6, Rhj7x6, Yhj7x6, Fij7x6, Mij7x6;
wire Tij7x6, Ajj7x6, Hjj7x6, Ojj7x6, Vjj7x6, Ckj7x6, Jkj7x6, Qkj7x6, Xkj7x6, Elj7x6;
wire Llj7x6, Slj7x6, Zlj7x6, Gmj7x6, Nmj7x6, Umj7x6, Bnj7x6, Inj7x6, Pnj7x6, Wnj7x6;
wire Doj7x6, Koj7x6, Roj7x6, Yoj7x6, Fpj7x6, Mpj7x6, Tpj7x6, Aqj7x6, Hqj7x6, Oqj7x6;
wire Vqj7x6, Crj7x6, Jrj7x6, Qrj7x6, Xrj7x6, Esj7x6, Lsj7x6, Ssj7x6, Zsj7x6, Gtj7x6;
wire Ntj7x6, Utj7x6, Buj7x6, Iuj7x6, Puj7x6, Wuj7x6, Dvj7x6, Kvj7x6, Rvj7x6, Yvj7x6;
wire Fwj7x6, Mwj7x6, Twj7x6, Axj7x6, Hxj7x6, Oxj7x6, Vxj7x6, Cyj7x6, Jyj7x6, Qyj7x6;
wire Xyj7x6, Ezj7x6, Lzj7x6, Szj7x6, Zzj7x6, G0k7x6, N0k7x6, U0k7x6, B1k7x6, I1k7x6;
wire P1k7x6, W1k7x6, D2k7x6, K2k7x6, R2k7x6, Y2k7x6, F3k7x6, M3k7x6, T3k7x6, A4k7x6;
wire H4k7x6, O4k7x6, V4k7x6, C5k7x6, J5k7x6, Q5k7x6, X5k7x6, E6k7x6, L6k7x6, S6k7x6;
wire Z6k7x6, G7k7x6, N7k7x6, U7k7x6, B8k7x6, I8k7x6, P8k7x6, W8k7x6, D9k7x6, K9k7x6;
wire R9k7x6, Y9k7x6, Fak7x6, Mak7x6, Tak7x6, Abk7x6, Hbk7x6, Obk7x6, Vbk7x6, Cck7x6;
wire Jck7x6, Qck7x6, Xck7x6, Edk7x6, Ldk7x6, Sdk7x6, Zdk7x6, Gek7x6, Nek7x6, Uek7x6;
wire Bfk7x6, Ifk7x6, Pfk7x6, Wfk7x6, Dgk7x6, Kgk7x6, Rgk7x6, Ygk7x6, Fhk7x6, Mhk7x6;
wire Thk7x6, Aik7x6, Hik7x6, Oik7x6, Vik7x6, Cjk7x6, Jjk7x6, Qjk7x6, Xjk7x6, Ekk7x6;
wire Lkk7x6, Skk7x6, Zkk7x6, Glk7x6, Nlk7x6, Ulk7x6, Bmk7x6, Imk7x6, Pmk7x6, Wmk7x6;
wire Dnk7x6, Knk7x6, Rnk7x6, Ynk7x6, Fok7x6, Mok7x6, Tok7x6, Apk7x6, Hpk7x6, Opk7x6;
wire Vpk7x6, Cqk7x6, Jqk7x6, Qqk7x6, Xqk7x6, Erk7x6, Lrk7x6, Srk7x6, Zrk7x6, Gsk7x6;
wire Nsk7x6, Usk7x6, Btk7x6, Itk7x6, Ptk7x6, Wtk7x6, Duk7x6, Kuk7x6, Ruk7x6, Yuk7x6;
wire Fvk7x6, Mvk7x6, Tvk7x6, Awk7x6, Hwk7x6, Owk7x6, Vwk7x6, Cxk7x6, Jxk7x6, Qxk7x6;
wire Xxk7x6, Eyk7x6, Lyk7x6, Syk7x6, Zyk7x6, Gzk7x6, Nzk7x6, Uzk7x6, B0l7x6, I0l7x6;
wire P0l7x6, W0l7x6, D1l7x6, K1l7x6, R1l7x6, Y1l7x6, F2l7x6, M2l7x6, T2l7x6, A3l7x6;
wire H3l7x6, O3l7x6, V3l7x6, C4l7x6, J4l7x6, Q4l7x6, X4l7x6, E5l7x6, L5l7x6, S5l7x6;
wire Z5l7x6, G6l7x6, N6l7x6, U6l7x6, B7l7x6, I7l7x6, P7l7x6, W7l7x6, D8l7x6, K8l7x6;
wire R8l7x6, Y8l7x6, F9l7x6, M9l7x6, T9l7x6, Aal7x6, Hal7x6, Oal7x6, Val7x6, Cbl7x6;
wire Jbl7x6, Qbl7x6, Xbl7x6, Ecl7x6, Lcl7x6, Scl7x6, Zcl7x6, Gdl7x6, Ndl7x6, Udl7x6;
wire Bel7x6, Iel7x6, Pel7x6, Wel7x6, Dfl7x6, Kfl7x6, Rfl7x6, Yfl7x6, Fgl7x6, Mgl7x6;
wire Tgl7x6, Ahl7x6, Hhl7x6, Ohl7x6, Vhl7x6, Cil7x6, Jil7x6, Qil7x6, Xil7x6, Ejl7x6;
wire Ljl7x6, Sjl7x6, Zjl7x6, Gkl7x6, Nkl7x6, Ukl7x6, Bll7x6, Ill7x6, Pll7x6, Wll7x6;
wire Dml7x6, Kml7x6, Rml7x6, Yml7x6, Fnl7x6, Mnl7x6, Tnl7x6, Aol7x6, Hol7x6, Ool7x6;
wire Vol7x6, Cpl7x6, Jpl7x6, Qpl7x6, Xpl7x6, Eql7x6, Lql7x6, Sql7x6, Zql7x6, Grl7x6;
wire Nrl7x6, Url7x6, Bsl7x6, Isl7x6, Psl7x6, Wsl7x6, Dtl7x6, Ktl7x6, Rtl7x6, Ytl7x6;
wire Ful7x6, Mul7x6, Tul7x6, Avl7x6, Hvl7x6, Ovl7x6, Vvl7x6, Cwl7x6, Jwl7x6, Qwl7x6;
wire Xwl7x6, Exl7x6, Lxl7x6, Sxl7x6, Zxl7x6, Gyl7x6, Nyl7x6, Uyl7x6, Bzl7x6, Izl7x6;
wire Pzl7x6, Wzl7x6, D0m7x6, K0m7x6, R0m7x6, Y0m7x6, F1m7x6, M1m7x6, T1m7x6, A2m7x6;
wire H2m7x6, O2m7x6, V2m7x6, C3m7x6, J3m7x6, Q3m7x6, X3m7x6, E4m7x6, L4m7x6, S4m7x6;
wire Z4m7x6, G5m7x6, N5m7x6, U5m7x6, B6m7x6, I6m7x6, P6m7x6, W6m7x6, D7m7x6, K7m7x6;
wire R7m7x6, Y7m7x6, F8m7x6, M8m7x6, T8m7x6, A9m7x6, H9m7x6, O9m7x6, V9m7x6, Cam7x6;
wire Jam7x6, Qam7x6, Xam7x6, Ebm7x6, Lbm7x6, Sbm7x6, Zbm7x6, Gcm7x6, Ncm7x6, Ucm7x6;
wire Bdm7x6, Idm7x6, Pdm7x6, Wdm7x6, Dem7x6, Kem7x6, Rem7x6, Yem7x6, Ffm7x6, Mfm7x6;
wire Tfm7x6, Agm7x6, Hgm7x6, Ogm7x6, Vgm7x6, Chm7x6, Jhm7x6, Qhm7x6, Xhm7x6, Eim7x6;
wire Lim7x6, Sim7x6, Zim7x6, Gjm7x6, Njm7x6, Ujm7x6, Bkm7x6, Ikm7x6, Pkm7x6, Wkm7x6;
wire Dlm7x6, Klm7x6, Rlm7x6, Ylm7x6, Fmm7x6, Mmm7x6, Tmm7x6, Anm7x6, Hnm7x6, Onm7x6;
wire Vnm7x6, Com7x6, Jom7x6, Qom7x6, Xom7x6, Epm7x6, Lpm7x6, Spm7x6, Zpm7x6, Gqm7x6;
wire Nqm7x6, Uqm7x6, Brm7x6, Irm7x6, Prm7x6, Wrm7x6, Dsm7x6, Ksm7x6, Rsm7x6, Ysm7x6;
wire Ftm7x6, Mtm7x6, Ttm7x6, Aum7x6, Hum7x6, Oum7x6, Vum7x6, Cvm7x6, Jvm7x6, Qvm7x6;
wire Xvm7x6, Ewm7x6, Lwm7x6, Swm7x6, Zwm7x6, Gxm7x6, Nxm7x6, Uxm7x6, Bym7x6, Iym7x6;
wire Pym7x6, Wym7x6, Dzm7x6, Kzm7x6, Rzm7x6, Yzm7x6, F0n7x6, M0n7x6, T0n7x6, A1n7x6;
wire H1n7x6, O1n7x6, V1n7x6, C2n7x6, J2n7x6, Q2n7x6, X2n7x6, E3n7x6, L3n7x6, S3n7x6;
wire Z3n7x6, G4n7x6, N4n7x6, U4n7x6, B5n7x6, I5n7x6, P5n7x6, W5n7x6, D6n7x6, K6n7x6;
wire R6n7x6, Y6n7x6, F7n7x6, M7n7x6, T7n7x6, A8n7x6, H8n7x6, O8n7x6, V8n7x6, C9n7x6;
wire J9n7x6, Q9n7x6, X9n7x6, Ean7x6, Lan7x6, San7x6, Zan7x6, Gbn7x6, Nbn7x6, Ubn7x6;
wire Bcn7x6, Icn7x6, Pcn7x6, Wcn7x6, Ddn7x6, Kdn7x6, Rdn7x6, Ydn7x6, Fen7x6, Men7x6;
wire Ten7x6, Afn7x6, Hfn7x6, Ofn7x6, Vfn7x6, Cgn7x6, Jgn7x6, Qgn7x6, Xgn7x6, Ehn7x6;
wire Lhn7x6, Shn7x6, Zhn7x6, Gin7x6, Nin7x6, Uin7x6, Bjn7x6, Ijn7x6, Pjn7x6, Wjn7x6;
wire Dkn7x6, Kkn7x6, Rkn7x6, Ykn7x6, Fln7x6, Mln7x6, Tln7x6, Amn7x6, Hmn7x6, Omn7x6;
wire Vmn7x6, Cnn7x6, Jnn7x6, Qnn7x6, Xnn7x6, Eon7x6, Lon7x6, Son7x6, Zon7x6, Gpn7x6;
wire Npn7x6, Upn7x6, Bqn7x6, Iqn7x6, Pqn7x6, Wqn7x6, Drn7x6, Krn7x6, Rrn7x6, Yrn7x6;
wire Fsn7x6, Msn7x6, Tsn7x6, Atn7x6, Htn7x6, Otn7x6, Vtn7x6, Cun7x6, Jun7x6, Qun7x6;
wire Xun7x6, Evn7x6, Lvn7x6, Svn7x6, Zvn7x6, Gwn7x6, Nwn7x6, Uwn7x6, Bxn7x6, Ixn7x6;
wire Pxn7x6, Wxn7x6, Dyn7x6, Kyn7x6, Ryn7x6, Yyn7x6, Fzn7x6, Mzn7x6, Tzn7x6, A0o7x6;
wire H0o7x6, O0o7x6, V0o7x6, C1o7x6, J1o7x6, Q1o7x6, X1o7x6, E2o7x6, L2o7x6, S2o7x6;
wire Z2o7x6, G3o7x6, N3o7x6, U3o7x6, B4o7x6, I4o7x6, P4o7x6, W4o7x6, D5o7x6, K5o7x6;
wire R5o7x6, Y5o7x6, F6o7x6, M6o7x6, T6o7x6, A7o7x6, H7o7x6, O7o7x6, V7o7x6, C8o7x6;
wire J8o7x6, Q8o7x6, X8o7x6, E9o7x6, L9o7x6, S9o7x6, Z9o7x6, Gao7x6, Nao7x6, Uao7x6;
wire Bbo7x6, Ibo7x6, Pbo7x6, Wbo7x6, Dco7x6, Kco7x6, Rco7x6, Yco7x6, Fdo7x6, Mdo7x6;
wire Tdo7x6, Aeo7x6, Heo7x6, Oeo7x6, Veo7x6, Cfo7x6, Jfo7x6, Qfo7x6, Xfo7x6, Ego7x6;
wire Lgo7x6, Sgo7x6, Zgo7x6, Gho7x6, Nho7x6, Uho7x6, Bio7x6, Iio7x6, Pio7x6, Wio7x6;
wire Djo7x6, Kjo7x6, Rjo7x6, Yjo7x6, Fko7x6, Mko7x6, Tko7x6, Alo7x6, Hlo7x6, Olo7x6;
wire Vlo7x6, Cmo7x6, Jmo7x6, Qmo7x6, Xmo7x6, Eno7x6, Lno7x6, Sno7x6, Zno7x6, Goo7x6;
wire Noo7x6, Uoo7x6, Bpo7x6, Ipo7x6, Ppo7x6, Wpo7x6, Dqo7x6, Kqo7x6, Rqo7x6, Yqo7x6;
wire Fro7x6, Mro7x6, Tro7x6, Aso7x6, Hso7x6, Oso7x6, Vso7x6, Cto7x6, Jto7x6, Qto7x6;
wire Xto7x6, Euo7x6, Luo7x6, Suo7x6, Zuo7x6, Gvo7x6, Nvo7x6, Uvo7x6, Bwo7x6, Iwo7x6;
wire Pwo7x6, Wwo7x6, Dxo7x6, Kxo7x6, Rxo7x6, Yxo7x6, Fyo7x6, Myo7x6, Tyo7x6, Azo7x6;
wire Hzo7x6, Ozo7x6, Vzo7x6, C0p7x6, J0p7x6, Q0p7x6, X0p7x6, E1p7x6, L1p7x6, S1p7x6;
wire Z1p7x6, G2p7x6, N2p7x6, U2p7x6, B3p7x6, I3p7x6, P3p7x6, W3p7x6, D4p7x6, K4p7x6;
wire R4p7x6, Y4p7x6, F5p7x6, M5p7x6, T5p7x6, A6p7x6, H6p7x6, O6p7x6, V6p7x6, C7p7x6;
wire J7p7x6, Q7p7x6, X7p7x6, E8p7x6, L8p7x6, S8p7x6, Z8p7x6, G9p7x6, N9p7x6, U9p7x6;
wire Bap7x6, Iap7x6, Pap7x6, Wap7x6, Dbp7x6, Kbp7x6, Rbp7x6, Ybp7x6, Fcp7x6, Mcp7x6;
wire Tcp7x6, Adp7x6, Hdp7x6, Odp7x6, Vdp7x6, Cep7x6, Jep7x6, Qep7x6, Xep7x6, Efp7x6;
wire Lfp7x6, Sfp7x6, Zfp7x6, Ggp7x6, Ngp7x6, Ugp7x6, Bhp7x6, Ihp7x6, Php7x6, Whp7x6;
wire Dip7x6, Kip7x6, Rip7x6, Yip7x6, Fjp7x6, Mjp7x6, Tjp7x6, Akp7x6, Hkp7x6, Okp7x6;
wire Vkp7x6, Clp7x6, Jlp7x6, Qlp7x6, Xlp7x6, Emp7x6, Lmp7x6, Smp7x6, Zmp7x6, Gnp7x6;
wire Nnp7x6, Unp7x6, Bop7x6, Iop7x6, Pop7x6, Wop7x6, Dpp7x6, Kpp7x6, Rpp7x6, Ypp7x6;
wire Fqp7x6, Mqp7x6, Tqp7x6, Arp7x6, Hrp7x6, Orp7x6, Vrp7x6, Csp7x6, Jsp7x6, Qsp7x6;
wire Xsp7x6, Etp7x6, Ltp7x6, Stp7x6, Ztp7x6, Gup7x6, Nup7x6, Uup7x6, Bvp7x6, Ivp7x6;
wire Pvp7x6, Wvp7x6, Dwp7x6, Kwp7x6, Rwp7x6, Ywp7x6, Fxp7x6, Mxp7x6, Txp7x6, Ayp7x6;
wire Hyp7x6, Oyp7x6, Vyp7x6, Czp7x6, Jzp7x6, Qzp7x6, Xzp7x6, E0q7x6, L0q7x6, S0q7x6;
wire Z0q7x6, G1q7x6, N1q7x6, U1q7x6, B2q7x6, I2q7x6, P2q7x6, W2q7x6, D3q7x6, K3q7x6;
wire R3q7x6, Y3q7x6, F4q7x6, M4q7x6, T4q7x6, A5q7x6, H5q7x6, O5q7x6, V5q7x6, C6q7x6;
wire J6q7x6, Q6q7x6, X6q7x6, E7q7x6, L7q7x6, S7q7x6, Z7q7x6, G8q7x6, N8q7x6, U8q7x6;
wire B9q7x6, I9q7x6, P9q7x6, W9q7x6, Daq7x6, Kaq7x6, Raq7x6, Yaq7x6, Fbq7x6, Mbq7x6;
wire Tbq7x6, Acq7x6, Hcq7x6, Ocq7x6, Vcq7x6, Cdq7x6, Jdq7x6, Qdq7x6, Xdq7x6, Eeq7x6;
wire Leq7x6, Seq7x6, Zeq7x6, Gfq7x6, Nfq7x6, Ufq7x6, Bgq7x6, Igq7x6, Pgq7x6, Wgq7x6;
wire Dhq7x6, Khq7x6, Rhq7x6, Yhq7x6, Fiq7x6, Miq7x6, Tiq7x6, Ajq7x6, Hjq7x6, Ojq7x6;
wire Vjq7x6, Ckq7x6, Jkq7x6, Qkq7x6, Xkq7x6, Elq7x6, Llq7x6, Slq7x6, Zlq7x6, Gmq7x6;
wire Nmq7x6, Umq7x6, Bnq7x6, Inq7x6, Pnq7x6, Wnq7x6, Doq7x6, Koq7x6, Roq7x6, Yoq7x6;
wire Fpq7x6, Mpq7x6, Tpq7x6, Aqq7x6, Hqq7x6, Oqq7x6, Vqq7x6, Crq7x6, Jrq7x6, Qrq7x6;
wire Xrq7x6, Esq7x6, Lsq7x6, Ssq7x6, Zsq7x6, Gtq7x6, Ntq7x6, Utq7x6, Buq7x6, Iuq7x6;
wire Puq7x6, Wuq7x6, Dvq7x6, Kvq7x6, Rvq7x6, Yvq7x6, Fwq7x6, Mwq7x6, Twq7x6, Axq7x6;
wire Hxq7x6, Oxq7x6, Vxq7x6, Cyq7x6, Jyq7x6, Qyq7x6, Xyq7x6, Ezq7x6, Lzq7x6, Szq7x6;
wire Zzq7x6, G0r7x6, N0r7x6, U0r7x6, B1r7x6, I1r7x6, P1r7x6, W1r7x6, D2r7x6, K2r7x6;
wire R2r7x6, Y2r7x6, F3r7x6, M3r7x6, T3r7x6, A4r7x6, H4r7x6, O4r7x6, V4r7x6, C5r7x6;
wire J5r7x6, Q5r7x6, X5r7x6, E6r7x6, L6r7x6, S6r7x6, Z6r7x6, G7r7x6, N7r7x6, U7r7x6;
wire B8r7x6, I8r7x6, P8r7x6, W8r7x6, D9r7x6, K9r7x6, R9r7x6, Y9r7x6, Far7x6, Mar7x6;
wire Tar7x6, Abr7x6, Hbr7x6, Obr7x6, Vbr7x6, Ccr7x6, Jcr7x6, Qcr7x6, Xcr7x6, Edr7x6;
wire Ldr7x6, Sdr7x6, Zdr7x6, Ger7x6, Ner7x6, Uer7x6, Bfr7x6, Ifr7x6, Pfr7x6, Wfr7x6;
wire Dgr7x6, Kgr7x6, Rgr7x6, Ygr7x6, Fhr7x6, Mhr7x6, Thr7x6, Air7x6, Hir7x6, Oir7x6;
wire Vir7x6, Cjr7x6, Jjr7x6, Qjr7x6, Xjr7x6, Ekr7x6, Lkr7x6, Skr7x6, Zkr7x6, Glr7x6;
wire Nlr7x6, Ulr7x6, Bmr7x6, Imr7x6, Pmr7x6, Wmr7x6, Dnr7x6, Knr7x6, Rnr7x6, Ynr7x6;
wire For7x6, Mor7x6, Tor7x6, Apr7x6, Hpr7x6, Opr7x6, Vpr7x6, Cqr7x6, Jqr7x6, Qqr7x6;
wire Xqr7x6, Err7x6, Lrr7x6, Srr7x6, Zrr7x6, Gsr7x6, Nsr7x6, Usr7x6, Btr7x6, Itr7x6;
wire Ptr7x6, Wtr7x6, Dur7x6, Kur7x6, Rur7x6, Yur7x6, Fvr7x6, Mvr7x6, Tvr7x6, Awr7x6;
wire Hwr7x6, Owr7x6, Vwr7x6, Cxr7x6, Jxr7x6, Qxr7x6, Xxr7x6, Eyr7x6, Lyr7x6, Syr7x6;
wire Zyr7x6, Gzr7x6, Nzr7x6, Uzr7x6, B0s7x6, I0s7x6, P0s7x6, W0s7x6, D1s7x6, K1s7x6;
wire R1s7x6, Y1s7x6, F2s7x6, M2s7x6, T2s7x6, A3s7x6, H3s7x6, O3s7x6, V3s7x6, C4s7x6;
wire J4s7x6, Q4s7x6, X4s7x6, E5s7x6, L5s7x6, S5s7x6, Z5s7x6, G6s7x6, N6s7x6, U6s7x6;
wire B7s7x6, I7s7x6, P7s7x6, W7s7x6, D8s7x6, K8s7x6, R8s7x6, Y8s7x6, F9s7x6, M9s7x6;
wire T9s7x6, Aas7x6, Has7x6, Oas7x6, Vas7x6, Cbs7x6, Jbs7x6, Qbs7x6, Xbs7x6, Ecs7x6;
wire Lcs7x6, Scs7x6, Zcs7x6, Gds7x6, Nds7x6, Uds7x6, Bes7x6, Ies7x6, Pes7x6, Wes7x6;
wire Dfs7x6, Kfs7x6, Rfs7x6, Yfs7x6, Fgs7x6, Mgs7x6, Tgs7x6, Ahs7x6, Hhs7x6, Ohs7x6;
wire Vhs7x6, Cis7x6, Jis7x6, Qis7x6, Xis7x6, Ejs7x6, Ljs7x6, Sjs7x6, Zjs7x6, Gks7x6;
wire Nks7x6, Uks7x6, Bls7x6, Ils7x6, Pls7x6, Wls7x6, Dms7x6, Kms7x6, Rms7x6, Yms7x6;
wire Fns7x6, Mns7x6, Tns7x6, Aos7x6, Hos7x6, Oos7x6, Vos7x6, Cps7x6, Jps7x6, Qps7x6;
wire Xps7x6, Eqs7x6, Lqs7x6, Sqs7x6, Zqs7x6, Grs7x6, Nrs7x6, Urs7x6, Bss7x6, Iss7x6;
wire Pss7x6, Wss7x6, Dts7x6, Kts7x6, Rts7x6, Yts7x6, Fus7x6, Mus7x6, Tus7x6, Avs7x6;
wire Hvs7x6, Ovs7x6, Vvs7x6, Cws7x6, Jws7x6, Qws7x6, Xws7x6, Exs7x6, Lxs7x6, Sxs7x6;
wire Zxs7x6, Gys7x6, Nys7x6, Uys7x6, Bzs7x6, Izs7x6, Pzs7x6, Wzs7x6, D0t7x6, K0t7x6;
wire R0t7x6, Y0t7x6, F1t7x6, M1t7x6, T1t7x6, A2t7x6, H2t7x6, O2t7x6, V2t7x6, C3t7x6;
wire J3t7x6, Q3t7x6, X3t7x6, E4t7x6, L4t7x6, S4t7x6, Z4t7x6, G5t7x6, N5t7x6, U5t7x6;
wire B6t7x6, I6t7x6, P6t7x6, W6t7x6, D7t7x6, K7t7x6, R7t7x6, Y7t7x6, F8t7x6, M8t7x6;
wire T8t7x6, A9t7x6, H9t7x6, O9t7x6, V9t7x6, Cat7x6, Jat7x6, Qat7x6, Xat7x6, Ebt7x6;
wire Lbt7x6, Sbt7x6, Zbt7x6, Gct7x6, Nct7x6, Uct7x6, Bdt7x6, Idt7x6, Pdt7x6, Wdt7x6;
wire Det7x6, Ket7x6, Ret7x6, Yet7x6, Fft7x6, Mft7x6, Tft7x6, Agt7x6, Hgt7x6, Ogt7x6;
wire Vgt7x6, Cht7x6, Jht7x6, Qht7x6, Xht7x6, Eit7x6, Lit7x6, Sit7x6, Zit7x6, Gjt7x6;
wire Njt7x6, Ujt7x6, Bkt7x6, Ikt7x6, Pkt7x6, Wkt7x6, Dlt7x6, Klt7x6, Rlt7x6, Ylt7x6;
wire Fmt7x6, Mmt7x6, Tmt7x6, Ant7x6, Hnt7x6, Ont7x6, Vnt7x6, Cot7x6, Jot7x6, Qot7x6;
wire Xot7x6, Ept7x6, Lpt7x6, Spt7x6, Zpt7x6, Gqt7x6, Nqt7x6, Uqt7x6, Brt7x6, Irt7x6;
wire Prt7x6, Wrt7x6, Dst7x6, Kst7x6, Rst7x6, Yst7x6, Ftt7x6, Mtt7x6, Ttt7x6, Aut7x6;
wire Hut7x6, Out7x6, Vut7x6, Cvt7x6, Jvt7x6, Qvt7x6, Xvt7x6, Ewt7x6, Lwt7x6, Swt7x6;
wire Zwt7x6, Gxt7x6, Nxt7x6, Uxt7x6, Byt7x6, Iyt7x6, Pyt7x6, Wyt7x6, Dzt7x6, Kzt7x6;
wire Rzt7x6, Yzt7x6, F0u7x6, M0u7x6, T0u7x6, A1u7x6, H1u7x6, O1u7x6, V1u7x6, C2u7x6;
wire J2u7x6, Q2u7x6, X2u7x6, E3u7x6, L3u7x6, S3u7x6, Z3u7x6, G4u7x6, N4u7x6, U4u7x6;
wire B5u7x6, I5u7x6, P5u7x6, W5u7x6, D6u7x6, K6u7x6, R6u7x6, Y6u7x6, F7u7x6, M7u7x6;
wire T7u7x6, A8u7x6, H8u7x6, O8u7x6, V8u7x6, C9u7x6, J9u7x6, Q9u7x6, X9u7x6, Eau7x6;
wire Lau7x6, Sau7x6, Zau7x6, Gbu7x6, Nbu7x6, Ubu7x6, Bcu7x6, Icu7x6, Pcu7x6, Wcu7x6;
wire Ddu7x6, Kdu7x6, Rdu7x6, Ydu7x6, Feu7x6, Meu7x6, Teu7x6, Afu7x6, Hfu7x6, Ofu7x6;
wire Vfu7x6, Cgu7x6, Jgu7x6, Qgu7x6, Xgu7x6, Ehu7x6, Lhu7x6, Shu7x6, Zhu7x6, Giu7x6;
wire Niu7x6, Uiu7x6, Bju7x6, Iju7x6, Pju7x6, Wju7x6, Dku7x6, Kku7x6, Rku7x6, Yku7x6;
wire Flu7x6, Mlu7x6, Tlu7x6, Amu7x6, Hmu7x6, Omu7x6, Vmu7x6, Cnu7x6, Jnu7x6, Qnu7x6;
wire Xnu7x6, Eou7x6, Lou7x6, Sou7x6, Zou7x6, Gpu7x6, Npu7x6, Upu7x6, Bqu7x6, Iqu7x6;
wire Pqu7x6, Wqu7x6, Dru7x6, Kru7x6, Rru7x6, Yru7x6, Fsu7x6, Msu7x6, Tsu7x6, Atu7x6;
wire Htu7x6, Otu7x6, Vtu7x6, Cuu7x6, Juu7x6, Quu7x6, Xuu7x6, Evu7x6, Lvu7x6, Svu7x6;
wire Zvu7x6, Gwu7x6, Nwu7x6, Uwu7x6, Bxu7x6, Ixu7x6, Pxu7x6, Wxu7x6, Dyu7x6, Kyu7x6;
wire Ryu7x6, Yyu7x6, Fzu7x6, Mzu7x6, Tzu7x6, A0v7x6, H0v7x6, O0v7x6, V0v7x6, C1v7x6;
wire J1v7x6, Q1v7x6, X1v7x6, E2v7x6, L2v7x6, S2v7x6, Z2v7x6, G3v7x6, N3v7x6, U3v7x6;
wire B4v7x6, I4v7x6, P4v7x6, W4v7x6, D5v7x6, K5v7x6, R5v7x6, Y5v7x6, F6v7x6, M6v7x6;
wire T6v7x6, A7v7x6, H7v7x6, O7v7x6, V7v7x6, C8v7x6, J8v7x6, Q8v7x6, X8v7x6, E9v7x6;
wire L9v7x6, S9v7x6, Z9v7x6, Gav7x6, Nav7x6, Uav7x6, Bbv7x6, Ibv7x6, Pbv7x6, Wbv7x6;
wire Dcv7x6, Kcv7x6, Rcv7x6, Ycv7x6, Fdv7x6, Mdv7x6, Tdv7x6, Aev7x6, Hev7x6, Oev7x6;
wire Vev7x6, Cfv7x6, Jfv7x6, Qfv7x6, Xfv7x6, Egv7x6, Lgv7x6, Sgv7x6, Zgv7x6, Ghv7x6;
wire Nhv7x6, Uhv7x6, Biv7x6, Iiv7x6, Piv7x6, Wiv7x6, Djv7x6, Kjv7x6, Rjv7x6, Yjv7x6;
wire Fkv7x6, Mkv7x6, Tkv7x6, Alv7x6, Hlv7x6, Olv7x6, Vlv7x6, Cmv7x6, Jmv7x6, Qmv7x6;
wire Xmv7x6, Env7x6, Lnv7x6, Snv7x6, Znv7x6, Gov7x6, Nov7x6, Uov7x6, Bpv7x6, Ipv7x6;
wire Ppv7x6, Wpv7x6, Dqv7x6, Kqv7x6, Rqv7x6, Yqv7x6, Frv7x6, Mrv7x6, Trv7x6, Asv7x6;
wire Hsv7x6, Osv7x6, Vsv7x6, Ctv7x6, Jtv7x6, Qtv7x6, Xtv7x6, Euv7x6, Luv7x6, Suv7x6;
wire Zuv7x6, Gvv7x6, Nvv7x6, Uvv7x6, Bwv7x6, Iwv7x6, Pwv7x6, Wwv7x6, Dxv7x6, Kxv7x6;
wire Rxv7x6, Yxv7x6, Fyv7x6, Myv7x6, Tyv7x6, Azv7x6, Hzv7x6, Ozv7x6, Vzv7x6, C0w7x6;
wire J0w7x6, Q0w7x6, X0w7x6, E1w7x6, L1w7x6, S1w7x6, Z1w7x6, G2w7x6, N2w7x6, U2w7x6;
wire B3w7x6, I3w7x6, P3w7x6, W3w7x6, D4w7x6, K4w7x6, R4w7x6, Y4w7x6, F5w7x6, M5w7x6;
wire T5w7x6, A6w7x6, H6w7x6, O6w7x6, V6w7x6, C7w7x6, J7w7x6, Q7w7x6, X7w7x6, E8w7x6;
wire L8w7x6, S8w7x6, Z8w7x6, G9w7x6, N9w7x6, U9w7x6, Baw7x6, Iaw7x6, Paw7x6, Waw7x6;
wire Dbw7x6, Kbw7x6, Rbw7x6, Ybw7x6, Fcw7x6, Mcw7x6, Tcw7x6, Adw7x6, Hdw7x6, Odw7x6;
wire Vdw7x6, Cew7x6, Jew7x6, Qew7x6, Xew7x6, Efw7x6, Lfw7x6, Sfw7x6, Zfw7x6, Ggw7x6;
wire Ngw7x6, Ugw7x6, Bhw7x6, Ihw7x6, Phw7x6, Whw7x6, Diw7x6, Kiw7x6, Riw7x6, Yiw7x6;
wire Fjw7x6, Mjw7x6, Tjw7x6, Akw7x6, Hkw7x6, Okw7x6, Vkw7x6, Clw7x6, Jlw7x6, Qlw7x6;
wire Xlw7x6, Emw7x6, Lmw7x6, Smw7x6, Zmw7x6, Gnw7x6, Nnw7x6, Unw7x6, Bow7x6, Iow7x6;
wire Pow7x6, Wow7x6, Dpw7x6, Kpw7x6, Rpw7x6, Ypw7x6, Fqw7x6, Mqw7x6, Tqw7x6, Arw7x6;
wire Hrw7x6, Orw7x6, Vrw7x6, Csw7x6, Jsw7x6, Qsw7x6, Xsw7x6, Etw7x6, Ltw7x6, Stw7x6;
wire Ztw7x6, Guw7x6, Nuw7x6, Uuw7x6, Bvw7x6, Ivw7x6, Pvw7x6, Wvw7x6, Dww7x6, Kww7x6;
wire Rww7x6, Yww7x6, Fxw7x6, Mxw7x6, Txw7x6, Ayw7x6, Hyw7x6, Oyw7x6, Vyw7x6, Czw7x6;
wire Jzw7x6, Qzw7x6, Xzw7x6, E0x7x6, L0x7x6, S0x7x6, Z0x7x6, G1x7x6, N1x7x6, U1x7x6;
wire B2x7x6, I2x7x6, P2x7x6, W2x7x6, D3x7x6, K3x7x6, R3x7x6, Y3x7x6, F4x7x6, M4x7x6;
wire T4x7x6, A5x7x6, H5x7x6, O5x7x6, V5x7x6, C6x7x6, J6x7x6, Q6x7x6, X6x7x6, E7x7x6;
wire L7x7x6, S7x7x6, Z7x7x6, G8x7x6, N8x7x6, U8x7x6, B9x7x6, I9x7x6, P9x7x6, W9x7x6;
wire Dax7x6, Kax7x6, Rax7x6, Yax7x6, Fbx7x6, Mbx7x6, Tbx7x6, Acx7x6, Hcx7x6, Ocx7x6;
wire Vcx7x6, Cdx7x6, Jdx7x6, Qdx7x6, Xdx7x6, Eex7x6, Lex7x6, Sex7x6, Zex7x6, Gfx7x6;
wire Nfx7x6, Ufx7x6, Bgx7x6, Igx7x6, Pgx7x6, Wgx7x6, Dhx7x6, Khx7x6, Rhx7x6, Yhx7x6;
wire Fix7x6, Mix7x6, Tix7x6, Ajx7x6, Hjx7x6, Ojx7x6, Vjx7x6, Ckx7x6, Jkx7x6, Qkx7x6;
wire Xkx7x6, Elx7x6, Llx7x6, Slx7x6, Zlx7x6, Gmx7x6, Nmx7x6, Umx7x6, Bnx7x6, Inx7x6;
wire Pnx7x6, Wnx7x6, Dox7x6, Kox7x6, Rox7x6, Yox7x6, Fpx7x6, Mpx7x6, Tpx7x6, Aqx7x6;
wire Hqx7x6, Oqx7x6, Vqx7x6, Crx7x6, Jrx7x6, Qrx7x6, Xrx7x6, Esx7x6, Lsx7x6, Ssx7x6;
wire Zsx7x6, Gtx7x6, Ntx7x6, Utx7x6, Bux7x6, Iux7x6, Pux7x6, Wux7x6, Dvx7x6, Kvx7x6;
wire Rvx7x6, Yvx7x6, Fwx7x6, Mwx7x6, Twx7x6, Axx7x6, Hxx7x6, Oxx7x6, Vxx7x6, Cyx7x6;
wire Jyx7x6, Qyx7x6, Xyx7x6, Ezx7x6, Lzx7x6, Szx7x6, Zzx7x6, G0y7x6, N0y7x6, U0y7x6;
wire B1y7x6, I1y7x6, P1y7x6, W1y7x6, D2y7x6, K2y7x6, R2y7x6, Y2y7x6, F3y7x6, M3y7x6;
wire T3y7x6, A4y7x6, H4y7x6, O4y7x6, V4y7x6, C5y7x6, J5y7x6, Q5y7x6, X5y7x6, E6y7x6;
wire L6y7x6, S6y7x6, Z6y7x6, G7y7x6, N7y7x6, U7y7x6, B8y7x6, I8y7x6, P8y7x6, W8y7x6;
wire D9y7x6, K9y7x6, R9y7x6, Y9y7x6, Fay7x6, May7x6, Tay7x6, Aby7x6, Hby7x6, Oby7x6;
wire Vby7x6, Ccy7x6, Jcy7x6, Qcy7x6, Xcy7x6, Edy7x6, Ldy7x6, Sdy7x6, Zdy7x6, Gey7x6;
wire Ney7x6, Uey7x6, Bfy7x6, Ify7x6, Pfy7x6, Wfy7x6, Dgy7x6, Kgy7x6, Rgy7x6, Ygy7x6;
wire Fhy7x6, Mhy7x6, Thy7x6, Aiy7x6, Hiy7x6, Oiy7x6, Viy7x6, Cjy7x6, Jjy7x6, Qjy7x6;
wire Xjy7x6, Eky7x6, Lky7x6, Sky7x6, Zky7x6, Gly7x6, Nly7x6, Uly7x6, Bmy7x6, Imy7x6;
wire Pmy7x6, Wmy7x6, Dny7x6, Kny7x6, Rny7x6, Yny7x6, Foy7x6, Moy7x6, Toy7x6, Apy7x6;
wire Hpy7x6, Opy7x6, Vpy7x6, Cqy7x6, Jqy7x6, Qqy7x6, Xqy7x6, Ery7x6, Lry7x6, Sry7x6;
wire Zry7x6, Gsy7x6, Nsy7x6, Usy7x6, Bty7x6, Ity7x6, Pty7x6, Wty7x6, Duy7x6, Kuy7x6;
wire Ruy7x6, Yuy7x6, Fvy7x6, Mvy7x6, Tvy7x6, Awy7x6, Hwy7x6, Owy7x6, Vwy7x6, Cxy7x6;
wire Jxy7x6, Qxy7x6, Xxy7x6, Eyy7x6, Lyy7x6, Syy7x6, Zyy7x6, Gzy7x6, Nzy7x6, Uzy7x6;
wire B0z7x6, I0z7x6, P0z7x6, W0z7x6, D1z7x6, K1z7x6, R1z7x6, Y1z7x6, F2z7x6, M2z7x6;
wire T2z7x6, A3z7x6, H3z7x6, O3z7x6, V3z7x6, C4z7x6, J4z7x6, Q4z7x6, X4z7x6, E5z7x6;
wire L5z7x6, S5z7x6, Z5z7x6, G6z7x6, N6z7x6, U6z7x6, B7z7x6, I7z7x6, P7z7x6, W7z7x6;
wire D8z7x6, K8z7x6, R8z7x6, Y8z7x6, F9z7x6, M9z7x6, T9z7x6, Aaz7x6, Haz7x6, Oaz7x6;
wire Vaz7x6, Cbz7x6, Jbz7x6, Qbz7x6, Xbz7x6, Ecz7x6, Lcz7x6, Scz7x6, Zcz7x6, Gdz7x6;
wire Ndz7x6, Udz7x6, Bez7x6, Iez7x6, Pez7x6, Wez7x6, Dfz7x6, Kfz7x6, Rfz7x6, Yfz7x6;
wire Fgz7x6, Mgz7x6, Tgz7x6, Ahz7x6, Hhz7x6, Ohz7x6, Vhz7x6, Ciz7x6, Jiz7x6, Qiz7x6;
wire Xiz7x6, Ejz7x6, Ljz7x6, Sjz7x6, Zjz7x6, Gkz7x6, Nkz7x6, Ukz7x6, Blz7x6, Ilz7x6;
wire Plz7x6, Wlz7x6, Dmz7x6, Kmz7x6, Rmz7x6, Ymz7x6, Fnz7x6, Mnz7x6, Tnz7x6, Aoz7x6;
wire Hoz7x6, Ooz7x6, Voz7x6, Cpz7x6, Jpz7x6, Qpz7x6, Xpz7x6, Eqz7x6, Lqz7x6, Sqz7x6;
wire Zqz7x6, Grz7x6, Nrz7x6, Urz7x6, Bsz7x6, Isz7x6, Psz7x6, Wsz7x6, Dtz7x6, Ktz7x6;
wire Rtz7x6, Ytz7x6, Fuz7x6, Muz7x6, Tuz7x6, Avz7x6, Hvz7x6, Ovz7x6, Vvz7x6, Cwz7x6;
wire Jwz7x6, Qwz7x6, Xwz7x6, Exz7x6, Lxz7x6, Sxz7x6, Zxz7x6, Gyz7x6, Nyz7x6, Uyz7x6;
wire Bzz7x6, Izz7x6, Pzz7x6, Wzz7x6, D008x6, K008x6, R008x6, Y008x6, F108x6, M108x6;
wire T108x6, A208x6, H208x6, O208x6, V208x6, C308x6, J308x6, Q308x6, X308x6, E408x6;
wire L408x6, S408x6, Z408x6, G508x6, N508x6, U508x6, B608x6, I608x6, P608x6, W608x6;
wire D708x6, K708x6, R708x6, Y708x6, F808x6, M808x6, T808x6, A908x6, H908x6, O908x6;
wire V908x6, Ca08x6, Ja08x6, Qa08x6, Xa08x6, Eb08x6, Lb08x6, Sb08x6, Zb08x6, Gc08x6;
wire Nc08x6, Uc08x6, Bd08x6, Id08x6, Pd08x6, Wd08x6, De08x6, Ke08x6, Re08x6, Ye08x6;
wire Ff08x6, Mf08x6, Tf08x6, Ag08x6, Hg08x6, Og08x6, Vg08x6, Ch08x6, Jh08x6, Qh08x6;
wire Xh08x6, Ei08x6, Li08x6, Si08x6, Zi08x6, Gj08x6, Nj08x6, Uj08x6, Bk08x6, Ik08x6;
wire Pk08x6, Wk08x6, Dl08x6, Kl08x6, Rl08x6, Yl08x6, Fm08x6, Mm08x6, Tm08x6, An08x6;
wire Hn08x6, On08x6, Vn08x6, Co08x6, Jo08x6, Qo08x6, Xo08x6, Ep08x6, Lp08x6, Sp08x6;
wire Zp08x6, Gq08x6, Nq08x6, Uq08x6, Br08x6, Ir08x6, Pr08x6, Wr08x6, Ds08x6, Ks08x6;
wire Rs08x6, Ys08x6, Ft08x6, Mt08x6, Tt08x6, Au08x6, Hu08x6, Ou08x6, Vu08x6, Cv08x6;
wire Jv08x6, Qv08x6, Xv08x6, Ew08x6, Lw08x6, Sw08x6, Zw08x6, Gx08x6, Nx08x6, Ux08x6;
wire By08x6, Iy08x6, Py08x6, Wy08x6, Dz08x6, Kz08x6, Rz08x6, Yz08x6, F018x6, M018x6;
wire T018x6, A118x6, H118x6, O118x6, V118x6, C218x6, J218x6, Q218x6, X218x6, E318x6;
wire L318x6, S318x6, Z318x6, G418x6, N418x6, U418x6, B518x6, I518x6, P518x6, W518x6;
wire D618x6, K618x6, R618x6, Y618x6, F718x6, M718x6, T718x6, A818x6, H818x6, O818x6;
wire V818x6, C918x6, J918x6, Q918x6, X918x6, Ea18x6, La18x6, Sa18x6, Za18x6, Gb18x6;
wire Nb18x6, Ub18x6, Bc18x6, Ic18x6, Pc18x6, Wc18x6, Dd18x6, Kd18x6, Rd18x6, Yd18x6;
wire Fe18x6, Me18x6, Te18x6, Af18x6, Hf18x6, Of18x6, Vf18x6, Cg18x6, Jg18x6, Qg18x6;
wire Xg18x6, Eh18x6, Lh18x6, Sh18x6, Zh18x6, Gi18x6, Ni18x6, Ui18x6, Bj18x6, Ij18x6;
wire Pj18x6, Wj18x6, Dk18x6, Kk18x6, Rk18x6, Yk18x6, Fl18x6, Ml18x6, Tl18x6, Am18x6;
wire Hm18x6, Om18x6, Vm18x6, Cn18x6, Jn18x6, Qn18x6, Xn18x6, Eo18x6, Lo18x6, So18x6;
wire Zo18x6, Gp18x6, Np18x6, Up18x6, Bq18x6, Iq18x6, Pq18x6, Wq18x6, Dr18x6, Kr18x6;
wire Rr18x6, Yr18x6, Fs18x6, Ms18x6, Ts18x6, At18x6, Ht18x6, Ot18x6, Vt18x6, Cu18x6;
wire Ju18x6, Qu18x6, Xu18x6, Ev18x6, Lv18x6, Sv18x6, Zv18x6, Gw18x6, Nw18x6, Uw18x6;
wire Bx18x6, Ix18x6, Px18x6, Wx18x6, Dy18x6, Ky18x6, Ry18x6, Yy18x6, Fz18x6, Mz18x6;
wire Tz18x6, A028x6, H028x6, O028x6, V028x6, C128x6, J128x6, Q128x6, X128x6, E228x6;
wire L228x6, S228x6, Z228x6, G328x6, N328x6, U328x6, B428x6, I428x6, P428x6, W428x6;
wire D528x6, K528x6, R528x6, Y528x6, F628x6, M628x6, T628x6, A728x6, H728x6, O728x6;
wire V728x6, C828x6, J828x6, Q828x6, X828x6, E928x6, L928x6, S928x6, Z928x6, Ga28x6;
wire Na28x6, Ua28x6, Bb28x6, Ib28x6, Pb28x6, Wb28x6, Dc28x6, Kc28x6, Rc28x6, Yc28x6;
wire Fd28x6, Md28x6, Td28x6, Ae28x6, He28x6, Oe28x6, Ve28x6, Cf28x6, Jf28x6, Qf28x6;
wire Xf28x6, Eg28x6, Lg28x6, Sg28x6, Zg28x6, Gh28x6, Nh28x6, Uh28x6, Bi28x6, Ii28x6;
wire Pi28x6, Wi28x6, Dj28x6, Kj28x6, Rj28x6, Yj28x6, Fk28x6, Mk28x6, Tk28x6, Al28x6;
wire Hl28x6, Ol28x6, Vl28x6, Cm28x6, Jm28x6, Qm28x6, Xm28x6, En28x6, Ln28x6, Sn28x6;
wire Zn28x6, Go28x6, No28x6, Uo28x6, Bp28x6, Ip28x6, Pp28x6, Wp28x6, Dq28x6, Kq28x6;
wire Rq28x6, Yq28x6, Fr28x6, Mr28x6, Tr28x6, As28x6, Hs28x6, Os28x6, Vs28x6, Ct28x6;
wire Jt28x6, Qt28x6, Xt28x6, Eu28x6, Lu28x6, Su28x6, Zu28x6, Gv28x6, Nv28x6, Uv28x6;
wire Bw28x6, Iw28x6, Pw28x6, Ww28x6, Dx28x6, Kx28x6, Rx28x6, Yx28x6, Fy28x6, My28x6;
wire Ty28x6, Az28x6, Hz28x6, Oz28x6, Vz28x6, C038x6, J038x6, Q038x6, X038x6, E138x6;
wire L138x6, S138x6, Z138x6, G238x6, N238x6, U238x6, B338x6, I338x6, P338x6, W338x6;
wire D438x6, K438x6, R438x6, Y438x6, F538x6, M538x6, T538x6, A638x6, H638x6, O638x6;
wire V638x6, C738x6, J738x6, Q738x6, X738x6, E838x6, L838x6, S838x6, Z838x6, G938x6;
wire N938x6, U938x6, Ba38x6, Ia38x6, Pa38x6, Wa38x6, Db38x6, Kb38x6, Rb38x6, Yb38x6;
wire Fc38x6, Mc38x6, Tc38x6, Ad38x6, Hd38x6, Od38x6, Vd38x6, Ce38x6, Je38x6, Qe38x6;
wire Xe38x6, Ef38x6, Lf38x6, Sf38x6, Zf38x6, Gg38x6, Ng38x6, Ug38x6, Bh38x6, Ih38x6;
wire Ph38x6, Wh38x6, Di38x6, Ki38x6, Ri38x6, Yi38x6, Fj38x6, Mj38x6, Tj38x6, Ak38x6;
wire Hk38x6, Ok38x6, Vk38x6, Cl38x6, Jl38x6, Ql38x6, Xl38x6, Em38x6, Lm38x6, Sm38x6;
wire Zm38x6, Gn38x6, Nn38x6, Un38x6, Bo38x6, Io38x6, Po38x6, Wo38x6, Dp38x6, Kp38x6;
wire Rp38x6, Yp38x6, Fq38x6, Mq38x6, Tq38x6, Ar38x6, Hr38x6, Or38x6, Vr38x6, Cs38x6;
wire Js38x6, Qs38x6, Xs38x6, Et38x6, Lt38x6, St38x6, Zt38x6, Gu38x6, Nu38x6, Uu38x6;
wire Bv38x6, Iv38x6, Pv38x6, Wv38x6, Dw38x6, Kw38x6, Rw38x6, Yw38x6, Fx38x6, Mx38x6;
wire Tx38x6, Ay38x6, Hy38x6, Oy38x6, Vy38x6, Cz38x6, Jz38x6, Qz38x6, Xz38x6, E048x6;
wire L048x6, S048x6, Z048x6, G148x6, N148x6, U148x6, B248x6, I248x6, P248x6, W248x6;
wire D348x6, K348x6, R348x6, Y348x6, F448x6, M448x6, T448x6, A548x6, H548x6, O548x6;
wire V548x6, C648x6, J648x6, Q648x6, X648x6, E748x6, L748x6, S748x6, Z748x6, G848x6;
wire N848x6, U848x6, B948x6, I948x6, P948x6, W948x6, Da48x6, Ka48x6, Ra48x6, Ya48x6;
wire Fb48x6, Mb48x6, Tb48x6, Ac48x6, Hc48x6, Oc48x6, Vc48x6, Cd48x6, Jd48x6, Qd48x6;
wire Xd48x6, Ee48x6, Le48x6, Se48x6, Ze48x6, Gf48x6, Nf48x6, Uf48x6, Bg48x6, Ig48x6;
wire Pg48x6, Wg48x6, Dh48x6, Kh48x6, Rh48x6, Yh48x6, Fi48x6, Mi48x6, Ti48x6, Aj48x6;
wire Hj48x6, Oj48x6, Vj48x6, Ck48x6, Jk48x6, Qk48x6, Xk48x6, El48x6, Ll48x6, Sl48x6;
wire Zl48x6, Gm48x6, Nm48x6, Um48x6, Bn48x6, In48x6, Pn48x6, Wn48x6, Do48x6, Ko48x6;
wire Ro48x6, Yo48x6, Fp48x6, Mp48x6, Tp48x6, Aq48x6, Hq48x6, Oq48x6, Vq48x6, Cr48x6;
wire Jr48x6, Qr48x6, Xr48x6, Es48x6, Ls48x6, Ss48x6, Zs48x6, Gt48x6, Nt48x6, Ut48x6;
wire Bu48x6, Iu48x6, Pu48x6, Wu48x6, Dv48x6, Kv48x6, Rv48x6, Yv48x6, Fw48x6, Mw48x6;
wire Tw48x6, Ax48x6, Hx48x6, Ox48x6, Vx48x6, Cy48x6, Jy48x6, Qy48x6, Xy48x6, Ez48x6;
wire Lz48x6, Sz48x6, Zz48x6, G058x6, N058x6, U058x6, B158x6, I158x6, P158x6, W158x6;
wire D258x6, K258x6, R258x6, Y258x6, F358x6, M358x6, T358x6, A458x6, H458x6, O458x6;
wire V458x6, C558x6, J558x6, Q558x6, X558x6, E658x6, L658x6, S658x6, Z658x6, G758x6;
wire N758x6, U758x6, B858x6, I858x6, P858x6, W858x6, D958x6, K958x6, R958x6, Y958x6;
wire Fa58x6, Ma58x6, Ta58x6, Ab58x6, Hb58x6, Ob58x6, Vb58x6, Cc58x6, Jc58x6, Qc58x6;
wire Xc58x6, Ed58x6, Ld58x6, Sd58x6, Zd58x6, Ge58x6, Ne58x6, Ue58x6, Bf58x6, If58x6;
wire Pf58x6, Wf58x6, Dg58x6, Kg58x6, Rg58x6, Yg58x6, Fh58x6, Mh58x6, Th58x6, Ai58x6;
wire Hi58x6, Oi58x6, Vi58x6, Cj58x6, Jj58x6, Qj58x6, Xj58x6, Ek58x6, Lk58x6, Sk58x6;
wire Zk58x6, Gl58x6, Nl58x6, Ul58x6, Bm58x6, Im58x6, Pm58x6, Wm58x6, Dn58x6, Kn58x6;
wire Rn58x6, Yn58x6, Fo58x6, Mo58x6, To58x6, Ap58x6, Hp58x6, Op58x6, Vp58x6, Cq58x6;
wire Jq58x6, Qq58x6, Xq58x6, Er58x6, Lr58x6, Sr58x6, Zr58x6, Gs58x6, Ns58x6, Us58x6;
wire Bt58x6, It58x6, Pt58x6, Wt58x6, Du58x6, Ku58x6, Ru58x6, Yu58x6, Fv58x6, Mv58x6;
wire Tv58x6, Aw58x6, Hw58x6, Ow58x6, Vw58x6, Cx58x6, Jx58x6, Qx58x6, Xx58x6, Ey58x6;
wire Ly58x6, Sy58x6, Zy58x6, Gz58x6, Nz58x6, Uz58x6, B068x6, I068x6, P068x6, W068x6;
wire D168x6, K168x6, R168x6, Y168x6, F268x6, M268x6, T268x6, A368x6, H368x6, O368x6;
wire V368x6, C468x6, J468x6, Q468x6, X468x6, E568x6, L568x6, S568x6, Z568x6, G668x6;
wire N668x6, U668x6, B768x6, I768x6, P768x6, W768x6, D868x6, K868x6, R868x6, Y868x6;
wire F968x6, M968x6, T968x6, Aa68x6, Ha68x6, Oa68x6, Va68x6, Cb68x6, Jb68x6, Qb68x6;
wire Xb68x6, Ec68x6, Lc68x6, Sc68x6, Zc68x6, Gd68x6, Nd68x6, Ud68x6, Be68x6, Ie68x6;
wire Pe68x6, We68x6, Df68x6, Kf68x6, Rf68x6, Yf68x6, Fg68x6, Mg68x6, Tg68x6, Ah68x6;
wire Hh68x6, Oh68x6, Vh68x6, Ci68x6, Ji68x6, Qi68x6, Xi68x6, Ej68x6, Lj68x6, Sj68x6;
wire Zj68x6, Gk68x6, Nk68x6, Uk68x6, Bl68x6, Il68x6, Pl68x6, Wl68x6, Dm68x6, Km68x6;
wire Rm68x6, Ym68x6, Fn68x6, Mn68x6, Tn68x6, Ao68x6, Ho68x6, Oo68x6, Vo68x6, Cp68x6;
wire Jp68x6, Qp68x6, Xp68x6, Eq68x6, Lq68x6, Sq68x6, Zq68x6, Gr68x6, Nr68x6, Ur68x6;
wire Bs68x6, Is68x6, Ps68x6, Ws68x6, Dt68x6, Kt68x6, Rt68x6, Yt68x6, Fu68x6, Mu68x6;
wire Tu68x6, Av68x6, Hv68x6, Ov68x6, Vv68x6, Cw68x6, Jw68x6, Qw68x6, Xw68x6, Ex68x6;
wire Lx68x6, Sx68x6, Zx68x6, Gy68x6, Ny68x6, Uy68x6, Bz68x6, Iz68x6, Pz68x6, Wz68x6;
wire D078x6, K078x6, R078x6, Y078x6, F178x6, M178x6, T178x6, A278x6, H278x6, O278x6;
wire V278x6, C378x6, J378x6, Q378x6, X378x6, E478x6, L478x6, S478x6, Z478x6, G578x6;
wire N578x6, U578x6, B678x6, I678x6, P678x6, W678x6, D778x6, K778x6, R778x6, Y778x6;
wire F878x6, M878x6, T878x6, A978x6, H978x6, O978x6, V978x6, Ca78x6, Ja78x6, Qa78x6;
wire Xa78x6, Eb78x6, Lb78x6, Sb78x6, Zb78x6, Gc78x6, Nc78x6, Uc78x6, Bd78x6, Id78x6;
wire Pd78x6, Wd78x6, De78x6, Ke78x6, Re78x6, Ye78x6, Ff78x6, Mf78x6, Tf78x6, Ag78x6;
wire Hg78x6, Og78x6, Vg78x6, Ch78x6, Jh78x6, Qh78x6, Xh78x6, Ei78x6, Li78x6, Si78x6;
wire Zi78x6, Gj78x6, Nj78x6, Uj78x6, Bk78x6, Ik78x6, Pk78x6, Wk78x6, Dl78x6, Kl78x6;
wire Rl78x6, Yl78x6, Fm78x6, Mm78x6, Tm78x6, An78x6, Hn78x6, On78x6, Vn78x6, Co78x6;
wire Jo78x6, Qo78x6, Xo78x6, Ep78x6, Lp78x6, Sp78x6, Zp78x6, Gq78x6, Nq78x6, Uq78x6;
wire Br78x6, Ir78x6, Pr78x6, Wr78x6, Ds78x6, Ks78x6, Rs78x6, Ys78x6, Ft78x6, Mt78x6;
wire Tt78x6, Au78x6, Hu78x6, Ou78x6, Vu78x6, Cv78x6, Jv78x6, Qv78x6, Xv78x6, Ew78x6;
wire Lw78x6, Sw78x6, Zw78x6, Gx78x6, Nx78x6, Ux78x6, By78x6, Iy78x6, Py78x6, Wy78x6;
wire Dz78x6, Kz78x6, Rz78x6, Yz78x6, F088x6, M088x6, T088x6, A188x6, H188x6, O188x6;
wire V188x6, C288x6, J288x6, Q288x6, X288x6, E388x6, L388x6, S388x6, Z388x6, G488x6;
wire N488x6, U488x6, B588x6, I588x6, P588x6, W588x6, D688x6, K688x6, R688x6, Y688x6;
wire F788x6, M788x6, T788x6, A888x6, H888x6, O888x6, V888x6, C988x6, J988x6, Q988x6;
wire X988x6, Ea88x6, La88x6, Sa88x6, Za88x6, Gb88x6, Nb88x6, Ub88x6, Bc88x6, Ic88x6;
wire Pc88x6, Wc88x6, Dd88x6, Kd88x6, Rd88x6, Yd88x6, Fe88x6, Me88x6, Te88x6, Af88x6;
wire Hf88x6, Of88x6, Vf88x6, Cg88x6, Jg88x6, Qg88x6, Xg88x6, Eh88x6, Lh88x6, Sh88x6;
wire Zh88x6, Gi88x6, Ni88x6, Ui88x6, Bj88x6, Ij88x6, Pj88x6, Wj88x6, Dk88x6, Kk88x6;
wire Rk88x6, Yk88x6, Fl88x6, Ml88x6, Tl88x6, Am88x6, Hm88x6, Om88x6, Vm88x6, Cn88x6;
wire Jn88x6, Qn88x6, Xn88x6, Eo88x6, Lo88x6, So88x6, Zo88x6, Gp88x6, Np88x6, Up88x6;
wire Bq88x6, Iq88x6, Pq88x6, Wq88x6, Dr88x6, Kr88x6, Rr88x6, Yr88x6, Fs88x6, Ms88x6;
wire Ts88x6, At88x6, Ht88x6, Ot88x6, Vt88x6, Cu88x6, Ju88x6, Qu88x6, Xu88x6, Ev88x6;
wire Lv88x6, Sv88x6, Zv88x6, Gw88x6, Nw88x6, Uw88x6, Bx88x6, Ix88x6, Px88x6, Wx88x6;
wire Dy88x6, Ky88x6, Ry88x6, Yy88x6, Fz88x6, Mz88x6, Tz88x6, A098x6, H098x6, O098x6;
wire V098x6, C198x6, J198x6, Q198x6, X198x6, E298x6, L298x6, S298x6, Z298x6, G398x6;
wire N398x6, U398x6, B498x6, I498x6, P498x6, W498x6, D598x6, K598x6, R598x6, Y598x6;
wire F698x6, M698x6, T698x6, A798x6, H798x6, O798x6, V798x6, C898x6, J898x6, Q898x6;
wire X898x6, E998x6, L998x6, S998x6, Z998x6, Ga98x6, Na98x6, Ua98x6, Bb98x6, Ib98x6;
wire Pb98x6, Wb98x6, Dc98x6, Kc98x6, Rc98x6, Yc98x6, Fd98x6, Md98x6, Td98x6, Ae98x6;
wire He98x6, Oe98x6, Ve98x6, Cf98x6, Jf98x6, Qf98x6, Xf98x6, Eg98x6, Lg98x6, Sg98x6;
wire Zg98x6, Gh98x6, Nh98x6, Uh98x6, Bi98x6, Ii98x6, Pi98x6, Wi98x6, Dj98x6, Kj98x6;
wire Rj98x6, Yj98x6, Fk98x6, Mk98x6, Tk98x6, Al98x6, Hl98x6, Ol98x6, Vl98x6, Cm98x6;
wire Jm98x6, Qm98x6, Xm98x6, En98x6, Ln98x6, Sn98x6, Zn98x6, Go98x6, No98x6, Uo98x6;
wire Bp98x6, Ip98x6, Pp98x6, Wp98x6, Dq98x6, Kq98x6, Rq98x6, Yq98x6, Fr98x6, Mr98x6;
wire Tr98x6, As98x6, Hs98x6, Os98x6, Vs98x6, Ct98x6, Jt98x6, Qt98x6, Xt98x6, Eu98x6;
wire Lu98x6, Su98x6, Zu98x6, Gv98x6, Nv98x6, Uv98x6, Bw98x6, Iw98x6, Pw98x6, Ww98x6;
wire Dx98x6, Kx98x6, Rx98x6, Yx98x6, Fy98x6, My98x6, Ty98x6, Az98x6, Hz98x6, Oz98x6;
wire Vz98x6, C0a8x6, J0a8x6, Q0a8x6, X0a8x6, E1a8x6, L1a8x6, S1a8x6, Z1a8x6, G2a8x6;
wire N2a8x6, U2a8x6, B3a8x6, I3a8x6, P3a8x6, W3a8x6, D4a8x6, K4a8x6, R4a8x6, Y4a8x6;
wire F5a8x6, M5a8x6, T5a8x6, A6a8x6, H6a8x6, O6a8x6, V6a8x6, C7a8x6, J7a8x6, Q7a8x6;
wire X7a8x6, E8a8x6, L8a8x6, S8a8x6, Z8a8x6, G9a8x6, N9a8x6, U9a8x6, Baa8x6, Iaa8x6;
wire Paa8x6, Waa8x6, Dba8x6, Kba8x6, Rba8x6, Yba8x6, Fca8x6, Mca8x6, Tca8x6, Ada8x6;
wire Hda8x6, Oda8x6, Vda8x6, Cea8x6, Jea8x6, Qea8x6, Xea8x6, Efa8x6, Lfa8x6, Sfa8x6;
wire Zfa8x6, Gga8x6, Nga8x6, Uga8x6, Bha8x6, Iha8x6, Pha8x6, Wha8x6, Dia8x6, Kia8x6;
wire Ria8x6, Yia8x6, Fja8x6, Mja8x6, Tja8x6, Aka8x6, Hka8x6, Oka8x6, Vka8x6, Cla8x6;
wire Jla8x6, Qla8x6, Xla8x6, Ema8x6, Lma8x6, Sma8x6, Zma8x6, Gna8x6, Nna8x6, Una8x6;
wire Boa8x6, Ioa8x6, Poa8x6, Woa8x6, Dpa8x6, Kpa8x6, Rpa8x6, Ypa8x6, Fqa8x6, Mqa8x6;
wire Tqa8x6, Ara8x6, Hra8x6, Ora8x6, Vra8x6, Csa8x6, Jsa8x6, Qsa8x6, Xsa8x6, Eta8x6;
wire Lta8x6, Sta8x6, Zta8x6, Gua8x6, Nua8x6, Uua8x6, Bva8x6, Iva8x6, Pva8x6, Wva8x6;
wire Dwa8x6, Kwa8x6, Rwa8x6, Ywa8x6, Fxa8x6, Mxa8x6, Txa8x6, Aya8x6, Hya8x6, Oya8x6;
wire Vya8x6, Cza8x6, Jza8x6, Qza8x6, Xza8x6, E0b8x6, L0b8x6, S0b8x6, Z0b8x6, G1b8x6;
wire N1b8x6, U1b8x6, B2b8x6, I2b8x6, P2b8x6, W2b8x6, D3b8x6, K3b8x6, R3b8x6, Y3b8x6;
wire F4b8x6, M4b8x6, T4b8x6, A5b8x6, H5b8x6, O5b8x6, V5b8x6, C6b8x6, J6b8x6, Q6b8x6;
wire X6b8x6, E7b8x6, L7b8x6, S7b8x6, Z7b8x6, G8b8x6, N8b8x6, U8b8x6, B9b8x6, I9b8x6;
wire P9b8x6, W9b8x6, Dab8x6, Kab8x6, Rab8x6, Yab8x6, Fbb8x6, Mbb8x6, Tbb8x6, Acb8x6;
wire Hcb8x6, Ocb8x6, Vcb8x6, Cdb8x6, Jdb8x6, Qdb8x6, Xdb8x6, Eeb8x6, Leb8x6, Seb8x6;
wire Zeb8x6, Gfb8x6, Nfb8x6, Ufb8x6, Bgb8x6, Igb8x6, Pgb8x6, Wgb8x6, Dhb8x6, Khb8x6;
wire Rhb8x6, Yhb8x6, Fib8x6, Mib8x6, Tib8x6, Ajb8x6, Hjb8x6, Ojb8x6, Vjb8x6, Ckb8x6;
wire Jkb8x6, Qkb8x6, Xkb8x6, Elb8x6, Llb8x6, Slb8x6, Zlb8x6, Gmb8x6, Nmb8x6, Umb8x6;
wire Bnb8x6, Inb8x6, Pnb8x6, Wnb8x6, Dob8x6, Kob8x6, Rob8x6, Yob8x6, Fpb8x6, Mpb8x6;
wire Tpb8x6, Aqb8x6, Hqb8x6, Oqb8x6, Vqb8x6, Crb8x6, Jrb8x6, Qrb8x6, Xrb8x6, Esb8x6;
wire Lsb8x6, Ssb8x6, Zsb8x6, Gtb8x6, Ntb8x6, Utb8x6, Bub8x6, Iub8x6, Pub8x6, Wub8x6;
wire Dvb8x6, Kvb8x6, Rvb8x6, Yvb8x6, Fwb8x6, Mwb8x6, Twb8x6, Axb8x6, Hxb8x6, Oxb8x6;
wire Vxb8x6, Cyb8x6, Jyb8x6, Qyb8x6, Xyb8x6, Ezb8x6, Lzb8x6, Szb8x6, Zzb8x6, G0c8x6;
wire N0c8x6, U0c8x6, B1c8x6, I1c8x6, P1c8x6, W1c8x6, D2c8x6, K2c8x6, R2c8x6, Y2c8x6;
wire F3c8x6, M3c8x6, T3c8x6, A4c8x6, H4c8x6, O4c8x6, V4c8x6, C5c8x6, J5c8x6, Q5c8x6;
wire X5c8x6, E6c8x6, L6c8x6, S6c8x6, Z6c8x6, G7c8x6, N7c8x6, U7c8x6, B8c8x6, I8c8x6;
wire P8c8x6, W8c8x6, D9c8x6, K9c8x6, R9c8x6, Y9c8x6, Fac8x6, Mac8x6, Tac8x6, Abc8x6;
wire Hbc8x6, Obc8x6, Vbc8x6, Ccc8x6, Jcc8x6, Qcc8x6, Xcc8x6, Edc8x6, Ldc8x6, Sdc8x6;
wire Zdc8x6, Gec8x6, Nec8x6, Uec8x6, Bfc8x6, Ifc8x6, Pfc8x6, Wfc8x6, Dgc8x6, Kgc8x6;
wire Rgc8x6, Ygc8x6, Fhc8x6, Mhc8x6, Thc8x6, Aic8x6, Hic8x6, Oic8x6, Vic8x6, Cjc8x6;
wire Jjc8x6, Qjc8x6, Xjc8x6, Ekc8x6, Lkc8x6, Skc8x6, Zkc8x6, Glc8x6, Nlc8x6, Ulc8x6;
wire Bmc8x6, Imc8x6, Pmc8x6, Wmc8x6, Dnc8x6, Knc8x6, Rnc8x6, Ync8x6, Foc8x6, Moc8x6;
wire Toc8x6, Apc8x6, Hpc8x6, Opc8x6, Vpc8x6, Cqc8x6, Jqc8x6, Qqc8x6, Xqc8x6, Erc8x6;
wire Lrc8x6, Src8x6, Zrc8x6, Gsc8x6, Nsc8x6, Usc8x6, Btc8x6, Itc8x6, Ptc8x6, Wtc8x6;
wire Duc8x6, Kuc8x6, Ruc8x6, Yuc8x6, Fvc8x6, Mvc8x6, Tvc8x6, Awc8x6, Hwc8x6, Owc8x6;
wire Vwc8x6, Cxc8x6, Jxc8x6, Qxc8x6, Xxc8x6, Eyc8x6, Lyc8x6, Syc8x6, Zyc8x6, Gzc8x6;
wire Nzc8x6, Uzc8x6, B0d8x6, I0d8x6, P0d8x6, W0d8x6, D1d8x6, K1d8x6, R1d8x6, Y1d8x6;
wire F2d8x6, M2d8x6, T2d8x6, A3d8x6, H3d8x6, O3d8x6, V3d8x6, C4d8x6, J4d8x6, Q4d8x6;
wire X4d8x6, E5d8x6, L5d8x6, S5d8x6, Z5d8x6, G6d8x6, N6d8x6, U6d8x6, B7d8x6, I7d8x6;
wire P7d8x6, W7d8x6, D8d8x6, K8d8x6, R8d8x6, Y8d8x6, F9d8x6, M9d8x6, T9d8x6, Aad8x6;
wire Had8x6, Oad8x6, Vad8x6, Cbd8x6, Jbd8x6, Qbd8x6, Xbd8x6, Ecd8x6, Lcd8x6, Scd8x6;
wire Zcd8x6, Gdd8x6, Ndd8x6, Udd8x6, Bed8x6, Ied8x6, Ped8x6, Wed8x6, Dfd8x6, Kfd8x6;
wire Rfd8x6, Yfd8x6, Fgd8x6, Mgd8x6, Tgd8x6, Ahd8x6, Hhd8x6, Ohd8x6, Vhd8x6, Cid8x6;
wire Jid8x6, Qid8x6, Xid8x6, Ejd8x6, Ljd8x6, Sjd8x6, Zjd8x6, Gkd8x6, Nkd8x6, Ukd8x6;
wire Bld8x6, Ild8x6, Pld8x6, Wld8x6, Dmd8x6, Kmd8x6, Rmd8x6, Ymd8x6, Fnd8x6, Mnd8x6;
wire Tnd8x6, Aod8x6, Hod8x6, Ood8x6, Vod8x6, Cpd8x6, Jpd8x6, Qpd8x6, Xpd8x6, Eqd8x6;
wire Lqd8x6, Sqd8x6, Zqd8x6, Grd8x6, Nrd8x6, Urd8x6, Bsd8x6, Isd8x6, Psd8x6, Wsd8x6;
wire Dtd8x6, Ktd8x6, Rtd8x6, Ytd8x6, Fud8x6, Mud8x6, Tud8x6, Avd8x6, Hvd8x6, Ovd8x6;
wire Vvd8x6, Cwd8x6, Jwd8x6, Qwd8x6, Xwd8x6, Exd8x6, Lxd8x6, Sxd8x6, Zxd8x6, Gyd8x6;
wire Nyd8x6, Uyd8x6, Bzd8x6, Izd8x6, Pzd8x6, Wzd8x6, D0e8x6, K0e8x6, R0e8x6, Y0e8x6;
wire F1e8x6, M1e8x6, T1e8x6, A2e8x6, H2e8x6, O2e8x6, V2e8x6, C3e8x6, J3e8x6, Q3e8x6;
wire X3e8x6, E4e8x6, L4e8x6, S4e8x6, Z4e8x6, G5e8x6, N5e8x6, U5e8x6, B6e8x6, I6e8x6;
wire P6e8x6, W6e8x6, D7e8x6, K7e8x6, R7e8x6, Y7e8x6, F8e8x6, M8e8x6, T8e8x6, A9e8x6;
wire H9e8x6, O9e8x6, V9e8x6, Cae8x6, Jae8x6, Qae8x6, Xae8x6, Ebe8x6, Lbe8x6, Sbe8x6;
wire Zbe8x6, Gce8x6, Nce8x6, Uce8x6, Bde8x6, Ide8x6, Pde8x6, Wde8x6, Dee8x6, Kee8x6;
wire Ree8x6, Yee8x6, Ffe8x6, Mfe8x6, Tfe8x6, Age8x6, Hge8x6, Oge8x6, Vge8x6, Che8x6;
wire Jhe8x6, Qhe8x6, Xhe8x6, Eie8x6, Lie8x6, Sie8x6, Zie8x6, Gje8x6, Nje8x6, Uje8x6;
wire Bke8x6, Ike8x6, Pke8x6, Qg3xx6, Xg3xx6, Eh3xx6, Lh3xx6, Sh3xx6, Zh3xx6, Gi3xx6;
wire Ni3xx6, Ui3xx6, Bj3xx6, Ij3xx6, Pj3xx6, Wj3xx6, Dk3xx6, Kk3xx6, Rk3xx6, Yk3xx6;
wire Fl3xx6, Ml3xx6, Tl3xx6, Am3xx6, Hm3xx6, Om3xx6, Vm3xx6, Cn3xx6, Jn3xx6, Qn3xx6;
wire Xn3xx6, Eo3xx6, Lo3xx6, So3xx6, Zo3xx6, Gp3xx6, Np3xx6, Up3xx6, Bq3xx6, Iq3xx6;
wire Pq3xx6, Wq3xx6, Dr3xx6, Kr3xx6, Rr3xx6, Yr3xx6, Fs3xx6, Ms3xx6, Ts3xx6, At3xx6;
wire Ht3xx6, Ot3xx6, Vt3xx6, Cu3xx6, Ju3xx6, Qu3xx6, Xu3xx6, Ev3xx6, Lv3xx6, Sv3xx6;
wire Zv3xx6, Gw3xx6, Nw3xx6, Uw3xx6, Bx3xx6, Ix3xx6, Px3xx6, Wx3xx6, Dy3xx6, Ky3xx6;
wire Ry3xx6, Yy3xx6, Fz3xx6, Mz3xx6, Tz3xx6, A04xx6, H04xx6, O04xx6, V04xx6, C14xx6;
wire J14xx6, Q14xx6, X14xx6, E24xx6, L24xx6, S24xx6, Z24xx6, G34xx6, N34xx6, U34xx6;
wire B44xx6, I44xx6, P44xx6, W44xx6, D54xx6, K54xx6, R54xx6, Y54xx6, F64xx6, M64xx6;
wire T64xx6, A74xx6, H74xx6, O74xx6, V74xx6, C84xx6, J84xx6, Q84xx6, X84xx6, E94xx6;
wire L94xx6, S94xx6, Z94xx6, Ga4xx6, Na4xx6, Ua4xx6, Bb4xx6, Ib4xx6, Pb4xx6, Wb4xx6;
wire Dc4xx6, Kc4xx6, Rc4xx6, Yc4xx6, Fd4xx6, Md4xx6, Td4xx6, Ae4xx6, He4xx6, Oe4xx6;
wire Ve4xx6, Cf4xx6, Jf4xx6, Qf4xx6, Xf4xx6, Eg4xx6, Lg4xx6, Sg4xx6, Zg4xx6, Gh4xx6;
wire Nh4xx6, Uh4xx6, Bi4xx6, Ii4xx6, Pi4xx6, Wi4xx6, Dj4xx6, Kj4xx6, Rj4xx6, Yj4xx6;
wire Fk4xx6, Mk4xx6, Tk4xx6, Al4xx6, Hl4xx6, Ol4xx6, Vl4xx6, Cm4xx6, Jm4xx6, Qm4xx6;
wire Xm4xx6, En4xx6, Ln4xx6, Sn4xx6, Zn4xx6, Go4xx6, No4xx6, Uo4xx6, Bp4xx6, Ip4xx6;
wire Pp4xx6, Wp4xx6, Dq4xx6, Kq4xx6, Rq4xx6, Yq4xx6, Fr4xx6, Mr4xx6, Tr4xx6, As4xx6;
wire Hs4xx6, Os4xx6, Vs4xx6, Ct4xx6, Jt4xx6, Qt4xx6, Xt4xx6, Eu4xx6, Lu4xx6, Su4xx6;
wire Zu4xx6, Gv4xx6, Nv4xx6, Uv4xx6, Bw4xx6, Iw4xx6, Pw4xx6, Ww4xx6, Dx4xx6, Kx4xx6;
wire Rx4xx6, Yx4xx6, Fy4xx6, My4xx6, Ty4xx6, Az4xx6, Hz4xx6, Oz4xx6, Vz4xx6, C05xx6;
wire J05xx6, Q05xx6, X05xx6, E15xx6, L15xx6, S15xx6, Z15xx6, G25xx6, N25xx6, U25xx6;
wire B35xx6, I35xx6, P35xx6, W35xx6, D45xx6, K45xx6, R45xx6, Y45xx6, F55xx6, M55xx6;
wire T55xx6, A65xx6, H65xx6, O65xx6, V65xx6, C75xx6, J75xx6, Q75xx6, X75xx6, E85xx6;
wire L85xx6, S85xx6, Z85xx6, G95xx6, N95xx6, U95xx6, Ba5xx6, Ia5xx6, Pa5xx6, Wa5xx6;
wire Db5xx6, Kb5xx6, Rb5xx6, Yb5xx6, Fc5xx6, Mc5xx6, Tc5xx6, Ad5xx6, Hd5xx6, Od5xx6;
wire Vd5xx6, Ce5xx6, Je5xx6, Qe5xx6, Xe5xx6, Ef5xx6, Lf5xx6, Sf5xx6, Zf5xx6, Gg5xx6;
wire Ng5xx6, Ug5xx6, Bh5xx6, Ih5xx6, Ph5xx6, Wh5xx6, Di5xx6, Ki5xx6, Ri5xx6, Yi5xx6;
wire Fj5xx6, Mj5xx6, Tj5xx6, Ak5xx6, Hk5xx6, Ok5xx6, Vk5xx6, Cl5xx6, Jl5xx6, Ql5xx6;
wire Xl5xx6, Em5xx6, Lm5xx6, Sm5xx6, Zm5xx6, Gn5xx6, Nn5xx6, Un5xx6, Bo5xx6, Io5xx6;
wire Po5xx6, Wo5xx6, Dp5xx6, Kp5xx6, Rp5xx6, Yp5xx6, Fq5xx6, Mq5xx6, Tq5xx6, Ar5xx6;
wire Hr5xx6, Or5xx6, Vr5xx6, Cs5xx6, Js5xx6, Qs5xx6, Xs5xx6, Et5xx6, Lt5xx6, St5xx6;
wire Zt5xx6, Gu5xx6, Nu5xx6, Uu5xx6, Bv5xx6, Iv5xx6, Pv5xx6, Wv5xx6, Dw5xx6, Kw5xx6;
wire Rw5xx6, Yw5xx6, Fx5xx6, Mx5xx6, Tx5xx6, Ay5xx6, Hy5xx6, Oy5xx6, Vy5xx6, Cz5xx6;
wire Jz5xx6, Qz5xx6, Xz5xx6, E06xx6, L06xx6, S06xx6, Z06xx6, G16xx6, N16xx6, U16xx6;
wire B26xx6, I26xx6, P26xx6, W26xx6, D36xx6, K36xx6, R36xx6, Y36xx6, F46xx6, M46xx6;
wire T46xx6, A56xx6, H56xx6, O56xx6, V56xx6, C66xx6, J66xx6, Q66xx6, X66xx6, E76xx6;
wire L76xx6, S76xx6, Z76xx6, G86xx6, N86xx6, U86xx6, B96xx6, I96xx6, P96xx6, W96xx6;
wire Da6xx6, Ka6xx6, Ra6xx6, Ya6xx6, Fb6xx6, Mb6xx6, Tb6xx6, Ac6xx6, Hc6xx6, Oc6xx6;
wire Vc6xx6, Cd6xx6, Jd6xx6, Qd6xx6, Xd6xx6, Ee6xx6, Le6xx6, Se6xx6, Ze6xx6, Gf6xx6;
wire Nf6xx6, Uf6xx6, Bg6xx6, Ig6xx6, Pg6xx6, Wg6xx6, Dh6xx6, Kh6xx6, Rh6xx6, Yh6xx6;
wire Fi6xx6, Mi6xx6, Ti6xx6, Aj6xx6, Hj6xx6, Oj6xx6, Vj6xx6, Ck6xx6, Jk6xx6, Qk6xx6;
wire Xk6xx6, El6xx6, Ll6xx6, Sl6xx6, Zl6xx6, Gm6xx6, Nm6xx6, Um6xx6, Bn6xx6, In6xx6;
wire Pn6xx6, Wn6xx6, Do6xx6, Ko6xx6, Ro6xx6, Yo6xx6, Fp6xx6, Mp6xx6, Tp6xx6, Aq6xx6;
wire Hq6xx6, Oq6xx6, Vq6xx6, Cr6xx6, Jr6xx6, Qr6xx6, Xr6xx6, Es6xx6, Ls6xx6, Ss6xx6;
wire Zs6xx6, Gt6xx6, Nt6xx6, Ut6xx6, Bu6xx6, Iu6xx6, Pu6xx6, Wu6xx6, Dv6xx6, Kv6xx6;
wire Rv6xx6, Yv6xx6, Fw6xx6, Mw6xx6, Tw6xx6, Ax6xx6, Hx6xx6, Ox6xx6, Vx6xx6, Cy6xx6;
wire Jy6xx6, Qy6xx6, Xy6xx6, Ez6xx6, Lz6xx6, Sz6xx6, Zz6xx6, G07xx6, N07xx6, U07xx6;
wire B17xx6, I17xx6, P17xx6, W17xx6, D27xx6, K27xx6, R27xx6, Y27xx6, F37xx6, M37xx6;
wire T37xx6, A47xx6, H47xx6, O47xx6, V47xx6, C57xx6, J57xx6, Q57xx6, X57xx6, E67xx6;
wire L67xx6, S67xx6, Z67xx6, G77xx6, N77xx6, U77xx6, B87xx6, I87xx6, P87xx6, W87xx6;
wire D97xx6, K97xx6, R97xx6, Y97xx6, Fa7xx6, Ma7xx6, Ta7xx6, Ab7xx6, Hb7xx6, Ob7xx6;
wire Vb7xx6, Cc7xx6, Jc7xx6, Qc7xx6, Xc7xx6, Ed7xx6, Ld7xx6, Sd7xx6, Zd7xx6, Ge7xx6;
wire Ne7xx6, Ue7xx6, Bf7xx6, If7xx6, Pf7xx6, Wf7xx6, Dg7xx6, Kg7xx6, Rg7xx6, Yg7xx6;
wire Fh7xx6, Mh7xx6, Th7xx6, Ai7xx6, Hi7xx6, Oi7xx6, Vi7xx6, Cj7xx6, Jj7xx6, Qj7xx6;
wire Xj7xx6, Ek7xx6, Lk7xx6, Sk7xx6, Zk7xx6, Gl7xx6, Nl7xx6, Ul7xx6, Bm7xx6, Im7xx6;
wire Pm7xx6, Wm7xx6, Dn7xx6, Kn7xx6, Rn7xx6, Yn7xx6, Fo7xx6, Mo7xx6, To7xx6, Ap7xx6;
wire Hp7xx6, Op7xx6, Vp7xx6, Cq7xx6, Jq7xx6, Qq7xx6, Xq7xx6, Er7xx6, Lr7xx6, Sr7xx6;
wire Zr7xx6, Gs7xx6, Ns7xx6, Us7xx6, Bt7xx6, It7xx6, Pt7xx6, Wt7xx6, Du7xx6, Ku7xx6;
wire Ru7xx6, Yu7xx6, Fv7xx6, Mv7xx6, Tv7xx6, Aw7xx6, Hw7xx6, Ow7xx6, Vw7xx6, Cx7xx6;
wire Jx7xx6, Qx7xx6, Xx7xx6, Ey7xx6, Ly7xx6, Sy7xx6, Zy7xx6, Gz7xx6, Nz7xx6, Uz7xx6;
wire B08xx6, I08xx6, P08xx6, W08xx6, D18xx6, K18xx6, R18xx6, Y18xx6, F28xx6, M28xx6;
wire T28xx6, A38xx6, H38xx6, O38xx6, V38xx6, C48xx6, J48xx6, Q48xx6, X48xx6, E58xx6;
wire L58xx6, S58xx6, Z58xx6, G68xx6, N68xx6, U68xx6, B78xx6, I78xx6, P78xx6, W78xx6;
wire D88xx6, K88xx6, R88xx6, Y88xx6, F98xx6, M98xx6, T98xx6, Aa8xx6, Ha8xx6, Oa8xx6;
wire Va8xx6, Cb8xx6, Jb8xx6, Qb8xx6, Xb8xx6, Ec8xx6, Lc8xx6, Sc8xx6, Zc8xx6, Gd8xx6;
wire Nd8xx6, Ud8xx6, Be8xx6, Ie8xx6, Pe8xx6, We8xx6, Df8xx6, Kf8xx6, Rf8xx6, Yf8xx6;
wire Fg8xx6, Mg8xx6, Tg8xx6, Ah8xx6, Hh8xx6, Oh8xx6, Vh8xx6, Ci8xx6, Ji8xx6, Qi8xx6;
wire Xi8xx6, Ej8xx6, Lj8xx6, Sj8xx6, Zj8xx6, Gk8xx6, Nk8xx6, Uk8xx6, Bl8xx6, Il8xx6;
wire Pl8xx6, Wl8xx6, Dm8xx6, Km8xx6, Rm8xx6, Ym8xx6, Fn8xx6, Mn8xx6, Tn8xx6, Ao8xx6;
wire Ho8xx6, Oo8xx6, Vo8xx6, Cp8xx6, Jp8xx6, Qp8xx6, Xp8xx6, Eq8xx6, Lq8xx6, Sq8xx6;
wire Zq8xx6, Gr8xx6, Nr8xx6, Ur8xx6, Bs8xx6, Is8xx6, Ps8xx6, Ws8xx6, Dt8xx6, Kt8xx6;
wire Rt8xx6, Yt8xx6, Fu8xx6, Mu8xx6, Tu8xx6, Av8xx6, Hv8xx6, Ov8xx6, Vv8xx6, Cw8xx6;
wire Jw8xx6, Qw8xx6, Xw8xx6, Ex8xx6, Lx8xx6, Sx8xx6, Zx8xx6, Gy8xx6, Ny8xx6, Uy8xx6;
wire Bz8xx6, Iz8xx6, Pz8xx6, Wz8xx6, D09xx6, K09xx6, R09xx6, Y09xx6, F19xx6, M19xx6;
wire T19xx6, A29xx6, H29xx6, O29xx6, V29xx6, C39xx6, J39xx6, Q39xx6, X39xx6, E49xx6;
wire L49xx6, S49xx6, Z49xx6, G59xx6, N59xx6, U59xx6, B69xx6, I69xx6, P69xx6, W69xx6;
wire D79xx6, K79xx6, R79xx6, Y79xx6, F89xx6, M89xx6, T89xx6, A99xx6, H99xx6, O99xx6;
wire V99xx6, Ca9xx6, Ja9xx6, Qa9xx6, Xa9xx6, Eb9xx6, Lb9xx6, Sb9xx6, Zb9xx6, Gc9xx6;
wire Nc9xx6, Uc9xx6, Bd9xx6, Id9xx6, Pd9xx6, Wd9xx6, De9xx6, Ke9xx6, Re9xx6, Ye9xx6;
wire Ff9xx6, Mf9xx6, Tf9xx6, Ag9xx6, Hg9xx6, Og9xx6, Vg9xx6, Ch9xx6, Jh9xx6, Qh9xx6;
wire Xh9xx6, Ei9xx6, Li9xx6, Si9xx6, Zi9xx6, Gj9xx6, Nj9xx6, Uj9xx6, Bk9xx6, Ik9xx6;
wire Pk9xx6, Wk9xx6, Dl9xx6, Kl9xx6, Rl9xx6, Yl9xx6, Fm9xx6, Mm9xx6, Tm9xx6, An9xx6;
wire Hn9xx6, On9xx6, Vn9xx6, Co9xx6, Jo9xx6, Qo9xx6, Xo9xx6, Ep9xx6, Lp9xx6, Sp9xx6;
wire Zp9xx6, Gq9xx6, Nq9xx6, Uq9xx6, Br9xx6, Ir9xx6, Pr9xx6, Wr9xx6, Ds9xx6, Ks9xx6;
wire Rs9xx6, Ys9xx6, Ft9xx6, Mt9xx6, Tt9xx6, Au9xx6, Hu9xx6, Ou9xx6, Vu9xx6, Cv9xx6;
wire Jv9xx6, Qv9xx6, Xv9xx6, Ew9xx6, Lw9xx6, Sw9xx6, Zw9xx6, Gx9xx6, Nx9xx6, Ux9xx6;
wire By9xx6, Iy9xx6, Py9xx6, Wy9xx6, Dz9xx6, Kz9xx6, Rz9xx6, Yz9xx6, F0axx6, M0axx6;
wire T0axx6, A1axx6, H1axx6, O1axx6, V1axx6, C2axx6, J2axx6, Q2axx6, X2axx6, E3axx6;
wire L3axx6, S3axx6, Z3axx6, G4axx6, N4axx6, U4axx6, B5axx6, I5axx6, P5axx6, W5axx6;
wire D6axx6, K6axx6, R6axx6, Y6axx6, F7axx6, M7axx6, T7axx6, A8axx6, H8axx6, O8axx6;
wire V8axx6, C9axx6, J9axx6, Q9axx6, X9axx6, Eaaxx6, Laaxx6, Saaxx6, Zaaxx6, Gbaxx6;
wire Nbaxx6, Ubaxx6, Bcaxx6, Icaxx6, Pcaxx6, Wcaxx6, Ddaxx6, Kdaxx6, Rdaxx6, Ydaxx6;
wire Feaxx6, Meaxx6, Teaxx6, Afaxx6, Hfaxx6, Ofaxx6, Vfaxx6, Cgaxx6, Jgaxx6, Qgaxx6;
wire Xgaxx6, Ehaxx6, Lhaxx6, Shaxx6, Zhaxx6, Giaxx6, Niaxx6, Uiaxx6, Bjaxx6, Ijaxx6;
wire Pjaxx6, Wjaxx6, Dkaxx6, Kkaxx6, Rkaxx6, Ykaxx6, Flaxx6, Mlaxx6, Tlaxx6, Amaxx6;
wire Hmaxx6, Omaxx6, Vmaxx6, Cnaxx6, Jnaxx6, Qnaxx6, Xnaxx6, Eoaxx6, Loaxx6, Soaxx6;
wire Zoaxx6, Gpaxx6, Npaxx6, Upaxx6, Bqaxx6, Iqaxx6, Pqaxx6, Wqaxx6, Draxx6, Kraxx6;
wire Rraxx6, Yraxx6, Fsaxx6, Msaxx6, Tsaxx6, Ataxx6, Htaxx6, Otaxx6, Vtaxx6, Cuaxx6;
wire Juaxx6, Quaxx6, Xuaxx6, Evaxx6, Lvaxx6, Svaxx6, Zvaxx6, Gwaxx6, Nwaxx6, Uwaxx6;
wire Bxaxx6, Ixaxx6, Pxaxx6, Wxaxx6, Dyaxx6, Kyaxx6, Ryaxx6, Yyaxx6, Fzaxx6, Mzaxx6;
wire Tzaxx6, A0bxx6, H0bxx6, O0bxx6, V0bxx6, C1bxx6, J1bxx6, Q1bxx6, X1bxx6, E2bxx6;
wire L2bxx6, S2bxx6, Z2bxx6, G3bxx6, N3bxx6, U3bxx6, B4bxx6, I4bxx6, P4bxx6, W4bxx6;
wire D5bxx6, K5bxx6, R5bxx6, Y5bxx6, F6bxx6, M6bxx6, T6bxx6, A7bxx6, H7bxx6, O7bxx6;
wire V7bxx6, C8bxx6, J8bxx6, Q8bxx6, X8bxx6, E9bxx6, L9bxx6, S9bxx6, Z9bxx6, Gabxx6;
wire Nabxx6, Uabxx6, Bbbxx6, Ibbxx6, Pbbxx6, Wbbxx6, Dcbxx6, Kcbxx6, Rcbxx6, Ycbxx6;
wire Fdbxx6, Mdbxx6, Tdbxx6, Aebxx6, Hebxx6, Oebxx6, Vebxx6, Cfbxx6, Jfbxx6, Qfbxx6;
wire Xfbxx6, Egbxx6, Lgbxx6, Sgbxx6, Zgbxx6, Ghbxx6, Nhbxx6, Uhbxx6, Bibxx6, Iibxx6;
wire Pibxx6, Wibxx6, Djbxx6, Kjbxx6, Rjbxx6, Yjbxx6, Fkbxx6, Mkbxx6, Tkbxx6, Albxx6;
wire Hlbxx6, Olbxx6, Vlbxx6, Cmbxx6, Jmbxx6, Qmbxx6, Xmbxx6, Enbxx6, Lnbxx6, Snbxx6;
wire Znbxx6, Gobxx6, Nobxx6, Uobxx6, Bpbxx6, Ipbxx6, Ppbxx6, Wpbxx6, Dqbxx6, Kqbxx6;
wire Rqbxx6, Yqbxx6, Frbxx6, Mrbxx6, Trbxx6, Asbxx6, Hsbxx6, Osbxx6, Vsbxx6, Ctbxx6;
wire Jtbxx6, Qtbxx6, Xtbxx6, Eubxx6, Lubxx6, Subxx6, Zubxx6, Gvbxx6, Nvbxx6, Uvbxx6;
wire Bwbxx6, Iwbxx6, Pwbxx6, Wwbxx6, Dxbxx6, Kxbxx6, Rxbxx6, Yxbxx6, Fybxx6, Mybxx6;
wire Tybxx6, Azbxx6, Hzbxx6, Ozbxx6, Vzbxx6, C0cxx6, J0cxx6, Q0cxx6, X0cxx6, E1cxx6;
wire L1cxx6, S1cxx6, Z1cxx6, G2cxx6, N2cxx6, U2cxx6, B3cxx6, I3cxx6, P3cxx6, W3cxx6;
wire D4cxx6, K4cxx6, R4cxx6, Y4cxx6, F5cxx6, M5cxx6, T5cxx6, A6cxx6, H6cxx6, O6cxx6;
wire V6cxx6, C7cxx6, J7cxx6, Q7cxx6, X7cxx6, E8cxx6, L8cxx6, S8cxx6, Z8cxx6, G9cxx6;
wire N9cxx6, U9cxx6, Bacxx6, Iacxx6, Pacxx6, Wacxx6, Dbcxx6, Kbcxx6, Rbcxx6, Ybcxx6;
wire Fccxx6, Mccxx6, Tccxx6, Adcxx6, Hdcxx6, Odcxx6, Vdcxx6, Cecxx6, Jecxx6, Qecxx6;
wire Xecxx6, Efcxx6, Lfcxx6, Sfcxx6, Zfcxx6, Ggcxx6, Ngcxx6, Ugcxx6, Bhcxx6, Ihcxx6;
wire Phcxx6, Whcxx6, Dicxx6, Kicxx6, Ricxx6, Yicxx6, Fjcxx6, Mjcxx6, Tjcxx6, Akcxx6;
wire Hkcxx6, Okcxx6, Vkcxx6, Clcxx6, Jlcxx6, Qlcxx6, Xlcxx6, Emcxx6, Lmcxx6, Smcxx6;
wire Zmcxx6, Gncxx6, Nncxx6, Uncxx6, Bocxx6, Iocxx6, Pocxx6, Wocxx6, Dpcxx6, Kpcxx6;
wire Rpcxx6, Ypcxx6, Fqcxx6, Mqcxx6, Tqcxx6, Arcxx6, Hrcxx6, Orcxx6, Vrcxx6, Cscxx6;
wire Jscxx6, Qscxx6, Xscxx6, Etcxx6, Ltcxx6, Stcxx6, Ztcxx6, Gucxx6, Nucxx6, Uucxx6;
wire Bvcxx6, Ivcxx6, Pvcxx6, Wvcxx6, Dwcxx6, Kwcxx6, Rwcxx6, Ywcxx6, Fxcxx6, Mxcxx6;
wire Txcxx6, Aycxx6, Hycxx6, Oycxx6, Vycxx6, Czcxx6, Jzcxx6, Qzcxx6, Xzcxx6, E0dxx6;
wire L0dxx6, S0dxx6, Z0dxx6, G1dxx6, N1dxx6, U1dxx6, B2dxx6, I2dxx6, P2dxx6, W2dxx6;
wire D3dxx6, K3dxx6, R3dxx6, Y3dxx6, F4dxx6, M4dxx6, T4dxx6, A5dxx6, H5dxx6, O5dxx6;
wire V5dxx6, C6dxx6, J6dxx6, Q6dxx6, X6dxx6, E7dxx6, L7dxx6, S7dxx6, Z7dxx6, G8dxx6;
wire N8dxx6, U8dxx6, B9dxx6, I9dxx6, P9dxx6, W9dxx6, Dadxx6, Kadxx6, Radxx6, Yadxx6;
wire Fbdxx6, Mbdxx6, Tbdxx6, Acdxx6, Hcdxx6, Ocdxx6, Vcdxx6, Cddxx6, Jddxx6, Qddxx6;
wire Xddxx6, Eedxx6, Ledxx6, Sedxx6, Zedxx6, Gfdxx6, Nfdxx6, Ufdxx6, Bgdxx6, Igdxx6;
wire Pgdxx6, Wgdxx6, Dhdxx6, Khdxx6, Rhdxx6, Yhdxx6, Fidxx6, Midxx6, Tidxx6, Ajdxx6;
wire Hjdxx6, Ojdxx6, Vjdxx6, Ckdxx6, Jkdxx6, Qkdxx6, Xkdxx6, Eldxx6, Lldxx6, Sldxx6;
wire Zldxx6, Gmdxx6, Nmdxx6, Umdxx6, Bndxx6, Indxx6, Pndxx6, Wndxx6, Dodxx6, Kodxx6;
wire Rodxx6, Yodxx6, Fpdxx6, Mpdxx6, Tpdxx6, Aqdxx6, Hqdxx6, Oqdxx6, Vqdxx6, Crdxx6;
wire Jrdxx6, Qrdxx6, Xrdxx6, Esdxx6, Lsdxx6, Ssdxx6, Zsdxx6, Gtdxx6, Ntdxx6, Utdxx6;
wire Budxx6, Iudxx6, Pudxx6, Wudxx6, Dvdxx6, Kvdxx6, Rvdxx6, Yvdxx6, Fwdxx6, Mwdxx6;
wire Twdxx6, Axdxx6, Hxdxx6, Oxdxx6, Vxdxx6, Cydxx6, Jydxx6, Qydxx6, Xydxx6, Ezdxx6;
wire Lzdxx6, Szdxx6, Zzdxx6, G0exx6, N0exx6, U0exx6, B1exx6, I1exx6, P1exx6, W1exx6;
wire D2exx6, K2exx6, R2exx6, Y2exx6, F3exx6, M3exx6, T3exx6, A4exx6, H4exx6, O4exx6;
wire V4exx6, C5exx6, J5exx6, Q5exx6, X5exx6, E6exx6, L6exx6, S6exx6, Z6exx6, G7exx6;
wire N7exx6, U7exx6, B8exx6, I8exx6, P8exx6, W8exx6, D9exx6, K9exx6, R9exx6, Y9exx6;
wire Faexx6, Maexx6, Taexx6, Abexx6, Hbexx6, Obexx6, Vbexx6, Ccexx6, Jcexx6, Qcexx6;
wire Xcexx6, Edexx6, Ldexx6, Sdexx6, Zdexx6, Geexx6, Neexx6, Ueexx6, Bfexx6, Ifexx6;
wire Pfexx6, Wfexx6, Dgexx6, Kgexx6, Rgexx6, Ygexx6, Fhexx6, Mhexx6, Thexx6, Aiexx6;
wire Hiexx6, Oiexx6, Viexx6, Cjexx6, Jjexx6, Qjexx6, Xjexx6, Ekexx6, Lkexx6, Skexx6;
wire Zkexx6, Glexx6, Nlexx6, Ulexx6, Bmexx6, Imexx6, Pmexx6, Wmexx6, Dnexx6, Knexx6;
wire Rnexx6, Ynexx6, Foexx6, Moexx6, Toexx6, Apexx6, Hpexx6, Opexx6, Vpexx6, Cqexx6;
wire Jqexx6, Qqexx6, Xqexx6, Erexx6, Lrexx6, Srexx6, Zrexx6, Gsexx6, Nsexx6, Usexx6;
wire Btexx6, Itexx6, Ptexx6, Wtexx6, Duexx6, Kuexx6, Ruexx6, Yuexx6, Fvexx6, Mvexx6;
wire Tvexx6, Awexx6, Hwexx6, Owexx6, Vwexx6, Cxexx6, Jxexx6, Qxexx6, Xxexx6, Eyexx6;
wire Lyexx6, Syexx6, Zyexx6, Gzexx6, Nzexx6, Uzexx6, B0fxx6, I0fxx6, P0fxx6, W0fxx6;
wire D1fxx6, K1fxx6, R1fxx6, Y1fxx6, F2fxx6, M2fxx6, T2fxx6, A3fxx6, H3fxx6, O3fxx6;
wire V3fxx6, C4fxx6, J4fxx6, Q4fxx6, X4fxx6, E5fxx6, L5fxx6, S5fxx6, Z5fxx6, G6fxx6;
wire N6fxx6, U6fxx6, B7fxx6, I7fxx6, P7fxx6, W7fxx6, D8fxx6, K8fxx6, R8fxx6, Y8fxx6;
wire F9fxx6, M9fxx6, T9fxx6, Aafxx6, Hafxx6, Oafxx6, Vafxx6, Cbfxx6, Jbfxx6, Qbfxx6;
wire Xbfxx6, Ecfxx6, Lcfxx6, Scfxx6, Zcfxx6, Gdfxx6, Ndfxx6, Udfxx6, Befxx6, Iefxx6;
wire Pefxx6, Wefxx6, Dffxx6, Kffxx6, Rffxx6, Yffxx6, Fgfxx6, Mgfxx6, Tgfxx6, Ahfxx6;
wire Hhfxx6, Ohfxx6, Vhfxx6, Cifxx6, Jifxx6, Qifxx6, Xifxx6, Ejfxx6, Ljfxx6, Sjfxx6;
wire Zjfxx6, Gkfxx6, Nkfxx6, Ukfxx6, Blfxx6, Ilfxx6, Plfxx6, Wlfxx6, Dmfxx6, Kmfxx6;
wire Rmfxx6, Ymfxx6, Fnfxx6, Mnfxx6, Tnfxx6, Aofxx6, Hofxx6, Oofxx6, Vofxx6, Cpfxx6;
wire Jpfxx6, Qpfxx6, Xpfxx6, Eqfxx6, Lqfxx6, Sqfxx6, Zqfxx6, Grfxx6, Nrfxx6, Urfxx6;
wire Bsfxx6, Isfxx6, Psfxx6, Wsfxx6, Dtfxx6, Ktfxx6, Rtfxx6, Ytfxx6, Fufxx6, Mufxx6;
wire Tufxx6, Avfxx6, Hvfxx6, Ovfxx6, Vvfxx6, Cwfxx6, Jwfxx6, Qwfxx6, Xwfxx6, Exfxx6;
wire Lxfxx6, Sxfxx6, Zxfxx6, Gyfxx6, Nyfxx6, Uyfxx6, Bzfxx6, Izfxx6, Pzfxx6, Wzfxx6;
wire D0gxx6, K0gxx6, R0gxx6, Y0gxx6, F1gxx6, M1gxx6, T1gxx6, A2gxx6, H2gxx6, O2gxx6;
wire V2gxx6, C3gxx6, J3gxx6, Q3gxx6, X3gxx6, E4gxx6, L4gxx6, S4gxx6, Z4gxx6, G5gxx6;
wire N5gxx6, U5gxx6, B6gxx6, I6gxx6, P6gxx6, W6gxx6, D7gxx6, K7gxx6, R7gxx6, Y7gxx6;
wire F8gxx6, M8gxx6, T8gxx6, A9gxx6, H9gxx6, O9gxx6, V9gxx6, Cagxx6, Jagxx6, Qagxx6;
wire Xagxx6, Ebgxx6, Lbgxx6, Sbgxx6, Zbgxx6, Gcgxx6, Ncgxx6, Ucgxx6, Bdgxx6, Idgxx6;
wire Pdgxx6, Wdgxx6, Degxx6, Kegxx6, Regxx6, Yegxx6, Ffgxx6, Mfgxx6, Tfgxx6, Aggxx6;
wire Hggxx6, Oggxx6, Vggxx6, Chgxx6, Jhgxx6, Qhgxx6, Xhgxx6, Eigxx6, Ligxx6, Sigxx6;
wire Zigxx6, Gjgxx6, Njgxx6, Ujgxx6, Bkgxx6, Ikgxx6, Pkgxx6, Wkgxx6, Dlgxx6, Klgxx6;
wire Rlgxx6, Ylgxx6, Fmgxx6, Mmgxx6, Tmgxx6, Angxx6, Hngxx6, Ongxx6, Vngxx6, Cogxx6;
wire Jogxx6, Qogxx6, Xogxx6, Epgxx6, Lpgxx6, Spgxx6, Zpgxx6, Gqgxx6, Nqgxx6, Uqgxx6;
wire Brgxx6, Irgxx6, Prgxx6, Wrgxx6, Dsgxx6, Ksgxx6, Rsgxx6, Ysgxx6, Ftgxx6, Mtgxx6;
wire Ttgxx6, Augxx6, Hugxx6, Ougxx6, Vugxx6, Cvgxx6, Jvgxx6, Qvgxx6, Xvgxx6, Ewgxx6;
wire Lwgxx6, Swgxx6, Zwgxx6, Gxgxx6, Nxgxx6, Uxgxx6, Bygxx6, Iygxx6, Pygxx6, Wygxx6;
wire Dzgxx6, Kzgxx6, Rzgxx6, Yzgxx6, F0hxx6, M0hxx6, T0hxx6, A1hxx6, H1hxx6, O1hxx6;
wire V1hxx6, C2hxx6, J2hxx6, Q2hxx6, X2hxx6, E3hxx6, L3hxx6, S3hxx6, Z3hxx6, G4hxx6;
wire N4hxx6, U4hxx6, B5hxx6, I5hxx6, P5hxx6, W5hxx6, D6hxx6, K6hxx6, R6hxx6, Y6hxx6;
wire F7hxx6, M7hxx6, T7hxx6, A8hxx6, H8hxx6, O8hxx6, V8hxx6, C9hxx6, J9hxx6, Q9hxx6;
wire X9hxx6, Eahxx6, Lahxx6, Sahxx6, Zahxx6, Gbhxx6, Nbhxx6, Ubhxx6, Bchxx6, Ichxx6;
wire Pchxx6, Wchxx6, Ddhxx6, Kdhxx6, Rdhxx6, Ydhxx6, Fehxx6, Mehxx6, Tehxx6, Afhxx6;
wire Hfhxx6, Ofhxx6, Vfhxx6, Cghxx6, Jghxx6, Qghxx6, Xghxx6, Ehhxx6, Lhhxx6, Shhxx6;
wire Zhhxx6, Gihxx6, Nihxx6, Uihxx6, Bjhxx6, Ijhxx6, Pjhxx6, Wjhxx6, Dkhxx6, Kkhxx6;
wire Rkhxx6, Ykhxx6, Flhxx6, Mlhxx6, Tlhxx6, Amhxx6, Hmhxx6, Omhxx6, Vmhxx6, Cnhxx6;
wire Jnhxx6, Qnhxx6, Xnhxx6, Eohxx6, Lohxx6, Sohxx6, Zohxx6, Gphxx6, Nphxx6, Uphxx6;
wire Bqhxx6, Iqhxx6, Pqhxx6, Wqhxx6, Drhxx6, Krhxx6, Rrhxx6, Yrhxx6, Fshxx6, Mshxx6;
wire Tshxx6, Athxx6, Hthxx6, Othxx6, Vthxx6, Cuhxx6, Juhxx6, Quhxx6, Xuhxx6, Evhxx6;
wire Lvhxx6, Svhxx6, Zvhxx6, Gwhxx6, Nwhxx6, Uwhxx6, Bxhxx6, Ixhxx6, Pxhxx6, Wxhxx6;
wire Dyhxx6, Kyhxx6, Ryhxx6, Yyhxx6, Fzhxx6, Mzhxx6, Tzhxx6, A0ixx6, H0ixx6, O0ixx6;
wire V0ixx6, C1ixx6, J1ixx6, Q1ixx6, X1ixx6, E2ixx6, L2ixx6, S2ixx6, Z2ixx6, G3ixx6;
wire N3ixx6, U3ixx6, B4ixx6, I4ixx6, P4ixx6, W4ixx6, D5ixx6, K5ixx6, R5ixx6, Y5ixx6;
wire F6ixx6, M6ixx6, T6ixx6, A7ixx6, H7ixx6, O7ixx6, V7ixx6, C8ixx6, J8ixx6, Q8ixx6;
wire X8ixx6, E9ixx6, L9ixx6, S9ixx6, Z9ixx6, Gaixx6, Naixx6, Uaixx6, Bbixx6, Ibixx6;
wire Pbixx6, Wbixx6, Dcixx6, Kcixx6, Rcixx6, Ycixx6, Fdixx6, Mdixx6, Tdixx6, Aeixx6;
wire Heixx6, Oeixx6, Veixx6, Cfixx6, Jfixx6, Qfixx6, Xfixx6, Egixx6, Lgixx6, Sgixx6;
wire Zgixx6, Ghixx6, Nhixx6, Uhixx6, Biixx6, Iiixx6, Piixx6, Wiixx6, Djixx6, Kjixx6;
wire Rjixx6, Yjixx6, Fkixx6, Mkixx6, Tkixx6, Alixx6, Hlixx6, Olixx6, Vlixx6, Cmixx6;
wire Jmixx6, Qmixx6, Xmixx6, Enixx6, Lnixx6, Snixx6, Znixx6, Goixx6, Noixx6, Uoixx6;
wire Bpixx6, Ipixx6, Ppixx6, Wpixx6, Dqixx6, Kqixx6, Rqixx6, Yqixx6, Frixx6, Mrixx6;
wire Trixx6, Asixx6, Hsixx6, Osixx6, Vsixx6, Ctixx6, Jtixx6, Qtixx6, Xtixx6, Euixx6;
wire Luixx6, Suixx6, Zuixx6, Gvixx6, Nvixx6, Uvixx6, Bwixx6, Iwixx6, Pwixx6, Wwixx6;
wire Dxixx6, Kxixx6, Rxixx6, Yxixx6, Fyixx6, Myixx6, Tyixx6, Azixx6, Hzixx6, Ozixx6;
wire Vzixx6, C0jxx6, J0jxx6, Q0jxx6, X0jxx6, E1jxx6, L1jxx6, S1jxx6, Z1jxx6, G2jxx6;
wire N2jxx6, U2jxx6, B3jxx6, I3jxx6, P3jxx6, W3jxx6, D4jxx6, K4jxx6, R4jxx6, Y4jxx6;
wire F5jxx6, M5jxx6, T5jxx6, A6jxx6, H6jxx6, O6jxx6, V6jxx6, C7jxx6, J7jxx6, Q7jxx6;
wire X7jxx6, E8jxx6, L8jxx6, S8jxx6, Z8jxx6, G9jxx6, N9jxx6, U9jxx6, Bajxx6, Iajxx6;
wire Pajxx6, Wajxx6, Dbjxx6, Kbjxx6, Rbjxx6, Ybjxx6, Fcjxx6, Mcjxx6, Tcjxx6, Adjxx6;
wire Hdjxx6, Odjxx6, Vdjxx6, Cejxx6, Jejxx6, Qejxx6, Xejxx6, Efjxx6, Lfjxx6, Sfjxx6;
wire Zfjxx6, Ggjxx6, Ngjxx6, Ugjxx6, Bhjxx6, Ihjxx6, Phjxx6, Whjxx6, Dijxx6, Kijxx6;
wire Rijxx6, Yijxx6, Fjjxx6, Mjjxx6, Tjjxx6, Akjxx6, Hkjxx6, Okjxx6, Vkjxx6, Cljxx6;
wire Jljxx6, Qljxx6, Xljxx6, Emjxx6, Lmjxx6, Smjxx6, Zmjxx6, Gnjxx6, Nnjxx6, Unjxx6;
wire Bojxx6, Iojxx6, Pojxx6, Wojxx6, Dpjxx6, Kpjxx6, Rpjxx6, Ypjxx6, Fqjxx6, Mqjxx6;
wire Tqjxx6, Arjxx6, Hrjxx6, Orjxx6, Vrjxx6, Csjxx6, Jsjxx6, Qsjxx6, Xsjxx6, Etjxx6;
wire Ltjxx6, Stjxx6, Ztjxx6, Gujxx6, Nujxx6, Uujxx6, Bvjxx6, Ivjxx6, Pvjxx6, Wvjxx6;
wire Dwjxx6, Kwjxx6, Rwjxx6, Ywjxx6, Fxjxx6, Mxjxx6, Txjxx6, Ayjxx6, Hyjxx6, Oyjxx6;
wire Vyjxx6, Czjxx6, Jzjxx6, Qzjxx6, Xzjxx6, E0kxx6, L0kxx6, S0kxx6, Z0kxx6, G1kxx6;
wire N1kxx6, U1kxx6, B2kxx6, I2kxx6, P2kxx6, W2kxx6, D3kxx6, K3kxx6, R3kxx6, Y3kxx6;
wire F4kxx6, M4kxx6, T4kxx6, A5kxx6, H5kxx6, O5kxx6, V5kxx6, C6kxx6, J6kxx6, Q6kxx6;
wire X6kxx6, E7kxx6, L7kxx6, S7kxx6, Z7kxx6, G8kxx6, N8kxx6, U8kxx6, B9kxx6, I9kxx6;
wire P9kxx6, W9kxx6, Dakxx6, Kakxx6, Rakxx6, Yakxx6, Fbkxx6, Mbkxx6, Tbkxx6, Ackxx6;
wire Hckxx6, Ockxx6, Vckxx6, Cdkxx6, Jdkxx6, Qdkxx6, Xdkxx6, Eekxx6, Lekxx6, Sekxx6;
wire Zekxx6, Gfkxx6, Nfkxx6, Ufkxx6, Bgkxx6, Igkxx6, Pgkxx6, Wgkxx6, Dhkxx6, Khkxx6;
wire Rhkxx6, Yhkxx6, Fikxx6, Mikxx6, Tikxx6, Ajkxx6, Hjkxx6, Ojkxx6, Vjkxx6, Ckkxx6;
wire Jkkxx6, Qkkxx6, Xkkxx6, Elkxx6, Llkxx6, Slkxx6, Zlkxx6, Gmkxx6, Nmkxx6, Umkxx6;
wire Bnkxx6, Inkxx6, Pnkxx6, Wnkxx6, Dokxx6, Kokxx6, Rokxx6, Yokxx6, Fpkxx6, Mpkxx6;
wire Tpkxx6, Aqkxx6, Hqkxx6, Oqkxx6, Vqkxx6, Crkxx6, Jrkxx6, Qrkxx6, Xrkxx6, Eskxx6;
wire Lskxx6, Sskxx6, Zskxx6, Gtkxx6, Ntkxx6, Utkxx6, Bukxx6, Iukxx6, Pukxx6, Wukxx6;
wire Dvkxx6, Kvkxx6, Rvkxx6, Yvkxx6, Fwkxx6, Mwkxx6, Twkxx6, Axkxx6, Hxkxx6, Oxkxx6;
wire Vxkxx6, Cykxx6, Jykxx6, Qykxx6, Xykxx6, Ezkxx6, Lzkxx6, Szkxx6, Zzkxx6, G0lxx6;
wire N0lxx6, U0lxx6, B1lxx6, I1lxx6, P1lxx6, W1lxx6, D2lxx6, K2lxx6, R2lxx6, Y2lxx6;
wire F3lxx6, M3lxx6, T3lxx6, A4lxx6, H4lxx6, O4lxx6, V4lxx6, C5lxx6, J5lxx6, Q5lxx6;
wire X5lxx6, E6lxx6, L6lxx6, S6lxx6, Z6lxx6, G7lxx6, N7lxx6, U7lxx6, B8lxx6, I8lxx6;
wire P8lxx6, W8lxx6, D9lxx6, K9lxx6, R9lxx6, Y9lxx6, Falxx6, Malxx6, Talxx6, Ablxx6;
wire Hblxx6, Oblxx6, Vblxx6, Cclxx6, Jclxx6, Qclxx6, Xclxx6, Edlxx6, Ldlxx6, Sdlxx6;
wire Zdlxx6, Gelxx6, Nelxx6, Uelxx6, Bflxx6, Iflxx6, Pflxx6, Wflxx6, Dglxx6, Kglxx6;
wire Rglxx6, Yglxx6, Fhlxx6, Mhlxx6, Thlxx6, Ailxx6, Hilxx6, Oilxx6, Vilxx6, Cjlxx6;
wire Jjlxx6, Qjlxx6, Xjlxx6, Eklxx6, Lklxx6, Sklxx6, Zklxx6, Gllxx6, Nllxx6, Ullxx6;
wire Bmlxx6, Imlxx6, Pmlxx6, Wmlxx6, Dnlxx6, Knlxx6, Rnlxx6, Ynlxx6, Folxx6, Molxx6;
wire Tolxx6, Aplxx6, Hplxx6, Oplxx6, Vplxx6, Cqlxx6, Jqlxx6, Qqlxx6, Xqlxx6, Erlxx6;
wire Lrlxx6, Srlxx6, Zrlxx6, Gslxx6, Nslxx6, Uslxx6, Btlxx6, Itlxx6, Ptlxx6, Wtlxx6;
wire Dulxx6, Kulxx6, Rulxx6, Yulxx6, Fvlxx6, Mvlxx6, Tvlxx6, Awlxx6, Hwlxx6, Owlxx6;
wire Vwlxx6, Cxlxx6, Jxlxx6, Qxlxx6, Xxlxx6, Eylxx6, Lylxx6, Sylxx6, Zylxx6, Gzlxx6;
wire Nzlxx6, Uzlxx6, B0mxx6, I0mxx6, P0mxx6, W0mxx6, D1mxx6, K1mxx6, R1mxx6, Y1mxx6;
wire F2mxx6, M2mxx6, T2mxx6, A3mxx6, H3mxx6, O3mxx6, V3mxx6, C4mxx6, J4mxx6, Q4mxx6;
wire X4mxx6, E5mxx6, L5mxx6, S5mxx6, Z5mxx6, G6mxx6, N6mxx6, U6mxx6, B7mxx6, I7mxx6;
wire P7mxx6, W7mxx6, D8mxx6, K8mxx6, R8mxx6, Y8mxx6, F9mxx6, M9mxx6, T9mxx6, Aamxx6;
wire Hamxx6, Oamxx6, Vamxx6, Cbmxx6, Jbmxx6, Qbmxx6, Xbmxx6, Ecmxx6, Lcmxx6, Scmxx6;
wire Zcmxx6, Gdmxx6, Ndmxx6, Udmxx6, Bemxx6, Iemxx6, Pemxx6, Wemxx6, Dfmxx6, Kfmxx6;
wire Rfmxx6, Yfmxx6, Fgmxx6, Mgmxx6, Tgmxx6, Ahmxx6, Hhmxx6, Ohmxx6, Vhmxx6, Cimxx6;
wire Jimxx6, Qimxx6, Ximxx6, Ejmxx6, Ljmxx6, Sjmxx6, Zjmxx6, Gkmxx6, Nkmxx6, Ukmxx6;
wire Blmxx6, Ilmxx6, Plmxx6, Wlmxx6, Dmmxx6, Kmmxx6, Rmmxx6, Ymmxx6, Fnmxx6, Mnmxx6;
wire Tnmxx6, Aomxx6, Homxx6, Oomxx6, Vomxx6, Cpmxx6, Jpmxx6, Qpmxx6, Xpmxx6, Eqmxx6;
wire Lqmxx6, Sqmxx6, Zqmxx6, Grmxx6, Nrmxx6, Urmxx6, Bsmxx6, Ismxx6, Psmxx6, Wsmxx6;
wire Dtmxx6, Ktmxx6, Rtmxx6, Ytmxx6, Fumxx6, Mumxx6, Tumxx6, Avmxx6, Hvmxx6, Ovmxx6;
wire Vvmxx6, Cwmxx6, Jwmxx6, Qwmxx6, Xwmxx6, Exmxx6, Lxmxx6, Sxmxx6, Zxmxx6, Gymxx6;
wire Nymxx6, Uymxx6, Bzmxx6, Izmxx6, Pzmxx6, Wzmxx6, D0nxx6, K0nxx6, R0nxx6, Y0nxx6;
wire F1nxx6, M1nxx6, T1nxx6, A2nxx6, H2nxx6, O2nxx6, V2nxx6, C3nxx6, J3nxx6, Q3nxx6;
wire X3nxx6, E4nxx6, L4nxx6, S4nxx6, Z4nxx6, G5nxx6, N5nxx6, U5nxx6, B6nxx6, I6nxx6;
wire P6nxx6, W6nxx6, D7nxx6, K7nxx6, R7nxx6, Y7nxx6, F8nxx6, M8nxx6, T8nxx6, A9nxx6;
wire H9nxx6, O9nxx6, V9nxx6, Canxx6, Janxx6, Qanxx6, Xanxx6, Ebnxx6, Lbnxx6, Sbnxx6;
wire Zbnxx6, Gcnxx6, Ncnxx6, Ucnxx6, Bdnxx6, Idnxx6, Pdnxx6, Wdnxx6, Denxx6, Kenxx6;
wire Renxx6, Yenxx6, Ffnxx6, Mfnxx6, Tfnxx6, Agnxx6, Hgnxx6, Ognxx6, Vgnxx6, Chnxx6;
wire Jhnxx6, Qhnxx6, Xhnxx6, Einxx6, Linxx6, Sinxx6, Zinxx6, Gjnxx6, Njnxx6, Ujnxx6;
wire Bknxx6, Iknxx6, Pknxx6, Wknxx6, Dlnxx6, Klnxx6, Rlnxx6, Ylnxx6, Fmnxx6, Mmnxx6;
wire Tmnxx6, Annxx6, Hnnxx6, Onnxx6, Vnnxx6, Conxx6, Jonxx6, Qonxx6, Xonxx6, Epnxx6;
wire Lpnxx6, Spnxx6, Zpnxx6, Gqnxx6, Nqnxx6, Uqnxx6, Brnxx6, Irnxx6, Prnxx6, Wrnxx6;
wire Dsnxx6, Ksnxx6, Rsnxx6, Ysnxx6, Ftnxx6, Mtnxx6, Ttnxx6, Aunxx6, Hunxx6, Ounxx6;
wire Vunxx6, Cvnxx6, Jvnxx6, Qvnxx6, Xvnxx6, Ewnxx6, Lwnxx6, Swnxx6, Zwnxx6, Gxnxx6;
wire Nxnxx6, Uxnxx6, Bynxx6, Iynxx6, Pynxx6, Wynxx6, Dznxx6, Kznxx6, Rznxx6, Yznxx6;
wire F0oxx6, M0oxx6, T0oxx6, A1oxx6, H1oxx6, O1oxx6, V1oxx6, C2oxx6, J2oxx6, Q2oxx6;
wire X2oxx6, E3oxx6, L3oxx6, S3oxx6, Z3oxx6, G4oxx6, N4oxx6, U4oxx6, B5oxx6, I5oxx6;
wire P5oxx6, W5oxx6, D6oxx6, K6oxx6, R6oxx6, Y6oxx6, F7oxx6, M7oxx6, T7oxx6, A8oxx6;
wire H8oxx6, O8oxx6, V8oxx6, C9oxx6, J9oxx6, Q9oxx6, X9oxx6, Eaoxx6, Laoxx6, Saoxx6;
wire Zaoxx6, Gboxx6, Nboxx6, Uboxx6, Bcoxx6, Icoxx6, Pcoxx6, Wcoxx6, Ddoxx6, Kdoxx6;
wire Rdoxx6, Ydoxx6, Feoxx6, Meoxx6, Teoxx6, Afoxx6, Hfoxx6, Ofoxx6, Vfoxx6, Cgoxx6;
wire Jgoxx6, Qgoxx6, Xgoxx6, Ehoxx6, Lhoxx6, Shoxx6, Zhoxx6, Gioxx6, Nioxx6, Uioxx6;
wire Bjoxx6, Ijoxx6, Pjoxx6, Wjoxx6, Dkoxx6, Kkoxx6, Rkoxx6, Ykoxx6, Floxx6, Mloxx6;
wire Tloxx6, Amoxx6, Hmoxx6, Omoxx6, Vmoxx6, Cnoxx6, Jnoxx6, Qnoxx6, Xnoxx6, Eooxx6;
wire Looxx6, Sooxx6, Zooxx6, Gpoxx6, Npoxx6, Upoxx6, Bqoxx6, Iqoxx6, Pqoxx6, Wqoxx6;
wire Droxx6, Kroxx6, Rroxx6, Yroxx6, Fsoxx6, Msoxx6, Tsoxx6, Atoxx6, Htoxx6, Otoxx6;
wire Vtoxx6, Cuoxx6, Juoxx6, Quoxx6, Xuoxx6, Evoxx6, Lvoxx6, Svoxx6, Zvoxx6, Gwoxx6;
wire Nwoxx6, Uwoxx6, Bxoxx6, Ixoxx6, Pxoxx6, Wxoxx6, Dyoxx6, Kyoxx6, Ryoxx6, Yyoxx6;
wire Fzoxx6, Mzoxx6, Tzoxx6, A0pxx6, H0pxx6, O0pxx6, V0pxx6, C1pxx6, J1pxx6, Q1pxx6;
wire X1pxx6, E2pxx6, L2pxx6, S2pxx6, Z2pxx6, G3pxx6, N3pxx6, U3pxx6, B4pxx6, I4pxx6;
wire P4pxx6, W4pxx6, D5pxx6, K5pxx6, R5pxx6, Y5pxx6, F6pxx6, M6pxx6, T6pxx6, A7pxx6;
wire H7pxx6, O7pxx6, V7pxx6, C8pxx6, J8pxx6, Q8pxx6, X8pxx6, E9pxx6, L9pxx6, S9pxx6;
wire Z9pxx6, Gapxx6, Napxx6, Uapxx6, Bbpxx6, Ibpxx6, Pbpxx6, Wbpxx6, Dcpxx6, Kcpxx6;
wire Rcpxx6, Ycpxx6, Fdpxx6, Mdpxx6, Tdpxx6, Aepxx6, Hepxx6, Oepxx6, Vepxx6, Cfpxx6;
wire Jfpxx6, Qfpxx6, Xfpxx6, Egpxx6, Lgpxx6, Sgpxx6, Zgpxx6, Ghpxx6, Nhpxx6, Uhpxx6;
wire Bipxx6, Iipxx6, Pipxx6, Wipxx6, Djpxx6, Kjpxx6, Rjpxx6, Yjpxx6, Fkpxx6, Mkpxx6;
wire Tkpxx6, Alpxx6, Hlpxx6, Olpxx6, Vlpxx6, Cmpxx6, Jmpxx6, Qmpxx6, Xmpxx6, Enpxx6;
wire Lnpxx6, Snpxx6, Znpxx6, Gopxx6, Nopxx6, Uopxx6, Bppxx6, Ippxx6, Pppxx6, Wppxx6;
wire Dqpxx6, Kqpxx6, Rqpxx6, Yqpxx6, Frpxx6, Mrpxx6, Trpxx6, Aspxx6, Hspxx6, Ospxx6;
wire Vspxx6, Ctpxx6, Jtpxx6, Qtpxx6, Xtpxx6, Eupxx6, Lupxx6, Supxx6, Zupxx6, Gvpxx6;
wire Nvpxx6, Uvpxx6, Bwpxx6, Iwpxx6, Pwpxx6, Wwpxx6, Dxpxx6, Kxpxx6, Rxpxx6, Yxpxx6;
wire Fypxx6, Mypxx6, Typxx6, Azpxx6, Hzpxx6, Ozpxx6, Vzpxx6, C0qxx6, J0qxx6, Q0qxx6;
wire X0qxx6, E1qxx6, L1qxx6, S1qxx6, Z1qxx6, G2qxx6, N2qxx6, U2qxx6, B3qxx6, I3qxx6;
wire P3qxx6, W3qxx6, D4qxx6, K4qxx6, R4qxx6, Y4qxx6, F5qxx6, M5qxx6, T5qxx6, A6qxx6;
wire H6qxx6, O6qxx6, V6qxx6, C7qxx6, J7qxx6, Q7qxx6, X7qxx6, E8qxx6, L8qxx6, S8qxx6;
wire Z8qxx6, G9qxx6, N9qxx6, U9qxx6, Baqxx6, Iaqxx6, Paqxx6, Waqxx6, Dbqxx6, Kbqxx6;
wire Rbqxx6, Ybqxx6, Fcqxx6, Mcqxx6, Tcqxx6, Adqxx6, Hdqxx6, Odqxx6, Vdqxx6, Ceqxx6;
wire Jeqxx6, Qeqxx6, Xeqxx6, Efqxx6, Lfqxx6, Sfqxx6, Zfqxx6, Ggqxx6, Ngqxx6, Ugqxx6;
wire Bhqxx6, Ihqxx6, Phqxx6, Whqxx6, Diqxx6, Kiqxx6, Riqxx6, Yiqxx6, Fjqxx6, Mjqxx6;
wire Tjqxx6, Akqxx6, Hkqxx6, Okqxx6, Vkqxx6, Clqxx6, Jlqxx6, Qlqxx6, Xlqxx6, Emqxx6;
wire Lmqxx6, Smqxx6, Zmqxx6, Gnqxx6, Nnqxx6, Unqxx6, Boqxx6, Ioqxx6, Poqxx6, Woqxx6;
wire Dpqxx6, Kpqxx6, Rpqxx6, Ypqxx6, Fqqxx6, Mqqxx6, Tqqxx6, Arqxx6, Hrqxx6, Orqxx6;
wire Vrqxx6, Csqxx6, Jsqxx6, Qsqxx6, Xsqxx6, Etqxx6, Ltqxx6, Stqxx6, Ztqxx6, Guqxx6;
wire Nuqxx6, Uuqxx6, Bvqxx6, Ivqxx6, Pvqxx6, Wvqxx6, Dwqxx6, Kwqxx6, Rwqxx6, Ywqxx6;
wire Fxqxx6, Mxqxx6, Txqxx6, Ayqxx6, Hyqxx6, Oyqxx6, Vyqxx6, Czqxx6, Jzqxx6, Qzqxx6;
wire Xzqxx6, E0rxx6, L0rxx6, S0rxx6, Z0rxx6, G1rxx6, N1rxx6, U1rxx6, B2rxx6, I2rxx6;
wire P2rxx6, W2rxx6, D3rxx6, K3rxx6, R3rxx6, Y3rxx6, F4rxx6, M4rxx6, T4rxx6, A5rxx6;
wire H5rxx6, O5rxx6, V5rxx6, C6rxx6, J6rxx6, Q6rxx6, X6rxx6, E7rxx6, L7rxx6, S7rxx6;
wire Z7rxx6, G8rxx6, N8rxx6, U8rxx6, B9rxx6, I9rxx6, P9rxx6, W9rxx6, Darxx6, Karxx6;
wire Rarxx6, Yarxx6, Fbrxx6, Mbrxx6, Tbrxx6, Acrxx6, Hcrxx6, Ocrxx6, Vcrxx6, Cdrxx6;
wire Jdrxx6, Qdrxx6, Xdrxx6, Eerxx6, Lerxx6, Serxx6, Zerxx6, Gfrxx6, Nfrxx6, Ufrxx6;
wire Bgrxx6, Igrxx6, Pgrxx6, Wgrxx6, Dhrxx6, Khrxx6, Rhrxx6, Yhrxx6, Firxx6, Mirxx6;
wire Tirxx6, Ajrxx6, Hjrxx6, Ojrxx6, Vjrxx6, Ckrxx6, Jkrxx6, Qkrxx6, Xkrxx6, Elrxx6;
wire Llrxx6, Slrxx6, Zlrxx6, Gmrxx6, Nmrxx6, Umrxx6, Bnrxx6, Inrxx6, Pnrxx6, Wnrxx6;
wire Dorxx6, Korxx6, Rorxx6, Yorxx6, Fprxx6, Mprxx6, Tprxx6, Aqrxx6, Hqrxx6, Oqrxx6;
wire Vqrxx6, Crrxx6, Jrrxx6, Qrrxx6, Xrrxx6, Esrxx6, Lsrxx6, Ssrxx6, Zsrxx6, Gtrxx6;
wire Ntrxx6, Utrxx6, Burxx6, Iurxx6, Purxx6, Wurxx6, Dvrxx6, Kvrxx6, Rvrxx6, Yvrxx6;
wire Fwrxx6, Mwrxx6, Twrxx6, Axrxx6, Hxrxx6, Oxrxx6, Vxrxx6, Cyrxx6, Jyrxx6, Qyrxx6;
wire Xyrxx6, Ezrxx6, Lzrxx6, Szrxx6, Zzrxx6, G0sxx6, N0sxx6, U0sxx6, B1sxx6, I1sxx6;
wire P1sxx6, W1sxx6, D2sxx6, K2sxx6, R2sxx6, Y2sxx6, F3sxx6, M3sxx6, T3sxx6, A4sxx6;
wire H4sxx6, O4sxx6, V4sxx6, C5sxx6, J5sxx6, Q5sxx6, X5sxx6, E6sxx6, L6sxx6, S6sxx6;
wire Z6sxx6, G7sxx6, N7sxx6, U7sxx6, B8sxx6, I8sxx6, P8sxx6, W8sxx6, D9sxx6, K9sxx6;
wire R9sxx6, Y9sxx6, Fasxx6, Masxx6, Tasxx6, Absxx6, Hbsxx6, Obsxx6, Vbsxx6, Ccsxx6;
wire Jcsxx6, Qcsxx6, Xcsxx6, Edsxx6, Ldsxx6, Sdsxx6, Zdsxx6, Gesxx6, Nesxx6, Uesxx6;
wire Bfsxx6, Ifsxx6, Pfsxx6, Wfsxx6, Dgsxx6, Kgsxx6, Rgsxx6, Ygsxx6, Fhsxx6, Mhsxx6;
wire Thsxx6, Aisxx6, Hisxx6, Oisxx6, Visxx6, Cjsxx6, Jjsxx6, Qjsxx6, Xjsxx6, Eksxx6;
wire Lksxx6, Sksxx6, Zksxx6, Glsxx6, Nlsxx6, Ulsxx6, Bmsxx6, Imsxx6, Pmsxx6, Wmsxx6;
wire Dnsxx6, Knsxx6, Rnsxx6, Ynsxx6, Fosxx6, Mosxx6, Tosxx6, Apsxx6, Hpsxx6, Opsxx6;
wire Vpsxx6, Cqsxx6, Jqsxx6, Qqsxx6, Xqsxx6, Ersxx6, Lrsxx6, Srsxx6, Zrsxx6, Gssxx6;
wire Nssxx6, Vssxx6, Dtsxx6, Ltsxx6, Ttsxx6, Busxx6, Jusxx6, Rusxx6, Zusxx6, Hvsxx6;
wire Pvsxx6, Xvsxx6, Fwsxx6, Nwsxx6, Vwsxx6, Dxsxx6, Lxsxx6, Txsxx6, Bysxx6, Jysxx6;
wire Rysxx6, Zysxx6, Hzsxx6, Pzsxx6, Xzsxx6, F0txx6, N0txx6, V0txx6, D1txx6, L1txx6;
wire T1txx6, B2txx6, J2txx6, R2txx6, Z2txx6, H3txx6, P3txx6, X3txx6, F4txx6, N4txx6;
wire V4txx6, D5txx6, L5txx6, T5txx6, B6txx6, J6txx6, R6txx6, Z6txx6, H7txx6, P7txx6;
wire X7txx6, F8txx6, N8txx6, V8txx6, D9txx6, L9txx6, T9txx6, Batxx6, Jatxx6, Ratxx6;
wire Zatxx6, Hbtxx6, Pbtxx6, Xbtxx6, Fctxx6, Nctxx6, Vctxx6, Ddtxx6, Ldtxx6, Tdtxx6;
wire Betxx6, Jetxx6, Retxx6, Zetxx6, Hftxx6, Pftxx6, Xftxx6, Fgtxx6, Ngtxx6, Vgtxx6;
wire Dhtxx6, Lhtxx6, Thtxx6, Bitxx6, Jitxx6, Ritxx6, Zitxx6, Hjtxx6, Pjtxx6, Xjtxx6;
wire Fktxx6, Nktxx6, Vktxx6, Dltxx6, Lltxx6, Tltxx6, Bmtxx6, Jmtxx6, Rmtxx6, Zmtxx6;
wire Hntxx6, Pntxx6, Xntxx6, Fotxx6, Notxx6, Votxx6, Dptxx6, Lptxx6, Tptxx6, Bqtxx6;
wire Jqtxx6, Rqtxx6, Zqtxx6, Hrtxx6, Prtxx6, Xrtxx6, Fstxx6, Nstxx6, Vstxx6, Dttxx6;
wire Lttxx6, Tttxx6, Butxx6, Jutxx6, Rutxx6, Zutxx6, Hvtxx6, Pvtxx6, Xvtxx6, Fwtxx6;
wire Nwtxx6, Vwtxx6, Dxtxx6, Lxtxx6, Txtxx6, Bytxx6, Jytxx6, Rytxx6, Zytxx6, Hztxx6;
wire Pztxx6, Xztxx6, F0uxx6, N0uxx6, V0uxx6, D1uxx6, L1uxx6, T1uxx6, B2uxx6, J2uxx6;
wire R2uxx6, Z2uxx6, H3uxx6, P3uxx6, X3uxx6, F4uxx6, N4uxx6, V4uxx6, D5uxx6, L5uxx6;
wire T5uxx6, B6uxx6, J6uxx6, R6uxx6, Z6uxx6, H7uxx6, P7uxx6, X7uxx6, F8uxx6, N8uxx6;
wire V8uxx6, D9uxx6, L9uxx6, T9uxx6, Bauxx6, Jauxx6, Rauxx6, Zauxx6, Hbuxx6, Pbuxx6;
wire Xbuxx6, Fcuxx6, Ncuxx6, Vcuxx6, Dduxx6, Lduxx6, Tduxx6, Beuxx6, Jeuxx6, Reuxx6;
wire Zeuxx6, Hfuxx6, Pfuxx6, Xfuxx6, Fguxx6, Nguxx6, Vguxx6, Dhuxx6, Lhuxx6, Thuxx6;
wire Biuxx6, Jiuxx6, Riuxx6, Ziuxx6, Hjuxx6, Pjuxx6, Xjuxx6, Fkuxx6, Nkuxx6, Vkuxx6;
wire Dluxx6, Lluxx6, Tluxx6, Bmuxx6, Jmuxx6, Rmuxx6, Zmuxx6, Hnuxx6, Pnuxx6, Xnuxx6;
wire Fouxx6, Nouxx6, Vouxx6, Dpuxx6, Lpuxx6, Tpuxx6, Bquxx6, Jquxx6, Rquxx6, Zquxx6;
wire Hruxx6, Pruxx6, Xruxx6, Fsuxx6, Nsuxx6, Vsuxx6, Dtuxx6, Ltuxx6, Ttuxx6, Buuxx6;
wire Juuxx6, Ruuxx6, Zuuxx6, Hvuxx6, Pvuxx6, Xvuxx6, Fwuxx6, Nwuxx6, Vwuxx6, Dxuxx6;
wire Lxuxx6, Txuxx6, Byuxx6, Jyuxx6, Ryuxx6, Zyuxx6, Hzuxx6, Pzuxx6, Xzuxx6, F0vxx6;
wire N0vxx6, V0vxx6, D1vxx6, L1vxx6, T1vxx6, B2vxx6, J2vxx6, R2vxx6, Z2vxx6, H3vxx6;
wire P3vxx6, X3vxx6, F4vxx6, N4vxx6, V4vxx6, D5vxx6, L5vxx6, T5vxx6, B6vxx6, J6vxx6;
wire R6vxx6, Z6vxx6, H7vxx6, P7vxx6, X7vxx6, F8vxx6, N8vxx6, V8vxx6, D9vxx6, L9vxx6;
wire T9vxx6, Bavxx6, Javxx6, Ravxx6, Zavxx6, Hbvxx6, Pbvxx6, Xbvxx6, Fcvxx6, Ncvxx6;
wire Vcvxx6, Ddvxx6, Ldvxx6, Tdvxx6, Bevxx6, Jevxx6, Revxx6, Zevxx6, Hfvxx6, Pfvxx6;
wire Xfvxx6, Fgvxx6, Ngvxx6, Vgvxx6, Dhvxx6, Lhvxx6, Thvxx6, Bivxx6, Jivxx6, Rivxx6;
wire Zivxx6, Hjvxx6, Pjvxx6, Xjvxx6, Fkvxx6, Nkvxx6, Vkvxx6, Dlvxx6, Llvxx6, Tlvxx6;
wire Bmvxx6, Jmvxx6, Rmvxx6, Zmvxx6, Hnvxx6, Pnvxx6, Xnvxx6, Fovxx6, Novxx6, Vovxx6;
wire Dpvxx6, Lpvxx6, Tpvxx6, Bqvxx6, Jqvxx6, Rqvxx6, Zqvxx6, Hrvxx6, Prvxx6, Xrvxx6;
wire Fsvxx6, Nsvxx6, Vsvxx6, Dtvxx6, Ltvxx6, Ttvxx6, Buvxx6, Juvxx6, Ruvxx6, Zuvxx6;
wire Hvvxx6, Pvvxx6, Xvvxx6, Fwvxx6, Nwvxx6, Vwvxx6, Dxvxx6, Lxvxx6, Txvxx6, Byvxx6;
wire Jyvxx6, Ryvxx6, Zyvxx6, Hzvxx6, Pzvxx6, Xzvxx6, F0wxx6, N0wxx6, V0wxx6, D1wxx6;
wire L1wxx6, T1wxx6, B2wxx6, J2wxx6, R2wxx6, Z2wxx6, H3wxx6, P3wxx6, X3wxx6, F4wxx6;
wire N4wxx6, V4wxx6, D5wxx6, L5wxx6, T5wxx6, B6wxx6, J6wxx6, R6wxx6, Z6wxx6, H7wxx6;
wire P7wxx6, X7wxx6, F8wxx6, N8wxx6, V8wxx6, D9wxx6, L9wxx6, T9wxx6, Bawxx6, Jawxx6;
wire Rawxx6, Zawxx6, Hbwxx6, Pbwxx6, Xbwxx6, Fcwxx6, Ncwxx6, Vcwxx6, Ddwxx6, Ldwxx6;
wire Tdwxx6, Bewxx6, Jewxx6, Rewxx6, Zewxx6, Hfwxx6, Pfwxx6, Xfwxx6, Fgwxx6, Ngwxx6;
wire Vgwxx6, Dhwxx6, Lhwxx6, Thwxx6, Biwxx6, Jiwxx6, Riwxx6, Ziwxx6, Hjwxx6, Pjwxx6;
wire Xjwxx6, Fkwxx6, Nkwxx6, Vkwxx6, Dlwxx6, Llwxx6, Tlwxx6, Bmwxx6, Jmwxx6, Rmwxx6;
wire Zmwxx6, Hnwxx6, Pnwxx6, Xnwxx6, Fowxx6, Nowxx6, Vowxx6, Dpwxx6, Lpwxx6, Tpwxx6;
wire Bqwxx6, Jqwxx6, Rqwxx6, Zqwxx6, Hrwxx6, Prwxx6, Xrwxx6, Fswxx6, Nswxx6, Vswxx6;
wire Dtwxx6, Ltwxx6, Ttwxx6, Buwxx6, Juwxx6, Ruwxx6, Zuwxx6, Hvwxx6, Pvwxx6, Xvwxx6;
wire Fwwxx6, Nwwxx6, Vwwxx6, Dxwxx6, Lxwxx6, Txwxx6, Bywxx6, Jywxx6, Rywxx6, Zywxx6;
wire Hzwxx6, Pzwxx6, Xzwxx6, F0xxx6, N0xxx6, V0xxx6, D1xxx6, L1xxx6, T1xxx6, B2xxx6;
wire J2xxx6, R2xxx6, Z2xxx6, H3xxx6, P3xxx6, X3xxx6, F4xxx6, N4xxx6, V4xxx6, D5xxx6;
wire L5xxx6, T5xxx6, B6xxx6, J6xxx6, R6xxx6, Z6xxx6, H7xxx6, P7xxx6, X7xxx6, F8xxx6;
wire N8xxx6, V8xxx6, D9xxx6, L9xxx6, T9xxx6, Baxxx6, Jaxxx6, Raxxx6, Zaxxx6, Hbxxx6;
wire Pbxxx6, Xbxxx6, Fcxxx6, Ncxxx6, Vcxxx6, Ddxxx6, Ldxxx6, Tdxxx6, Bexxx6, Jexxx6;
wire Rexxx6, Zexxx6, Hfxxx6, Pfxxx6, Xfxxx6, Fgxxx6, Ngxxx6, Vgxxx6, Dhxxx6, Lhxxx6;
wire Thxxx6, Bixxx6, Jixxx6, Rixxx6, Zixxx6, Hjxxx6, Pjxxx6, Xjxxx6, Fkxxx6, Nkxxx6;
wire Vkxxx6, Dlxxx6, Llxxx6, Tlxxx6, Bmxxx6, Jmxxx6, Rmxxx6, Zmxxx6, Hnxxx6, Pnxxx6;
wire Xnxxx6, Foxxx6, Noxxx6, Voxxx6, Dpxxx6, Lpxxx6, Tpxxx6, Bqxxx6, Jqxxx6, Rqxxx6;
wire Zqxxx6, Hrxxx6, Prxxx6, Xrxxx6, Fsxxx6, Nsxxx6, Vsxxx6, Dtxxx6, Ltxxx6, Ttxxx6;
wire Buxxx6, Juxxx6, Ruxxx6, Zuxxx6, Hvxxx6, Pvxxx6, Xvxxx6, Fwxxx6, Nwxxx6, Vwxxx6;
wire Dxxxx6, Lxxxx6, Txxxx6, Byxxx6, Jyxxx6, Ryxxx6, Zyxxx6, Hzxxx6, Pzxxx6, Xzxxx6;
wire F0yxx6, N0yxx6, V0yxx6, D1yxx6, L1yxx6, T1yxx6, B2yxx6, J2yxx6, R2yxx6, Z2yxx6;
wire H3yxx6, P3yxx6, X3yxx6, F4yxx6, N4yxx6, V4yxx6, D5yxx6, L5yxx6, T5yxx6, B6yxx6;
wire J6yxx6, R6yxx6, Z6yxx6, H7yxx6, P7yxx6, X7yxx6, F8yxx6, N8yxx6, V8yxx6, D9yxx6;
wire L9yxx6, T9yxx6, Bayxx6, Jayxx6, Rayxx6, Zayxx6, Hbyxx6, Pbyxx6, Xbyxx6, Fcyxx6;
wire Ncyxx6, Vcyxx6, Ddyxx6, Ldyxx6, Tdyxx6, Beyxx6, Jeyxx6, Reyxx6, Zeyxx6, Hfyxx6;
wire Pfyxx6, Xfyxx6, Fgyxx6, Ngyxx6, Vgyxx6, Dhyxx6, Lhyxx6, Thyxx6, Biyxx6, Jiyxx6;
wire Riyxx6, Ziyxx6, Hjyxx6, Pjyxx6, Xjyxx6, Fkyxx6, Nkyxx6, Vkyxx6, Dlyxx6, Llyxx6;
wire Tlyxx6, Bmyxx6, Jmyxx6, Rmyxx6, Zmyxx6, Hnyxx6, Pnyxx6, Xnyxx6, Foyxx6, Noyxx6;
wire Voyxx6, Dpyxx6, Lpyxx6, Tpyxx6, Bqyxx6, Jqyxx6, Rqyxx6, Zqyxx6, Hryxx6, Pryxx6;
wire Xryxx6, Fsyxx6, Nsyxx6, Vsyxx6, Dtyxx6, Ltyxx6, Ttyxx6, Buyxx6, Juyxx6, Ruyxx6;
wire Zuyxx6, Hvyxx6, Pvyxx6, Xvyxx6, Fwyxx6, Nwyxx6, Vwyxx6, Dxyxx6, Lxyxx6, Txyxx6;
wire Byyxx6, Jyyxx6, Ryyxx6, Zyyxx6, Hzyxx6, Pzyxx6, Xzyxx6, F0zxx6, N0zxx6, V0zxx6;
wire D1zxx6, L1zxx6, T1zxx6, B2zxx6, J2zxx6, R2zxx6, Z2zxx6, H3zxx6, P3zxx6, X3zxx6;
wire F4zxx6, N4zxx6, V4zxx6, D5zxx6, L5zxx6, T5zxx6, B6zxx6, J6zxx6, R6zxx6, Z6zxx6;
wire H7zxx6, P7zxx6, X7zxx6, F8zxx6, N8zxx6, V8zxx6, D9zxx6, L9zxx6, T9zxx6, Bazxx6;
wire Jazxx6, Razxx6, Zazxx6, Hbzxx6, Pbzxx6, Xbzxx6, Fczxx6, Nczxx6, Vczxx6, Ddzxx6;
wire Ldzxx6, Tdzxx6, Bezxx6, Jezxx6, Rezxx6, Zezxx6, Hfzxx6, Pfzxx6, Xfzxx6, Fgzxx6;
wire Ngzxx6, Vgzxx6, Dhzxx6, Lhzxx6, Thzxx6, Bizxx6, Jizxx6, Rizxx6, Zizxx6, Hjzxx6;
wire Pjzxx6, Xjzxx6, Fkzxx6, Nkzxx6, Vkzxx6, Dlzxx6, Llzxx6, Tlzxx6, Bmzxx6, Jmzxx6;
wire Rmzxx6, Zmzxx6, Hnzxx6, Pnzxx6, Xnzxx6, Fozxx6, Nozxx6, Vozxx6, Dpzxx6, Lpzxx6;
wire Tpzxx6, Bqzxx6, Jqzxx6, Rqzxx6, Zqzxx6, Hrzxx6, Przxx6, Xrzxx6, Fszxx6, Nszxx6;
wire Vszxx6, Dtzxx6, Ltzxx6, Ttzxx6, Buzxx6, Juzxx6, Ruzxx6, Zuzxx6, Hvzxx6, Pvzxx6;
wire Xvzxx6, Fwzxx6, Nwzxx6, Vwzxx6, Dxzxx6, Lxzxx6, Txzxx6, Byzxx6, Jyzxx6, Ryzxx6;
wire Zyzxx6, Hzzxx6, Pzzxx6, Xzzxx6, F00yx6, N00yx6, V00yx6, D10yx6, L10yx6, T10yx6;
wire B20yx6, J20yx6, R20yx6, Z20yx6, H30yx6, P30yx6, X30yx6, F40yx6, N40yx6, V40yx6;
wire D50yx6, L50yx6, T50yx6, B60yx6, J60yx6, R60yx6, Z60yx6, H70yx6, P70yx6, X70yx6;
wire F80yx6, N80yx6, V80yx6, D90yx6, L90yx6, T90yx6, Ba0yx6, Ja0yx6, Ra0yx6, Za0yx6;
wire Hb0yx6, Pb0yx6, Xb0yx6, Fc0yx6, Nc0yx6, Vc0yx6, Dd0yx6, Ld0yx6, Td0yx6, Be0yx6;
wire Je0yx6, Re0yx6, Ze0yx6, Hf0yx6, Pf0yx6, Xf0yx6, Fg0yx6, Ng0yx6, Vg0yx6, Dh0yx6;
wire Lh0yx6, Th0yx6, Bi0yx6, Ji0yx6, Ri0yx6, Zi0yx6, Hj0yx6, Pj0yx6, Xj0yx6, Fk0yx6;
wire Nk0yx6, Vk0yx6, Dl0yx6, Ll0yx6, Tl0yx6, Bm0yx6, Jm0yx6, Rm0yx6, Zm0yx6, Hn0yx6;
wire Pn0yx6, Xn0yx6, Fo0yx6, No0yx6, Vo0yx6, Dp0yx6, Lp0yx6, Tp0yx6, Bq0yx6, Jq0yx6;
wire Rq0yx6, Zq0yx6, Hr0yx6, Pr0yx6, Xr0yx6, Fs0yx6, Ns0yx6, Vs0yx6, Dt0yx6, Lt0yx6;
wire Tt0yx6, Bu0yx6, Ju0yx6, Ru0yx6, Zu0yx6, Hv0yx6, Pv0yx6, Xv0yx6, Fw0yx6, Nw0yx6;
wire Vw0yx6, Dx0yx6, Lx0yx6, Tx0yx6, By0yx6, Jy0yx6, Ry0yx6, Zy0yx6, Hz0yx6, Pz0yx6;
wire Xz0yx6, F01yx6, N01yx6, V01yx6, D11yx6, L11yx6, T11yx6, B21yx6, J21yx6, R21yx6;
wire Z21yx6, H31yx6, P31yx6, X31yx6, F41yx6, N41yx6, V41yx6, D51yx6, L51yx6, T51yx6;
wire B61yx6, J61yx6, R61yx6, Z61yx6, H71yx6, P71yx6, X71yx6, F81yx6, N81yx6, V81yx6;
wire D91yx6, L91yx6, T91yx6, Ba1yx6, Ja1yx6, Ra1yx6, Za1yx6, Hb1yx6, Pb1yx6, Xb1yx6;
wire Fc1yx6, Nc1yx6, Vc1yx6, Dd1yx6, Ld1yx6, Td1yx6, Be1yx6, Je1yx6, Re1yx6, Ze1yx6;
wire Hf1yx6, Pf1yx6, Xf1yx6, Fg1yx6, Ng1yx6, Vg1yx6, Dh1yx6, Lh1yx6, Th1yx6, Bi1yx6;
wire Ji1yx6, Ri1yx6, Zi1yx6, Hj1yx6, Pj1yx6, Xj1yx6, Fk1yx6, Nk1yx6, Vk1yx6, Dl1yx6;
wire Ll1yx6, Tl1yx6, Bm1yx6, Jm1yx6, Rm1yx6, Zm1yx6, Hn1yx6, Pn1yx6, Xn1yx6, Fo1yx6;
wire No1yx6, Vo1yx6, Dp1yx6, Lp1yx6, Tp1yx6, Bq1yx6, Jq1yx6, Rq1yx6, Zq1yx6, Hr1yx6;
wire Pr1yx6, Xr1yx6, Fs1yx6, Ns1yx6, Vs1yx6, Dt1yx6, Lt1yx6, Tt1yx6, Bu1yx6, Ju1yx6;
wire Ru1yx6, Zu1yx6, Hv1yx6, Pv1yx6, Xv1yx6, Fw1yx6, Nw1yx6, Vw1yx6, Dx1yx6, Lx1yx6;
wire Tx1yx6, By1yx6, Jy1yx6, Ry1yx6, Zy1yx6, Hz1yx6, Pz1yx6, Xz1yx6, F02yx6, N02yx6;
wire V02yx6, D12yx6, L12yx6, T12yx6, B22yx6, J22yx6, R22yx6, Z22yx6, H32yx6, P32yx6;
wire X32yx6, F42yx6, N42yx6, V42yx6, D52yx6, L52yx6, T52yx6, B62yx6, J62yx6, R62yx6;
wire Z62yx6, H72yx6, P72yx6, X72yx6, F82yx6, N82yx6, V82yx6, D92yx6, L92yx6, T92yx6;
wire Ba2yx6, Ja2yx6, Ra2yx6, Za2yx6, Hb2yx6, Pb2yx6, Xb2yx6, Fc2yx6, Nc2yx6, Vc2yx6;
wire Dd2yx6, Ld2yx6, Td2yx6, Be2yx6, Je2yx6, Re2yx6, Ze2yx6, Hf2yx6, Pf2yx6, Xf2yx6;
wire Fg2yx6, Ng2yx6, Vg2yx6, Dh2yx6, Lh2yx6, Th2yx6, Bi2yx6, Ji2yx6, Ri2yx6, Zi2yx6;
wire Hj2yx6, Pj2yx6, Xj2yx6, Fk2yx6, Nk2yx6, Vk2yx6, Dl2yx6, Ll2yx6, Tl2yx6, Bm2yx6;
wire Jm2yx6, Rm2yx6, Zm2yx6, Hn2yx6, Pn2yx6, Xn2yx6, Fo2yx6, No2yx6, Vo2yx6, Dp2yx6;
wire Lp2yx6, Tp2yx6, Bq2yx6, Jq2yx6, Rq2yx6, Zq2yx6, Hr2yx6, Pr2yx6, Xr2yx6, Fs2yx6;
wire Ns2yx6, Vs2yx6, Dt2yx6, Lt2yx6, Tt2yx6, Bu2yx6, Ju2yx6, Ru2yx6, Zu2yx6, Hv2yx6;
wire Pv2yx6, Xv2yx6, Fw2yx6, Nw2yx6, Vw2yx6, Dx2yx6, Lx2yx6, Tx2yx6, By2yx6, Jy2yx6;
wire Ry2yx6, Zy2yx6, Hz2yx6, Pz2yx6, Xz2yx6, F03yx6, N03yx6, V03yx6, D13yx6, L13yx6;
wire T13yx6, B23yx6, J23yx6, R23yx6, Z23yx6, H33yx6, P33yx6, X33yx6, F43yx6, N43yx6;
wire V43yx6, D53yx6, L53yx6, T53yx6, B63yx6, J63yx6, R63yx6, Z63yx6, H73yx6, P73yx6;
wire X73yx6, F83yx6, N83yx6, V83yx6, D93yx6, L93yx6, T93yx6, Ba3yx6, Ja3yx6, Ra3yx6;
wire Za3yx6, Hb3yx6, Pb3yx6, Xb3yx6, Fc3yx6, Nc3yx6, Vc3yx6, Dd3yx6, Ld3yx6, Td3yx6;
wire Be3yx6, Je3yx6, Re3yx6, Ze3yx6, Hf3yx6, Pf3yx6, Xf3yx6, Fg3yx6, Ng3yx6, Vg3yx6;
wire Dh3yx6, Lh3yx6, Th3yx6, Bi3yx6, Ji3yx6, Ri3yx6, Zi3yx6, Hj3yx6, Pj3yx6, Xj3yx6;
wire Fk3yx6, Nk3yx6, Vk3yx6, Dl3yx6, Ll3yx6, Tl3yx6, Bm3yx6, Jm3yx6, Rm3yx6, Zm3yx6;
wire Hn3yx6, Pn3yx6, Xn3yx6, Fo3yx6, No3yx6, Vo3yx6, Dp3yx6, Lp3yx6, Tp3yx6, Bq3yx6;
wire Jq3yx6, Rq3yx6, Zq3yx6, Hr3yx6, Pr3yx6, Xr3yx6, Fs3yx6, Ns3yx6, Vs3yx6, Dt3yx6;
wire Lt3yx6, Tt3yx6, Bu3yx6, Ju3yx6, Ru3yx6, Zu3yx6, Hv3yx6, Pv3yx6, Xv3yx6, Fw3yx6;
wire Nw3yx6, Vw3yx6, Dx3yx6, Lx3yx6, Tx3yx6, By3yx6, Jy3yx6, Ry3yx6, Zy3yx6, Hz3yx6;
wire Pz3yx6, Xz3yx6, F04yx6, N04yx6, V04yx6, D14yx6, L14yx6, T14yx6, B24yx6, J24yx6;
wire R24yx6, Z24yx6, H34yx6, P34yx6, X34yx6, F44yx6, N44yx6, V44yx6, D54yx6, L54yx6;
wire T54yx6, B64yx6, J64yx6, R64yx6, Z64yx6, H74yx6, P74yx6, X74yx6, F84yx6, N84yx6;
wire V84yx6, D94yx6, L94yx6, T94yx6, Ba4yx6, Ja4yx6, Ra4yx6, Za4yx6, Hb4yx6, Pb4yx6;
wire Xb4yx6, Fc4yx6, Nc4yx6, Vc4yx6, Dd4yx6, Ld4yx6, Td4yx6, Be4yx6, Je4yx6, Re4yx6;
wire Ze4yx6, Hf4yx6, Pf4yx6, Xf4yx6, Fg4yx6, Ng4yx6, Vg4yx6, Dh4yx6, Lh4yx6, Th4yx6;
wire Bi4yx6, Ji4yx6, Ri4yx6, Zi4yx6, Hj4yx6, Pj4yx6, Xj4yx6, Fk4yx6, Nk4yx6, Vk4yx6;
wire Dl4yx6, Ll4yx6, Tl4yx6, Bm4yx6, Jm4yx6, Rm4yx6, Zm4yx6, Hn4yx6, Pn4yx6, Xn4yx6;
wire Fo4yx6, No4yx6, Vo4yx6, Dp4yx6, Lp4yx6, Tp4yx6, Bq4yx6, Jq4yx6, Rq4yx6, Zq4yx6;
wire Hr4yx6, Pr4yx6, Xr4yx6, Fs4yx6, Ns4yx6, Vs4yx6, Dt4yx6, Lt4yx6, Tt4yx6, Bu4yx6;
wire Ju4yx6, Ru4yx6, Zu4yx6, Hv4yx6, Pv4yx6, Xv4yx6, Fw4yx6, Nw4yx6, Vw4yx6, Dx4yx6;
wire Lx4yx6, Tx4yx6, By4yx6, Jy4yx6, Ry4yx6, Zy4yx6, Hz4yx6, Pz4yx6, Xz4yx6, F05yx6;
wire N05yx6, V05yx6, D15yx6, L15yx6, T15yx6, B25yx6, J25yx6, R25yx6, Z25yx6, H35yx6;
wire P35yx6, X35yx6, F45yx6, N45yx6, V45yx6, D55yx6, L55yx6, T55yx6, B65yx6, J65yx6;
wire R65yx6, Z65yx6, H75yx6, P75yx6, X75yx6, F85yx6, N85yx6, V85yx6, D95yx6, L95yx6;
wire T95yx6, Ba5yx6, Ja5yx6, Ra5yx6, Za5yx6, Hb5yx6, Pb5yx6, Xb5yx6, Fc5yx6, Nc5yx6;
wire Vc5yx6, Dd5yx6, Ld5yx6, Td5yx6, Be5yx6, Je5yx6, Re5yx6, Ze5yx6, Hf5yx6, Pf5yx6;
wire Xf5yx6, Fg5yx6, Ng5yx6, Vg5yx6, Dh5yx6, Lh5yx6, Th5yx6, Bi5yx6, Ji5yx6, Ri5yx6;
wire Zi5yx6, Hj5yx6, Pj5yx6, Xj5yx6, Fk5yx6, Nk5yx6, Vk5yx6, Dl5yx6, Ll5yx6, Tl5yx6;
wire Bm5yx6, Jm5yx6, Rm5yx6, Zm5yx6, Hn5yx6, Pn5yx6, Xn5yx6, Fo5yx6, No5yx6, Vo5yx6;
wire Dp5yx6, Lp5yx6, Tp5yx6, Bq5yx6, Jq5yx6, Rq5yx6, Zq5yx6, Hr5yx6, Pr5yx6, Xr5yx6;
wire Fs5yx6, Ns5yx6, Vs5yx6, Dt5yx6, Lt5yx6, Tt5yx6, Bu5yx6, Ju5yx6, Ru5yx6, Zu5yx6;
wire Hv5yx6, Pv5yx6, Xv5yx6, Fw5yx6, Nw5yx6, Vw5yx6, Dx5yx6, Lx5yx6, Tx5yx6, By5yx6;
wire Jy5yx6, Ry5yx6, Zy5yx6, Hz5yx6, Pz5yx6, Xz5yx6, F06yx6, N06yx6, V06yx6, D16yx6;
wire L16yx6, T16yx6, B26yx6, J26yx6, R26yx6, Z26yx6, H36yx6, P36yx6, X36yx6, F46yx6;
wire N46yx6, V46yx6, D56yx6, L56yx6, T56yx6, B66yx6, J66yx6, R66yx6, Z66yx6, H76yx6;
wire P76yx6, X76yx6, F86yx6, N86yx6, V86yx6, D96yx6, L96yx6, T96yx6, Ba6yx6, Ja6yx6;
wire Ra6yx6, Za6yx6, Hb6yx6, Pb6yx6, Xb6yx6, Fc6yx6, Nc6yx6, Vc6yx6, Dd6yx6, Ld6yx6;
wire Td6yx6, Be6yx6, Je6yx6, Re6yx6, Ze6yx6, Hf6yx6, Pf6yx6, Xf6yx6, Fg6yx6, Ng6yx6;
wire Vg6yx6, Dh6yx6, Lh6yx6, Th6yx6, Bi6yx6, Ji6yx6, Ri6yx6, Zi6yx6, Hj6yx6, Pj6yx6;
wire Xj6yx6, Fk6yx6, Nk6yx6, Vk6yx6, Dl6yx6, Ll6yx6, Tl6yx6, Bm6yx6, Jm6yx6, Rm6yx6;
wire Zm6yx6, Hn6yx6, Pn6yx6, Xn6yx6, Fo6yx6, No6yx6, Vo6yx6, Dp6yx6, Lp6yx6, Tp6yx6;
wire Bq6yx6, Jq6yx6, Rq6yx6, Zq6yx6, Hr6yx6, Pr6yx6, Xr6yx6, Fs6yx6, Ns6yx6, Vs6yx6;
wire Dt6yx6, Lt6yx6, Tt6yx6, Bu6yx6, Ju6yx6, Ru6yx6, Zu6yx6, Hv6yx6, Pv6yx6, Xv6yx6;
wire Fw6yx6, Nw6yx6, Vw6yx6, Dx6yx6, Lx6yx6, Tx6yx6, By6yx6, Jy6yx6, Ry6yx6, Zy6yx6;
wire Hz6yx6, Pz6yx6, Xz6yx6, F07yx6, N07yx6, V07yx6, D17yx6, L17yx6, T17yx6, B27yx6;
wire J27yx6, R27yx6, Z27yx6, H37yx6, P37yx6, X37yx6, F47yx6, N47yx6, V47yx6, D57yx6;
wire L57yx6, T57yx6, B67yx6, J67yx6, R67yx6, Z67yx6, H77yx6, P77yx6, X77yx6, F87yx6;
wire N87yx6, V87yx6, D97yx6, L97yx6, T97yx6, Ba7yx6, Ja7yx6, Ra7yx6, Za7yx6, Hb7yx6;
wire Pb7yx6, Xb7yx6, Fc7yx6, Nc7yx6, Vc7yx6, Dd7yx6, Ld7yx6, Td7yx6, Be7yx6, Je7yx6;
wire Re7yx6, Ze7yx6, Hf7yx6, Pf7yx6, Xf7yx6, Fg7yx6, Ng7yx6, Vg7yx6, Dh7yx6, Lh7yx6;
wire Th7yx6, Bi7yx6, Ji7yx6, Ri7yx6, Zi7yx6, Hj7yx6, Pj7yx6, Xj7yx6, Fk7yx6, Nk7yx6;
wire Vk7yx6, Dl7yx6, Ll7yx6, Tl7yx6, Bm7yx6, Jm7yx6, Rm7yx6, Zm7yx6, Hn7yx6, Pn7yx6;
wire Xn7yx6, Fo7yx6, No7yx6, Vo7yx6, Dp7yx6, Lp7yx6, Tp7yx6, Bq7yx6, Jq7yx6, Rq7yx6;
wire Zq7yx6, Hr7yx6, Pr7yx6, Xr7yx6, Fs7yx6, Ns7yx6, Vs7yx6, Dt7yx6, Lt7yx6, Tt7yx6;
wire Bu7yx6, Ju7yx6, Ru7yx6, Zu7yx6, Hv7yx6, Pv7yx6, Xv7yx6, Fw7yx6, Nw7yx6, Vw7yx6;
wire Dx7yx6, Lx7yx6, Tx7yx6, By7yx6, Jy7yx6, Ry7yx6, Zy7yx6, Hz7yx6, Pz7yx6, Xz7yx6;
wire F08yx6, N08yx6, V08yx6, D18yx6, L18yx6, T18yx6, B28yx6, J28yx6, R28yx6, Z28yx6;
wire H38yx6, P38yx6, X38yx6, F48yx6, N48yx6, V48yx6, D58yx6, L58yx6, T58yx6, B68yx6;
wire J68yx6, R68yx6, Z68yx6, H78yx6, P78yx6, X78yx6, F88yx6, N88yx6, V88yx6, D98yx6;
wire L98yx6, T98yx6, Ba8yx6, Ja8yx6, Ra8yx6, Za8yx6, Hb8yx6, Pb8yx6, Xb8yx6, Fc8yx6;
wire Nc8yx6, Vc8yx6, Dd8yx6, Ld8yx6, Td8yx6, Be8yx6, Je8yx6, Re8yx6, Ze8yx6, Hf8yx6;
wire Pf8yx6, Xf8yx6, Fg8yx6, Ng8yx6, Vg8yx6, Dh8yx6, Lh8yx6, Th8yx6, Bi8yx6, Ji8yx6;
wire Ri8yx6, Zi8yx6, Hj8yx6, Pj8yx6, Xj8yx6, Fk8yx6, Nk8yx6, Vk8yx6, Dl8yx6, Ll8yx6;
wire Tl8yx6, Bm8yx6, Jm8yx6, Rm8yx6, Zm8yx6, Hn8yx6, Pn8yx6, Xn8yx6, Fo8yx6, No8yx6;
wire Vo8yx6, Dp8yx6, Lp8yx6, Tp8yx6, Bq8yx6, Jq8yx6, Rq8yx6, Zq8yx6, Hr8yx6, Pr8yx6;
wire Xr8yx6, Fs8yx6, Ns8yx6, Vs8yx6, Dt8yx6, Lt8yx6, Tt8yx6, Bu8yx6, Ju8yx6, Ru8yx6;
wire Zu8yx6, Hv8yx6, Pv8yx6, Xv8yx6, Fw8yx6, Nw8yx6, Vw8yx6, Dx8yx6, Lx8yx6, Tx8yx6;
wire By8yx6, Jy8yx6, Ry8yx6, Zy8yx6, Hz8yx6, Pz8yx6, Xz8yx6, F09yx6, N09yx6, V09yx6;
wire D19yx6, L19yx6, T19yx6, B29yx6, J29yx6, R29yx6, Z29yx6, H39yx6, P39yx6, X39yx6;
wire F49yx6, N49yx6, V49yx6, D59yx6, L59yx6, T59yx6, B69yx6, J69yx6, R69yx6, Z69yx6;
wire H79yx6, P79yx6, X79yx6, F89yx6, N89yx6, V89yx6, D99yx6, L99yx6, T99yx6, Ba9yx6;
wire Ja9yx6, Ra9yx6, Za9yx6, Hb9yx6, Pb9yx6, Xb9yx6, Fc9yx6, Nc9yx6, Vc9yx6, Dd9yx6;
wire Ld9yx6, Td9yx6, Be9yx6, Je9yx6, Re9yx6, Ze9yx6, Hf9yx6, Pf9yx6, Xf9yx6, Fg9yx6;
wire Ng9yx6, Vg9yx6, Dh9yx6, Lh9yx6, Th9yx6, Bi9yx6, Ji9yx6, Ri9yx6, Zi9yx6, Hj9yx6;
wire Pj9yx6, Xj9yx6, Fk9yx6, Nk9yx6, Vk9yx6, Dl9yx6, Ll9yx6, Tl9yx6, Bm9yx6, Jm9yx6;
wire Rm9yx6, Zm9yx6, Hn9yx6, Pn9yx6, Xn9yx6, Fo9yx6, No9yx6, Vo9yx6, Dp9yx6, Lp9yx6;
wire Tp9yx6, Bq9yx6, Jq9yx6, Rq9yx6, Zq9yx6, Hr9yx6, Pr9yx6, Xr9yx6, Fs9yx6, Ns9yx6;
wire Vs9yx6, Dt9yx6, Lt9yx6, Tt9yx6, Bu9yx6, Ju9yx6, Ru9yx6, Zu9yx6, Hv9yx6, Pv9yx6;
wire Xv9yx6, Fw9yx6, Nw9yx6, Vw9yx6, Dx9yx6, Lx9yx6, Tx9yx6, By9yx6, Jy9yx6, Ry9yx6;
wire Zy9yx6, Hz9yx6, Pz9yx6, Xz9yx6, F0ayx6, N0ayx6, V0ayx6, D1ayx6, L1ayx6, T1ayx6;
wire B2ayx6, J2ayx6, R2ayx6, Z2ayx6, H3ayx6, P3ayx6, X3ayx6, F4ayx6, N4ayx6, V4ayx6;
wire D5ayx6, L5ayx6, T5ayx6, B6ayx6, J6ayx6, R6ayx6, Z6ayx6, H7ayx6, P7ayx6, X7ayx6;
wire F8ayx6, N8ayx6, V8ayx6, D9ayx6, L9ayx6, T9ayx6, Baayx6, Jaayx6, Raayx6, Zaayx6;
wire Hbayx6, Pbayx6, Xbayx6, Fcayx6, Ncayx6, Vcayx6, Ddayx6, Ldayx6, Tdayx6, Beayx6;
wire Jeayx6, Reayx6, Zeayx6, Hfayx6, Pfayx6, Xfayx6, Fgayx6, Ngayx6, Vgayx6, Dhayx6;
wire Lhayx6, Thayx6, Biayx6, Jiayx6, Riayx6, Ziayx6, Hjayx6, Pjayx6, Xjayx6, Fkayx6;
wire Nkayx6, Vkayx6, Dlayx6, Llayx6, Tlayx6, Bmayx6, Jmayx6, Rmayx6, Zmayx6, Hnayx6;
wire Pnayx6, Xnayx6, Foayx6, Noayx6, Voayx6, Dpayx6, Lpayx6, Tpayx6, Bqayx6, Jqayx6;
wire Rqayx6, Zqayx6, Hrayx6, Prayx6, Xrayx6, Fsayx6, Nsayx6, Vsayx6, Dtayx6, Ltayx6;
wire Ttayx6, Buayx6, Juayx6, Ruayx6, Zuayx6, Hvayx6, Pvayx6, Xvayx6, Fwayx6, Nwayx6;
wire Vwayx6, Dxayx6, Lxayx6, Txayx6, Byayx6, Jyayx6, Ryayx6, Zyayx6, Hzayx6, Pzayx6;
wire Xzayx6, F0byx6, N0byx6, V0byx6, D1byx6, L1byx6, T1byx6, B2byx6, J2byx6, R2byx6;
wire Z2byx6, H3byx6, P3byx6, X3byx6, F4byx6, N4byx6, V4byx6, D5byx6, L5byx6, T5byx6;
wire B6byx6, J6byx6, R6byx6, Z6byx6, H7byx6, P7byx6, X7byx6, F8byx6, N8byx6, V8byx6;
wire D9byx6, L9byx6, T9byx6, Babyx6, Jabyx6, Rabyx6, Zabyx6, Hbbyx6, Pbbyx6, Xbbyx6;
wire Fcbyx6, Ncbyx6, Vcbyx6, Ddbyx6, Ldbyx6, Tdbyx6, Bebyx6, Jebyx6, Rebyx6, Zebyx6;
wire Hfbyx6, Pfbyx6, Xfbyx6, Fgbyx6, Ngbyx6, Vgbyx6, Dhbyx6, Lhbyx6, Thbyx6, Bibyx6;
wire Jibyx6, Ribyx6, Zibyx6, Hjbyx6, Pjbyx6, Xjbyx6, Fkbyx6, Nkbyx6, Vkbyx6, Dlbyx6;
wire Llbyx6, Tlbyx6, Bmbyx6, Jmbyx6, Rmbyx6, Zmbyx6, Hnbyx6, Pnbyx6, Xnbyx6, Fobyx6;
wire Nobyx6, Vobyx6, Dpbyx6, Lpbyx6, Tpbyx6, Bqbyx6, Jqbyx6, Rqbyx6, Zqbyx6, Hrbyx6;
wire Prbyx6, Xrbyx6, Fsbyx6, Nsbyx6, Vsbyx6, Dtbyx6, Ltbyx6, Ttbyx6, Bubyx6, Jubyx6;
wire Rubyx6, Zubyx6, Hvbyx6, Pvbyx6, Xvbyx6, Fwbyx6, Nwbyx6, Vwbyx6, Dxbyx6, Lxbyx6;
wire Txbyx6, Bybyx6, Jybyx6, Rybyx6, Zybyx6, Hzbyx6, Pzbyx6, Xzbyx6, F0cyx6, N0cyx6;
wire V0cyx6, D1cyx6, L1cyx6, T1cyx6, B2cyx6, J2cyx6, R2cyx6, Z2cyx6, H3cyx6, P3cyx6;
wire X3cyx6, F4cyx6, N4cyx6, V4cyx6, D5cyx6, L5cyx6, T5cyx6, B6cyx6, J6cyx6, R6cyx6;
wire Z6cyx6, H7cyx6, P7cyx6, X7cyx6, F8cyx6, N8cyx6, V8cyx6, D9cyx6, L9cyx6, T9cyx6;
wire Bacyx6, Jacyx6, Racyx6, Zacyx6, Hbcyx6, Pbcyx6, Xbcyx6, Fccyx6, Nccyx6, Vccyx6;
wire Ddcyx6, Ldcyx6, Tdcyx6, Becyx6, Jecyx6, Recyx6, Zecyx6, Hfcyx6, Pfcyx6, Xfcyx6;
wire Fgcyx6, Ngcyx6, Vgcyx6, Dhcyx6, Lhcyx6, Thcyx6, Bicyx6, Jicyx6, Ricyx6, Zicyx6;
wire Hjcyx6, Pjcyx6, Xjcyx6, Fkcyx6, Nkcyx6, Vkcyx6, Dlcyx6, Llcyx6, Tlcyx6, Bmcyx6;
wire Jmcyx6, Rmcyx6, Zmcyx6, Hncyx6, Pncyx6, Xncyx6, Focyx6, Nocyx6, Vocyx6, Dpcyx6;
wire Lpcyx6, Tpcyx6, Bqcyx6, Jqcyx6, Rqcyx6, Zqcyx6, Hrcyx6, Prcyx6, Xrcyx6, Fscyx6;
wire Nscyx6, Vscyx6, Dtcyx6, Ltcyx6, Ttcyx6, Bucyx6, Jucyx6, Rucyx6, Zucyx6, Hvcyx6;
wire Pvcyx6, Xvcyx6, Fwcyx6, Nwcyx6, Vwcyx6, Dxcyx6, Lxcyx6, Txcyx6, Bycyx6, Jycyx6;
wire Rycyx6, Zycyx6, Hzcyx6, Pzcyx6, Xzcyx6, F0dyx6, N0dyx6, V0dyx6, D1dyx6, L1dyx6;
wire T1dyx6, B2dyx6, J2dyx6, R2dyx6, Z2dyx6, H3dyx6, P3dyx6, X3dyx6, F4dyx6, N4dyx6;
wire V4dyx6, D5dyx6, L5dyx6, T5dyx6, B6dyx6, J6dyx6, R6dyx6, Z6dyx6, H7dyx6, P7dyx6;
wire X7dyx6, F8dyx6, N8dyx6, V8dyx6, D9dyx6, L9dyx6, T9dyx6, Badyx6, Jadyx6, Radyx6;
wire Zadyx6, Hbdyx6, Pbdyx6, Xbdyx6, Fcdyx6, Ncdyx6, Vcdyx6, Dddyx6, Lddyx6, Tddyx6;
wire Bedyx6, Jedyx6, Redyx6, Zedyx6, Hfdyx6, Pfdyx6, Xfdyx6, Fgdyx6, Ngdyx6, Vgdyx6;
wire Dhdyx6, Lhdyx6, Thdyx6, Bidyx6, Jidyx6, Ridyx6, Zidyx6, Hjdyx6, Pjdyx6, Xjdyx6;
wire Fkdyx6, Nkdyx6, Vkdyx6, Dldyx6, Lldyx6, Tldyx6, Bmdyx6, Jmdyx6, Rmdyx6, Zmdyx6;
wire Hndyx6, Pndyx6, Xndyx6, Fodyx6, Nodyx6, Vodyx6, Dpdyx6, Lpdyx6, Tpdyx6, Bqdyx6;
wire Jqdyx6, Rqdyx6, Zqdyx6, Hrdyx6, Prdyx6, Xrdyx6, Fsdyx6, Nsdyx6, Vsdyx6, Dtdyx6;
wire Ltdyx6, Ttdyx6, Budyx6, Judyx6, Rudyx6, Zudyx6, Hvdyx6, Pvdyx6, Xvdyx6, Fwdyx6;
wire Nwdyx6, Vwdyx6, Dxdyx6, Lxdyx6, Txdyx6, Bydyx6, Jydyx6, Rydyx6, Zydyx6, Hzdyx6;
wire Pzdyx6, Xzdyx6, F0eyx6, N0eyx6, V0eyx6, D1eyx6, L1eyx6, T1eyx6, B2eyx6, J2eyx6;
wire R2eyx6, Z2eyx6, H3eyx6, P3eyx6, X3eyx6, F4eyx6, N4eyx6, V4eyx6, D5eyx6, L5eyx6;
wire T5eyx6, B6eyx6, J6eyx6, R6eyx6, Z6eyx6, H7eyx6, P7eyx6, X7eyx6, F8eyx6, N8eyx6;
wire V8eyx6, D9eyx6, L9eyx6, T9eyx6, Baeyx6, Jaeyx6, Raeyx6, Zaeyx6, Hbeyx6, Pbeyx6;
wire Xbeyx6, Fceyx6, Nceyx6, Vceyx6, Ddeyx6, Ldeyx6, Tdeyx6, Beeyx6, Jeeyx6, Reeyx6;
wire Zeeyx6, Hfeyx6, Pfeyx6, Xfeyx6, Fgeyx6, Ngeyx6, Vgeyx6, Dheyx6, Lheyx6, Theyx6;
wire Bieyx6, Jieyx6, Rieyx6, Zieyx6, Hjeyx6, Pjeyx6, Xjeyx6, Fkeyx6, Nkeyx6, Vkeyx6;
wire Dleyx6, Lleyx6, Tleyx6, Bmeyx6, Jmeyx6, Rmeyx6, Zmeyx6, Hneyx6, Pneyx6, Xneyx6;
wire Foeyx6, Noeyx6, Voeyx6, Dpeyx6, Lpeyx6, Tpeyx6, Bqeyx6, Jqeyx6, Rqeyx6, Zqeyx6;
wire Hreyx6, Preyx6, Xreyx6, Fseyx6, Nseyx6, Vseyx6, Dteyx6, Lteyx6, Tteyx6, Bueyx6;
wire Jueyx6, Rueyx6, Zueyx6, Hveyx6, Pveyx6, Xveyx6, Fweyx6, Nweyx6, Vweyx6, Dxeyx6;
wire Lxeyx6, Txeyx6, Byeyx6, Jyeyx6, Ryeyx6, Zyeyx6, Hzeyx6, Pzeyx6, Xzeyx6, F0fyx6;
wire N0fyx6, V0fyx6, D1fyx6, L1fyx6, T1fyx6, B2fyx6, J2fyx6, R2fyx6, Z2fyx6, H3fyx6;
wire P3fyx6, X3fyx6, F4fyx6, N4fyx6, V4fyx6, D5fyx6, L5fyx6, T5fyx6, B6fyx6, J6fyx6;
wire R6fyx6, Z6fyx6, H7fyx6, P7fyx6, X7fyx6, F8fyx6, N8fyx6, V8fyx6, D9fyx6, L9fyx6;
wire T9fyx6, Bafyx6, Jafyx6, Rafyx6, Zafyx6, Hbfyx6, Pbfyx6, Xbfyx6, Fcfyx6, Ncfyx6;
wire Vcfyx6, Ddfyx6, Ldfyx6, Tdfyx6, Befyx6, Jefyx6, Refyx6, Zefyx6, Hffyx6, Pffyx6;
wire Xffyx6, Fgfyx6, Ngfyx6, Vgfyx6, Dhfyx6, Lhfyx6, Thfyx6, Bifyx6, Jifyx6, Rifyx6;
wire Zifyx6, Hjfyx6, Pjfyx6, Xjfyx6, Fkfyx6, Nkfyx6, Vkfyx6, Dlfyx6, Llfyx6, Tlfyx6;
wire Bmfyx6, Jmfyx6, Rmfyx6, Zmfyx6, Hnfyx6, Pnfyx6, Xnfyx6, Fofyx6, Nofyx6, Vofyx6;
wire Dpfyx6, Lpfyx6, Tpfyx6, Bqfyx6, Jqfyx6, Rqfyx6, Zqfyx6, Hrfyx6, Prfyx6, Xrfyx6;
wire Fsfyx6, Nsfyx6, Vsfyx6, Dtfyx6, Ltfyx6, Ttfyx6, Bufyx6, Jufyx6, Rufyx6, Zufyx6;
wire Hvfyx6, Pvfyx6, Xvfyx6, Fwfyx6, Nwfyx6, Vwfyx6, Dxfyx6, Lxfyx6, Txfyx6, Byfyx6;
wire Jyfyx6, Ryfyx6, Zyfyx6, Hzfyx6, Pzfyx6, Xzfyx6, F0gyx6, N0gyx6, V0gyx6, D1gyx6;
wire L1gyx6, T1gyx6, B2gyx6, J2gyx6, R2gyx6, Z2gyx6, H3gyx6, P3gyx6, X3gyx6, F4gyx6;
wire N4gyx6, V4gyx6, D5gyx6, L5gyx6, T5gyx6, B6gyx6, J6gyx6, R6gyx6, Z6gyx6, H7gyx6;
wire P7gyx6, X7gyx6, F8gyx6, N8gyx6, V8gyx6, D9gyx6, L9gyx6, T9gyx6, Bagyx6, Jagyx6;
wire Ragyx6, Zagyx6, Hbgyx6, Pbgyx6, Xbgyx6, Fcgyx6, Ncgyx6, Vcgyx6, Ddgyx6, Ldgyx6;
wire Tdgyx6, Begyx6, Jegyx6, Regyx6, Zegyx6, Hfgyx6, Pfgyx6, Xfgyx6, Fggyx6, Nggyx6;
wire Vggyx6, Dhgyx6, Lhgyx6, Thgyx6, Bigyx6, Jigyx6, Rigyx6, Zigyx6, Hjgyx6, Pjgyx6;
wire Xjgyx6, Fkgyx6, Nkgyx6, Vkgyx6, Dlgyx6, Llgyx6, Tlgyx6, Bmgyx6, Jmgyx6, Rmgyx6;
wire Zmgyx6, Hngyx6, Pngyx6, Xngyx6, Fogyx6, Nogyx6, Vogyx6, Dpgyx6, Lpgyx6, Tpgyx6;
wire Bqgyx6, Jqgyx6, Rqgyx6, Zqgyx6, Hrgyx6, Prgyx6, Xrgyx6, Fsgyx6, Nsgyx6, Vsgyx6;
wire Dtgyx6, Ltgyx6, Ttgyx6, Bugyx6, Jugyx6, Rugyx6, Zugyx6, Hvgyx6, Pvgyx6, Xvgyx6;
wire Fwgyx6, Nwgyx6, Vwgyx6, Dxgyx6, Lxgyx6, Txgyx6, Bygyx6, Jygyx6, Rygyx6, Zygyx6;
wire Hzgyx6, Pzgyx6, Xzgyx6, F0hyx6, N0hyx6, V0hyx6, D1hyx6, L1hyx6, T1hyx6, B2hyx6;
wire J2hyx6, R2hyx6, Z2hyx6, H3hyx6, P3hyx6, X3hyx6, F4hyx6, N4hyx6, V4hyx6, D5hyx6;
wire L5hyx6, T5hyx6, B6hyx6, J6hyx6, R6hyx6, Z6hyx6, H7hyx6, P7hyx6, X7hyx6, F8hyx6;
wire N8hyx6, V8hyx6, D9hyx6, L9hyx6, T9hyx6, Bahyx6, Jahyx6, Rahyx6, Zahyx6, Hbhyx6;
wire Pbhyx6, Xbhyx6, Fchyx6, Nchyx6, Vchyx6, Ddhyx6, Ldhyx6, Tdhyx6, Behyx6, Jehyx6;
wire Rehyx6, Zehyx6, Hfhyx6, Pfhyx6, Xfhyx6, Fghyx6, Nghyx6, Vghyx6, Dhhyx6, Lhhyx6;
wire Thhyx6, Bihyx6, Jihyx6, Rihyx6, Zihyx6, Hjhyx6, Pjhyx6, Xjhyx6, Fkhyx6, Nkhyx6;
wire Vkhyx6, Dlhyx6, Llhyx6, Tlhyx6, Bmhyx6, Jmhyx6, Rmhyx6, Zmhyx6, Hnhyx6, Pnhyx6;
wire Xnhyx6, Fohyx6, Nohyx6, Vohyx6, Dphyx6, Lphyx6, Tphyx6, Bqhyx6, Jqhyx6, Rqhyx6;
wire Zqhyx6, Hrhyx6, Prhyx6, Xrhyx6, Fshyx6, Nshyx6, Vshyx6, Dthyx6, Lthyx6, Tthyx6;
wire Buhyx6, Juhyx6, Ruhyx6, Zuhyx6, Hvhyx6, Pvhyx6, Xvhyx6, Fwhyx6, Nwhyx6, Vwhyx6;
wire Dxhyx6, Lxhyx6, Txhyx6, Byhyx6, Jyhyx6, Ryhyx6, Zyhyx6, Hzhyx6, Pzhyx6, Xzhyx6;
wire F0iyx6, N0iyx6, V0iyx6, D1iyx6, L1iyx6, T1iyx6, B2iyx6, J2iyx6, R2iyx6, Z2iyx6;
wire H3iyx6, P3iyx6, X3iyx6, F4iyx6, N4iyx6, V4iyx6, D5iyx6, L5iyx6, T5iyx6, B6iyx6;
wire J6iyx6, R6iyx6, Z6iyx6, H7iyx6, P7iyx6, X7iyx6, F8iyx6, N8iyx6, V8iyx6, D9iyx6;
wire L9iyx6, T9iyx6, Baiyx6, Jaiyx6, Raiyx6, Zaiyx6, Hbiyx6, Pbiyx6, Xbiyx6, Fciyx6;
wire Nciyx6, Vciyx6, Ddiyx6, Ldiyx6, Tdiyx6, Beiyx6, Jeiyx6, Reiyx6, Zeiyx6, Hfiyx6;
wire Pfiyx6, Xfiyx6, Fgiyx6, Ngiyx6, Vgiyx6, Dhiyx6, Lhiyx6, Thiyx6, Biiyx6, Jiiyx6;
wire Riiyx6, Ziiyx6, Hjiyx6, Pjiyx6, Xjiyx6, Fkiyx6, Nkiyx6, Vkiyx6, Dliyx6, Lliyx6;
wire Tliyx6, Bmiyx6, Jmiyx6, Rmiyx6, Zmiyx6, Hniyx6, Pniyx6, Xniyx6, Foiyx6, Noiyx6;
wire Voiyx6, Dpiyx6, Lpiyx6, Tpiyx6, Bqiyx6, Jqiyx6, Rqiyx6, Zqiyx6, Hriyx6, Priyx6;
wire Xriyx6, Fsiyx6, Nsiyx6, Vsiyx6, Dtiyx6, Ltiyx6, Ttiyx6, Buiyx6, Juiyx6, Ruiyx6;
wire Zuiyx6, Hviyx6, Pviyx6, Xviyx6, Fwiyx6, Nwiyx6, Vwiyx6, Dxiyx6, Lxiyx6, Txiyx6;
wire Byiyx6, Jyiyx6, Ryiyx6, Zyiyx6, Hziyx6, Pziyx6, Xziyx6, F0jyx6, N0jyx6, V0jyx6;
wire D1jyx6, L1jyx6, T1jyx6, B2jyx6, J2jyx6, R2jyx6, Z2jyx6, H3jyx6, P3jyx6, X3jyx6;
wire F4jyx6, N4jyx6, V4jyx6, D5jyx6, L5jyx6, T5jyx6, B6jyx6, J6jyx6, R6jyx6, Z6jyx6;
wire H7jyx6, P7jyx6, X7jyx6, F8jyx6, N8jyx6, V8jyx6, D9jyx6, L9jyx6, T9jyx6, Bajyx6;
wire Jajyx6, Rajyx6, Zajyx6, Hbjyx6, Pbjyx6, Xbjyx6, Fcjyx6, Ncjyx6, Vcjyx6, Ddjyx6;
wire Ldjyx6, Tdjyx6, Bejyx6, Jejyx6, Rejyx6, Zejyx6, Hfjyx6, Pfjyx6, Xfjyx6, Fgjyx6;
wire Ngjyx6, Vgjyx6, Dhjyx6, Lhjyx6, Thjyx6, Bijyx6, Jijyx6, Rijyx6, Zijyx6, Hjjyx6;
wire Pjjyx6, Xjjyx6, Fkjyx6, Nkjyx6, Vkjyx6, Dljyx6, Lljyx6, Tljyx6, Bmjyx6, Jmjyx6;
wire Rmjyx6, Zmjyx6, Hnjyx6, Pnjyx6, Xnjyx6, Fojyx6, Nojyx6, Vojyx6, Dpjyx6, Lpjyx6;
wire Tpjyx6, Bqjyx6, Jqjyx6, Rqjyx6, Zqjyx6, Hrjyx6, Prjyx6, Xrjyx6, Fsjyx6, Nsjyx6;
wire Vsjyx6, Dtjyx6, Ltjyx6, Ttjyx6, Bujyx6, Jujyx6, Rujyx6, Zujyx6, Hvjyx6, Pvjyx6;
wire Xvjyx6, Fwjyx6, Nwjyx6, Vwjyx6, Dxjyx6, Lxjyx6, Txjyx6, Byjyx6, Jyjyx6, Ryjyx6;
wire Zyjyx6, Hzjyx6, Pzjyx6, Xzjyx6, F0kyx6, N0kyx6, V0kyx6, D1kyx6, L1kyx6, T1kyx6;
wire B2kyx6, J2kyx6, R2kyx6, Z2kyx6, H3kyx6, P3kyx6, X3kyx6, F4kyx6, N4kyx6, V4kyx6;
wire D5kyx6, L5kyx6, T5kyx6, B6kyx6, J6kyx6, R6kyx6, Z6kyx6, H7kyx6, P7kyx6, X7kyx6;
wire F8kyx6, N8kyx6, V8kyx6, D9kyx6, L9kyx6, T9kyx6, Bakyx6, Jakyx6, Rakyx6, Zakyx6;
wire Hbkyx6, Pbkyx6, Xbkyx6, Fckyx6, Nckyx6, Vckyx6, Ddkyx6, Ldkyx6, Tdkyx6, Bekyx6;
wire Jekyx6, Rekyx6, Zekyx6, Hfkyx6, Pfkyx6, Xfkyx6, Fgkyx6, Ngkyx6, Vgkyx6, Dhkyx6;
wire Lhkyx6, Thkyx6, Bikyx6, Jikyx6, Rikyx6, Zikyx6, Hjkyx6, Pjkyx6, Xjkyx6, Fkkyx6;
wire Nkkyx6, Vkkyx6, Dlkyx6, Llkyx6, Tlkyx6, Bmkyx6, Jmkyx6, Rmkyx6, Zmkyx6, Hnkyx6;
wire Pnkyx6, Xnkyx6, Fokyx6, Nokyx6, Vokyx6, Dpkyx6, Lpkyx6, Tpkyx6, Bqkyx6, Jqkyx6;
wire Rqkyx6, Zqkyx6, Hrkyx6, Prkyx6, Xrkyx6, Fskyx6, Nskyx6, Vskyx6, Dtkyx6, Ltkyx6;
wire Ttkyx6, Bukyx6, Jukyx6, Rukyx6, Zukyx6, Hvkyx6, Pvkyx6, Xvkyx6, Fwkyx6, Nwkyx6;
wire Vwkyx6, Dxkyx6, Lxkyx6, Txkyx6, Bykyx6, Jykyx6, Rykyx6, Zykyx6, Hzkyx6, Pzkyx6;
wire Xzkyx6, F0lyx6, N0lyx6, V0lyx6, D1lyx6, L1lyx6, T1lyx6, B2lyx6, J2lyx6, R2lyx6;
wire Z2lyx6, H3lyx6, P3lyx6, X3lyx6, F4lyx6, N4lyx6, V4lyx6, D5lyx6, L5lyx6, T5lyx6;
wire B6lyx6, J6lyx6, R6lyx6, Z6lyx6, H7lyx6, P7lyx6, X7lyx6, F8lyx6, N8lyx6, V8lyx6;
wire D9lyx6, L9lyx6, T9lyx6, Balyx6, Jalyx6, Ralyx6, Zalyx6, Hblyx6, Pblyx6, Xblyx6;
wire Fclyx6, Nclyx6, Vclyx6, Ddlyx6, Ldlyx6, Tdlyx6, Belyx6, Jelyx6, Relyx6, Zelyx6;
wire Hflyx6, Pflyx6, Xflyx6, Fglyx6, Nglyx6, Vglyx6, Dhlyx6, Lhlyx6, Thlyx6, Bilyx6;
wire Jilyx6, Rilyx6, Zilyx6, Hjlyx6, Pjlyx6, Xjlyx6, Fklyx6, Nklyx6, Vklyx6, Dllyx6;
wire Lllyx6, Tllyx6, Bmlyx6, Jmlyx6, Rmlyx6, Zmlyx6, Hnlyx6, Pnlyx6, Xnlyx6, Folyx6;
wire Nolyx6, Volyx6, Dplyx6, Lplyx6, Tplyx6, Bqlyx6, Jqlyx6, Rqlyx6, Zqlyx6, Hrlyx6;
wire Prlyx6, Xrlyx6, Fslyx6, Nslyx6, Vslyx6, Dtlyx6, Ltlyx6, Ttlyx6, Bulyx6, Julyx6;
wire Rulyx6, Zulyx6, Hvlyx6, Pvlyx6, Xvlyx6, Fwlyx6, Nwlyx6, Vwlyx6, Dxlyx6, Lxlyx6;
wire Txlyx6, Bylyx6, Jylyx6, Rylyx6, Zylyx6, Hzlyx6, Pzlyx6, Xzlyx6, F0myx6, N0myx6;
wire V0myx6, D1myx6, L1myx6, T1myx6, B2myx6, J2myx6, R2myx6, Z2myx6, H3myx6, P3myx6;
wire X3myx6, F4myx6, N4myx6, V4myx6, D5myx6, L5myx6, T5myx6, B6myx6, J6myx6, R6myx6;
wire Z6myx6, H7myx6, P7myx6, X7myx6, F8myx6, N8myx6, V8myx6, D9myx6, L9myx6, T9myx6;
wire Bamyx6, Jamyx6, Ramyx6, Zamyx6, Hbmyx6, Pbmyx6, Xbmyx6, Fcmyx6, Ncmyx6, Vcmyx6;
wire Ddmyx6, Ldmyx6, Tdmyx6, Bemyx6, Jemyx6, Remyx6, Zemyx6, Hfmyx6, Pfmyx6, Xfmyx6;
wire Fgmyx6, Ngmyx6, Vgmyx6, Dhmyx6, Lhmyx6, Thmyx6, Bimyx6, Jimyx6, Rimyx6, Zimyx6;
wire Hjmyx6, Pjmyx6, Xjmyx6, Fkmyx6, Nkmyx6, Vkmyx6, Dlmyx6, Llmyx6, Tlmyx6, Bmmyx6;
wire Jmmyx6, Rmmyx6, Zmmyx6, Hnmyx6, Pnmyx6, Xnmyx6, Fomyx6, Nomyx6, Vomyx6, Dpmyx6;
wire Lpmyx6, Tpmyx6, Bqmyx6, Jqmyx6, Rqmyx6, Zqmyx6, Hrmyx6, Prmyx6, Xrmyx6, Fsmyx6;
wire Nsmyx6, Vsmyx6, Dtmyx6, Ltmyx6, Ttmyx6, Bumyx6, Jumyx6, Rumyx6, Zumyx6, Hvmyx6;
wire Pvmyx6, Xvmyx6, Fwmyx6, Nwmyx6, Vwmyx6, Dxmyx6, Lxmyx6, Txmyx6, Bymyx6, Jymyx6;
wire Rymyx6, Zymyx6, Hzmyx6, Pzmyx6, Xzmyx6, F0nyx6, N0nyx6, V0nyx6, D1nyx6, L1nyx6;
wire T1nyx6, B2nyx6, J2nyx6, R2nyx6, Z2nyx6, H3nyx6, P3nyx6, X3nyx6, F4nyx6, N4nyx6;
wire V4nyx6, D5nyx6, L5nyx6, T5nyx6, B6nyx6, J6nyx6, R6nyx6, Z6nyx6, H7nyx6, P7nyx6;
wire X7nyx6, F8nyx6, N8nyx6, V8nyx6, D9nyx6, L9nyx6, T9nyx6, Banyx6, Janyx6, Ranyx6;
wire Zanyx6, Hbnyx6, Pbnyx6, Xbnyx6, Fcnyx6, Ncnyx6, Vcnyx6, Ddnyx6, Ldnyx6, Tdnyx6;
wire Benyx6, Jenyx6, Renyx6, Zenyx6, Hfnyx6, Pfnyx6, Xfnyx6, Fgnyx6, Ngnyx6, Vgnyx6;
wire Dhnyx6, Lhnyx6, Thnyx6, Binyx6, Jinyx6, Rinyx6, Zinyx6, Hjnyx6, Pjnyx6, Xjnyx6;
wire Fknyx6, Nknyx6, Vknyx6, Dlnyx6, Llnyx6, Tlnyx6, Bmnyx6, Jmnyx6, Rmnyx6, Zmnyx6;
wire Hnnyx6, Pnnyx6, Xnnyx6, Fonyx6, Nonyx6, Vonyx6, Dpnyx6, Lpnyx6, Tpnyx6, Bqnyx6;
wire Jqnyx6, Rqnyx6, Zqnyx6, Hrnyx6, Prnyx6, Xrnyx6, Fsnyx6, Nsnyx6, Vsnyx6, Dtnyx6;
wire Ltnyx6, Ttnyx6, Bunyx6, Junyx6, Runyx6, Zunyx6, Hvnyx6, Pvnyx6, Xvnyx6, Fwnyx6;
wire Nwnyx6, Vwnyx6, Dxnyx6, Lxnyx6, Txnyx6, Bynyx6, Jynyx6, Rynyx6, Zynyx6, Hznyx6;
wire Pznyx6, Xznyx6, F0oyx6, N0oyx6, V0oyx6, D1oyx6, L1oyx6, T1oyx6, B2oyx6, J2oyx6;
wire R2oyx6, Z2oyx6, H3oyx6, P3oyx6, X3oyx6, F4oyx6, N4oyx6, V4oyx6, D5oyx6, L5oyx6;
wire T5oyx6, B6oyx6, J6oyx6, R6oyx6, Z6oyx6, H7oyx6, P7oyx6, X7oyx6, F8oyx6, N8oyx6;
wire V8oyx6, D9oyx6, L9oyx6, T9oyx6, Baoyx6, Jaoyx6, Raoyx6, Zaoyx6, Hboyx6, Pboyx6;
wire Xboyx6, Fcoyx6, Ncoyx6, Vcoyx6, Ddoyx6, Ldoyx6, Tdoyx6, Beoyx6, Jeoyx6, Reoyx6;
wire Zeoyx6, Hfoyx6, Pfoyx6, Xfoyx6, Fgoyx6, Ngoyx6, Vgoyx6, Dhoyx6, Lhoyx6, Thoyx6;
wire Bioyx6, Jioyx6, Rioyx6, Zioyx6, Hjoyx6, Pjoyx6, Xjoyx6, Fkoyx6, Nkoyx6, Vkoyx6;
wire Dloyx6, Lloyx6, Tloyx6, Bmoyx6, Jmoyx6, Rmoyx6, Zmoyx6, Hnoyx6, Pnoyx6, Xnoyx6;
wire Fooyx6, Nooyx6, Vooyx6, Dpoyx6, Lpoyx6, Tpoyx6, Bqoyx6, Jqoyx6, Rqoyx6, Zqoyx6;
wire Hroyx6, Proyx6, Xroyx6, Fsoyx6, Nsoyx6, Vsoyx6, Dtoyx6, Ltoyx6, Ttoyx6, Buoyx6;
wire Juoyx6, Ruoyx6, Zuoyx6, Hvoyx6, Pvoyx6, Xvoyx6, Fwoyx6, Nwoyx6, Vwoyx6, Dxoyx6;
wire Lxoyx6, Txoyx6, Byoyx6, Jyoyx6, Ryoyx6, Zyoyx6, Hzoyx6, Pzoyx6, Xzoyx6, F0pyx6;
wire N0pyx6, V0pyx6, D1pyx6, L1pyx6, T1pyx6, B2pyx6, J2pyx6, R2pyx6, Z2pyx6, H3pyx6;
wire P3pyx6, X3pyx6, F4pyx6, N4pyx6, V4pyx6, D5pyx6, L5pyx6, T5pyx6, B6pyx6, J6pyx6;
wire R6pyx6, Z6pyx6, H7pyx6, P7pyx6, X7pyx6, F8pyx6, N8pyx6, V8pyx6, D9pyx6, L9pyx6;
wire T9pyx6, Bapyx6, Japyx6, Rapyx6, Zapyx6, Hbpyx6, Pbpyx6, Xbpyx6, Fcpyx6, Ncpyx6;
wire Vcpyx6, Ddpyx6, Ldpyx6, Tdpyx6, Bepyx6, Jepyx6, Repyx6, Zepyx6, Hfpyx6, Pfpyx6;
wire Xfpyx6, Fgpyx6, Ngpyx6, Vgpyx6, Dhpyx6, Lhpyx6, Thpyx6, Bipyx6, Jipyx6, Ripyx6;
wire Zipyx6, Hjpyx6, Pjpyx6, Xjpyx6, Fkpyx6, Nkpyx6, Vkpyx6, Dlpyx6, Llpyx6, Tlpyx6;
wire Bmpyx6, Jmpyx6, Rmpyx6, Zmpyx6, Hnpyx6, Pnpyx6, Xnpyx6, Fopyx6, Nopyx6, Vopyx6;
wire Dppyx6, Lppyx6, Tppyx6, Bqpyx6, Jqpyx6, Rqpyx6, Zqpyx6, Hrpyx6, Prpyx6, Xrpyx6;
wire Fspyx6, Nspyx6, Vspyx6, Dtpyx6, Ltpyx6, Ttpyx6, Bupyx6, Jupyx6, Rupyx6, Zupyx6;
wire Hvpyx6, Pvpyx6, Xvpyx6, Fwpyx6, Nwpyx6, Vwpyx6, Dxpyx6, Lxpyx6, Txpyx6, Bypyx6;
wire Jypyx6, Rypyx6, Zypyx6, Hzpyx6, Pzpyx6, Xzpyx6, F0qyx6, N0qyx6, V0qyx6, D1qyx6;
wire L1qyx6, T1qyx6, B2qyx6, J2qyx6, R2qyx6, Z2qyx6, H3qyx6, P3qyx6, X3qyx6, F4qyx6;
wire N4qyx6, V4qyx6, D5qyx6, L5qyx6, T5qyx6, B6qyx6, J6qyx6, R6qyx6, Z6qyx6, H7qyx6;
wire P7qyx6, X7qyx6, F8qyx6, N8qyx6, V8qyx6, D9qyx6, L9qyx6, T9qyx6, Baqyx6, Jaqyx6;
wire Raqyx6, Zaqyx6, Hbqyx6, Pbqyx6, Xbqyx6, Fcqyx6, Ncqyx6, Vcqyx6, Ddqyx6, Ldqyx6;
wire Tdqyx6, Beqyx6, Jeqyx6, Reqyx6, Zeqyx6, Hfqyx6, Pfqyx6, Xfqyx6, Fgqyx6, Ngqyx6;
wire Vgqyx6, Dhqyx6, Lhqyx6, Thqyx6, Biqyx6, Jiqyx6, Riqyx6, Ziqyx6, Hjqyx6, Pjqyx6;
wire Xjqyx6, Fkqyx6, Nkqyx6, Vkqyx6, Dlqyx6, Llqyx6, Tlqyx6, Bmqyx6, Jmqyx6, Rmqyx6;
wire Zmqyx6, Hnqyx6, Pnqyx6, Xnqyx6, Foqyx6, Noqyx6, Voqyx6, Dpqyx6, Lpqyx6, Tpqyx6;
wire Bqqyx6, Jqqyx6, Rqqyx6, Zqqyx6, Hrqyx6, Prqyx6, Xrqyx6, Fsqyx6, Nsqyx6, Vsqyx6;
wire Dtqyx6, Ltqyx6, Ttqyx6, Buqyx6, Juqyx6, Ruqyx6, Zuqyx6, Hvqyx6, Pvqyx6, Xvqyx6;
wire Fwqyx6, Nwqyx6, Vwqyx6, Dxqyx6, Lxqyx6, Txqyx6, Byqyx6, Jyqyx6, Ryqyx6, Zyqyx6;
wire Hzqyx6, Pzqyx6, Xzqyx6, F0ryx6, N0ryx6, V0ryx6, D1ryx6, L1ryx6, T1ryx6, B2ryx6;
wire J2ryx6, R2ryx6, Z2ryx6, H3ryx6, P3ryx6, X3ryx6, F4ryx6, N4ryx6, V4ryx6, D5ryx6;
wire L5ryx6, T5ryx6, B6ryx6, J6ryx6, R6ryx6, Z6ryx6, H7ryx6, P7ryx6, X7ryx6, F8ryx6;
wire N8ryx6, V8ryx6, D9ryx6, L9ryx6, T9ryx6, Baryx6, Jaryx6, Raryx6, Zaryx6, Hbryx6;
wire Pbryx6, Xbryx6, Fcryx6, Ncryx6, Vcryx6, Ddryx6, Ldryx6, Tdryx6, Beryx6, Jeryx6;
wire Reryx6, Zeryx6, Hfryx6, Pfryx6, Xfryx6, Fgryx6, Ngryx6, Vgryx6, Dhryx6, Lhryx6;
wire Thryx6, Biryx6, Jiryx6, Riryx6, Ziryx6, Hjryx6, Pjryx6, Xjryx6, Fkryx6, Nkryx6;
wire Vkryx6, Dlryx6, Llryx6, Tlryx6, Bmryx6, Jmryx6, Rmryx6, Zmryx6, Hnryx6, Pnryx6;
wire Xnryx6, Foryx6, Noryx6, Voryx6, Dpryx6, Lpryx6, Tpryx6, Bqryx6, Jqryx6, Rqryx6;
wire Zqryx6, Hrryx6, Prryx6, Xrryx6, Fsryx6, Nsryx6, Vsryx6, Dtryx6, Ltryx6, Ttryx6;
wire Buryx6, Juryx6, Ruryx6, Zuryx6, Hvryx6, Pvryx6, Xvryx6, Fwryx6, Nwryx6, Vwryx6;
wire Dxryx6, Lxryx6, Txryx6, Byryx6, Jyryx6, Ryryx6, Zyryx6, Hzryx6, Pzryx6, Xzryx6;
wire F0syx6, N0syx6, V0syx6, D1syx6, L1syx6, T1syx6, B2syx6, J2syx6, R2syx6, Z2syx6;
wire H3syx6, P3syx6, X3syx6, F4syx6, N4syx6, V4syx6, D5syx6, L5syx6, T5syx6, B6syx6;
wire J6syx6, R6syx6, Z6syx6, H7syx6, P7syx6, X7syx6, F8syx6, N8syx6, V8syx6, D9syx6;
wire L9syx6, T9syx6, Basyx6, Jasyx6, Rasyx6, Zasyx6, Hbsyx6, Pbsyx6, Xbsyx6, Fcsyx6;
wire Ncsyx6, Vcsyx6, Ddsyx6, Ldsyx6, Tdsyx6, Besyx6, Jesyx6, Resyx6, Zesyx6, Hfsyx6;
wire Pfsyx6, Xfsyx6, Fgsyx6, Ngsyx6, Vgsyx6, Dhsyx6, Lhsyx6, Thsyx6, Bisyx6, Jisyx6;
wire Risyx6, Zisyx6, Hjsyx6, Pjsyx6, Xjsyx6, Fksyx6, Nksyx6, Vksyx6, Dlsyx6, Llsyx6;
wire Tlsyx6, Bmsyx6, Jmsyx6, Rmsyx6, Zmsyx6, Hnsyx6, Pnsyx6, Xnsyx6, Fosyx6, Nosyx6;
wire Vosyx6, Dpsyx6, Lpsyx6, Tpsyx6, Bqsyx6, Jqsyx6, Rqsyx6, Zqsyx6, Hrsyx6, Prsyx6;
wire Xrsyx6, Fssyx6, Nssyx6, Vssyx6, Dtsyx6, Ltsyx6, Ttsyx6, Busyx6, Jusyx6, Rusyx6;
wire Zusyx6, Hvsyx6, Pvsyx6, Xvsyx6, Fwsyx6, Nwsyx6, Vwsyx6, Dxsyx6, Lxsyx6, Txsyx6;
wire Bysyx6, Jysyx6, Rysyx6, Zysyx6, Hzsyx6, Pzsyx6, Xzsyx6, F0tyx6, N0tyx6, V0tyx6;
wire D1tyx6, L1tyx6, T1tyx6, B2tyx6, J2tyx6, R2tyx6, Z2tyx6, H3tyx6, P3tyx6, X3tyx6;
wire F4tyx6, N4tyx6, V4tyx6, D5tyx6, L5tyx6, T5tyx6, B6tyx6, J6tyx6, R6tyx6, Z6tyx6;
wire H7tyx6, P7tyx6, X7tyx6, F8tyx6, N8tyx6, V8tyx6, D9tyx6, L9tyx6, T9tyx6, Batyx6;
wire Jatyx6, Ratyx6, Zatyx6, Hbtyx6, Pbtyx6, Xbtyx6, Fctyx6, Nctyx6, Vctyx6, Ddtyx6;
wire Ldtyx6, Tdtyx6, Betyx6, Jetyx6, Retyx6, Zetyx6, Hftyx6, Pftyx6, Xftyx6, Fgtyx6;
wire Ngtyx6, Vgtyx6, Dhtyx6, Lhtyx6, Thtyx6, Bityx6, Jityx6, Rityx6, Zityx6, Hjtyx6;
wire Pjtyx6, Xjtyx6, Fktyx6, Nktyx6, Vktyx6, Dltyx6, Lltyx6, Tltyx6, Bmtyx6, Jmtyx6;
wire Rmtyx6, Zmtyx6, Hntyx6, Pntyx6, Xntyx6, Fotyx6, Notyx6, Votyx6, Dptyx6, Lptyx6;
wire Tptyx6, Bqtyx6, Jqtyx6, Rqtyx6, Zqtyx6, Hrtyx6, Prtyx6, Xrtyx6, Fstyx6, Nstyx6;
wire Vstyx6, Dttyx6, Lttyx6, Tttyx6, Butyx6, Jutyx6, Rutyx6, Zutyx6, Hvtyx6, Pvtyx6;
wire Xvtyx6, Fwtyx6, Nwtyx6, Vwtyx6, Dxtyx6, Lxtyx6, Txtyx6, Bytyx6, Jytyx6, Rytyx6;
wire Zytyx6, Hztyx6, Pztyx6, Xztyx6, F0uyx6, N0uyx6, V0uyx6, D1uyx6, L1uyx6, T1uyx6;
wire B2uyx6, J2uyx6, R2uyx6, Z2uyx6, H3uyx6, P3uyx6, X3uyx6, F4uyx6, N4uyx6, V4uyx6;
wire D5uyx6, L5uyx6, T5uyx6, B6uyx6, J6uyx6, R6uyx6, Z6uyx6, H7uyx6, P7uyx6, X7uyx6;
wire F8uyx6, N8uyx6, V8uyx6, D9uyx6, L9uyx6, T9uyx6, Bauyx6, Jauyx6, Rauyx6, Zauyx6;
wire Hbuyx6, Pbuyx6, Xbuyx6, Fcuyx6, Ncuyx6, Vcuyx6, Dduyx6, Lduyx6, Tduyx6, Beuyx6;
wire Jeuyx6, Reuyx6, Zeuyx6, Hfuyx6, Pfuyx6, Xfuyx6, Fguyx6, Nguyx6, Vguyx6, Dhuyx6;
wire Lhuyx6, Thuyx6, Biuyx6, Jiuyx6, Riuyx6, Ziuyx6, Hjuyx6, Pjuyx6, Xjuyx6, Fkuyx6;
wire Nkuyx6, Vkuyx6, Dluyx6, Lluyx6, Tluyx6, Bmuyx6, Jmuyx6, Rmuyx6, Zmuyx6, Hnuyx6;
wire Pnuyx6, Xnuyx6, Fouyx6, Nouyx6, Vouyx6, Dpuyx6, Lpuyx6, Tpuyx6, Bquyx6, Jquyx6;
wire Rquyx6, Zquyx6, Hruyx6, Pruyx6, Xruyx6, Fsuyx6, Nsuyx6, Vsuyx6, Dtuyx6, Ltuyx6;
wire Ttuyx6, Buuyx6, Juuyx6, Ruuyx6, Zuuyx6, Hvuyx6, Pvuyx6, Xvuyx6, Fwuyx6, Nwuyx6;
wire Vwuyx6, Dxuyx6, Lxuyx6, Txuyx6, Byuyx6, Jyuyx6, Ryuyx6, Zyuyx6, Hzuyx6, Pzuyx6;
wire Xzuyx6, F0vyx6, N0vyx6, V0vyx6, D1vyx6, L1vyx6, T1vyx6, B2vyx6, J2vyx6, R2vyx6;
wire Z2vyx6, H3vyx6, P3vyx6, X3vyx6, F4vyx6, N4vyx6, V4vyx6, D5vyx6, L5vyx6, T5vyx6;
wire B6vyx6, J6vyx6, R6vyx6, Z6vyx6, H7vyx6, P7vyx6, X7vyx6, F8vyx6, N8vyx6, V8vyx6;
wire D9vyx6, L9vyx6, T9vyx6, Bavyx6, Javyx6, Ravyx6, Zavyx6, Hbvyx6, Pbvyx6, Xbvyx6;
wire Fcvyx6, Ncvyx6, Vcvyx6, Ddvyx6, Ldvyx6, Tdvyx6, Bevyx6, Jevyx6, Revyx6, Zevyx6;
wire Hfvyx6, Pfvyx6, Xfvyx6, Fgvyx6, Ngvyx6, Vgvyx6, Dhvyx6, Lhvyx6, Thvyx6, Bivyx6;
wire Jivyx6, Rivyx6, Zivyx6, Hjvyx6, Pjvyx6, Xjvyx6, Fkvyx6, Nkvyx6, Vkvyx6, Dlvyx6;
wire Llvyx6, Tlvyx6, Bmvyx6, Jmvyx6, Rmvyx6, Zmvyx6, Hnvyx6, Pnvyx6, Xnvyx6, Fovyx6;
wire Novyx6, Vovyx6, Dpvyx6, Lpvyx6, Tpvyx6, Bqvyx6, Jqvyx6, Rqvyx6, Zqvyx6, Hrvyx6;
wire Prvyx6, Xrvyx6, Fsvyx6, Nsvyx6, Vsvyx6, Dtvyx6, Ltvyx6, Ttvyx6, Buvyx6, Juvyx6;
wire Ruvyx6, Zuvyx6, Hvvyx6, Pvvyx6, Xvvyx6, Fwvyx6, Nwvyx6, Vwvyx6, Dxvyx6, Lxvyx6;
wire Txvyx6, Byvyx6, Jyvyx6, Ryvyx6, Zyvyx6, Hzvyx6, Pzvyx6, Xzvyx6, F0wyx6, N0wyx6;
wire V0wyx6, D1wyx6, L1wyx6, T1wyx6, B2wyx6, J2wyx6, R2wyx6, Z2wyx6, H3wyx6, P3wyx6;
wire X3wyx6, F4wyx6, N4wyx6, V4wyx6, D5wyx6, L5wyx6, T5wyx6, B6wyx6, J6wyx6, R6wyx6;
wire Z6wyx6, H7wyx6, P7wyx6, X7wyx6, F8wyx6, N8wyx6, V8wyx6, D9wyx6, L9wyx6, T9wyx6;
wire Bawyx6, Jawyx6, Rawyx6, Zawyx6, Hbwyx6, Pbwyx6, Xbwyx6, Fcwyx6, Ncwyx6, Vcwyx6;
wire Ddwyx6, Ldwyx6, Tdwyx6, Bewyx6, Jewyx6, Rewyx6, Zewyx6, Hfwyx6, Pfwyx6, Xfwyx6;
wire Fgwyx6, Ngwyx6, Vgwyx6, Dhwyx6, Lhwyx6, Thwyx6, Biwyx6, Jiwyx6, Riwyx6, Ziwyx6;
wire Hjwyx6, Pjwyx6, Xjwyx6, Fkwyx6, Nkwyx6, Vkwyx6, Dlwyx6, Llwyx6, Tlwyx6, Bmwyx6;
wire Jmwyx6, Rmwyx6, Zmwyx6, Hnwyx6, Pnwyx6, Xnwyx6, Fowyx6, Nowyx6, Vowyx6, Dpwyx6;
wire Lpwyx6, Tpwyx6, Bqwyx6, Jqwyx6, Rqwyx6, Zqwyx6, Hrwyx6, Prwyx6, Xrwyx6, Fswyx6;
wire Nswyx6, Vswyx6, Dtwyx6, Ltwyx6, Ttwyx6, Buwyx6, Juwyx6, Ruwyx6, Zuwyx6, Hvwyx6;
wire Pvwyx6, Xvwyx6, Fwwyx6, Nwwyx6, Vwwyx6, Dxwyx6, Lxwyx6, Txwyx6, Bywyx6, Jywyx6;
wire Rywyx6, Zywyx6, Hzwyx6, Pzwyx6, Xzwyx6, F0xyx6, N0xyx6, V0xyx6, D1xyx6, L1xyx6;
wire T1xyx6, B2xyx6, J2xyx6, R2xyx6, Z2xyx6, H3xyx6, P3xyx6, X3xyx6, F4xyx6, N4xyx6;
wire V4xyx6, D5xyx6, L5xyx6, T5xyx6, B6xyx6, J6xyx6, R6xyx6, Z6xyx6, H7xyx6, P7xyx6;
wire X7xyx6, F8xyx6, N8xyx6, V8xyx6, D9xyx6, L9xyx6, T9xyx6, Baxyx6, Jaxyx6, Raxyx6;
wire Zaxyx6, Hbxyx6, Pbxyx6, Xbxyx6, Fcxyx6, Ncxyx6, Vcxyx6, Ddxyx6, Ldxyx6, Tdxyx6;
wire Bexyx6, Jexyx6, Rexyx6, Zexyx6, Hfxyx6, Pfxyx6, Xfxyx6, Fgxyx6, Ngxyx6, Vgxyx6;
wire Dhxyx6, Lhxyx6, Thxyx6, Bixyx6, Jixyx6, Rixyx6, Zixyx6, Hjxyx6, Pjxyx6, Xjxyx6;
wire Fkxyx6, Nkxyx6, Vkxyx6, Dlxyx6, Llxyx6, Tlxyx6, Bmxyx6, Jmxyx6, Rmxyx6, Zmxyx6;
wire Hnxyx6, Pnxyx6, Xnxyx6, Foxyx6, Noxyx6, Voxyx6, Dpxyx6, Lpxyx6, Tpxyx6, Bqxyx6;
wire Jqxyx6, Rqxyx6, Zqxyx6, Hrxyx6, Prxyx6, Xrxyx6, Fsxyx6, Nsxyx6, Vsxyx6, Dtxyx6;
wire Ltxyx6, Ttxyx6, Buxyx6, Juxyx6, Ruxyx6, Zuxyx6, Hvxyx6, Pvxyx6, Xvxyx6, Fwxyx6;
wire Nwxyx6, Vwxyx6, Dxxyx6, Lxxyx6, Txxyx6, Byxyx6, Jyxyx6, Ryxyx6, Zyxyx6, Hzxyx6;
wire Pzxyx6, Xzxyx6, F0yyx6, N0yyx6, V0yyx6, D1yyx6, L1yyx6, T1yyx6, B2yyx6, J2yyx6;
wire R2yyx6, Z2yyx6, H3yyx6, P3yyx6, X3yyx6, F4yyx6, N4yyx6, V4yyx6, D5yyx6, L5yyx6;
wire T5yyx6, B6yyx6, J6yyx6, R6yyx6, Z6yyx6, H7yyx6, P7yyx6, X7yyx6, F8yyx6, N8yyx6;
wire V8yyx6, D9yyx6, L9yyx6, T9yyx6, Bayyx6, Jayyx6, Rayyx6, Zayyx6, Hbyyx6, Pbyyx6;
wire Xbyyx6, Fcyyx6, Ncyyx6, Vcyyx6, Ddyyx6, Ldyyx6, Tdyyx6, Beyyx6, Jeyyx6, Reyyx6;
wire Zeyyx6, Hfyyx6, Pfyyx6, Xfyyx6, Fgyyx6, Ngyyx6, Vgyyx6, Dhyyx6, Lhyyx6, Thyyx6;
wire Biyyx6, Jiyyx6, Riyyx6, Ziyyx6, Hjyyx6, Pjyyx6, Xjyyx6, Fkyyx6, Nkyyx6, Vkyyx6;
wire Dlyyx6, Llyyx6, Tlyyx6, Bmyyx6, Jmyyx6, Rmyyx6, Zmyyx6, Hnyyx6, Pnyyx6, Xnyyx6;
wire Foyyx6, Noyyx6, Voyyx6, Dpyyx6, Lpyyx6, Tpyyx6, Bqyyx6, Jqyyx6, Rqyyx6, Zqyyx6;
wire Hryyx6, Pryyx6, Xryyx6, Fsyyx6, Nsyyx6, Vsyyx6, Dtyyx6, Ltyyx6, Ttyyx6, Buyyx6;
wire Juyyx6, Ruyyx6, Zuyyx6, Hvyyx6, Pvyyx6, Xvyyx6, Fwyyx6, Nwyyx6, Vwyyx6, Dxyyx6;
wire Lxyyx6, Txyyx6, Byyyx6, Jyyyx6, Ryyyx6, Zyyyx6, Hzyyx6, Pzyyx6, Xzyyx6, F0zyx6;
wire N0zyx6, V0zyx6, D1zyx6, L1zyx6, T1zyx6, B2zyx6, J2zyx6, R2zyx6, Z2zyx6, H3zyx6;
wire P3zyx6, X3zyx6, F4zyx6, N4zyx6, V4zyx6, D5zyx6, L5zyx6, T5zyx6, B6zyx6, J6zyx6;
wire R6zyx6, Z6zyx6, H7zyx6, P7zyx6, X7zyx6, F8zyx6, N8zyx6, V8zyx6, D9zyx6, L9zyx6;
wire T9zyx6, Bazyx6, Jazyx6, Razyx6, Zazyx6, Hbzyx6, Pbzyx6, Xbzyx6, Fczyx6, Nczyx6;
wire Vczyx6, Ddzyx6, Ldzyx6, Tdzyx6, Bezyx6, Jezyx6, Rezyx6, Zezyx6, Hfzyx6, Pfzyx6;
wire Xfzyx6, Fgzyx6, Ngzyx6, Vgzyx6, Dhzyx6, Lhzyx6, Thzyx6, Bizyx6, Jizyx6, Rizyx6;
wire Zizyx6, Hjzyx6, Pjzyx6, Xjzyx6, Fkzyx6, Nkzyx6, Vkzyx6, Dlzyx6, Llzyx6, Tlzyx6;
wire Bmzyx6, Jmzyx6, Rmzyx6, Zmzyx6, Hnzyx6, Pnzyx6, Xnzyx6, Fozyx6, Nozyx6, Vozyx6;
wire Dpzyx6, Lpzyx6, Tpzyx6, Bqzyx6, Jqzyx6, Rqzyx6, Zqzyx6, Hrzyx6, Przyx6, Xrzyx6;
wire Fszyx6, Nszyx6, Vszyx6, Dtzyx6, Ltzyx6, Ttzyx6, Buzyx6, Juzyx6, Ruzyx6, Zuzyx6;
wire Hvzyx6, Pvzyx6, Xvzyx6, Fwzyx6, Nwzyx6, Vwzyx6, Dxzyx6, Lxzyx6, Txzyx6, Byzyx6;
wire Jyzyx6, Ryzyx6, Zyzyx6, Hzzyx6, Pzzyx6, Xzzyx6, F00zx6, N00zx6, V00zx6, D10zx6;
wire L10zx6, T10zx6, B20zx6, J20zx6, R20zx6, Z20zx6, H30zx6, P30zx6, X30zx6, F40zx6;
wire N40zx6, V40zx6, D50zx6, L50zx6, T50zx6, B60zx6, J60zx6, R60zx6, Z60zx6, H70zx6;
wire P70zx6, X70zx6, F80zx6, N80zx6, V80zx6, D90zx6, L90zx6, T90zx6, Ba0zx6, Ja0zx6;
wire Ra0zx6, Za0zx6, Hb0zx6, Pb0zx6, Xb0zx6, Fc0zx6, Nc0zx6, Vc0zx6, Dd0zx6, Ld0zx6;
wire Td0zx6, Be0zx6, Je0zx6, Re0zx6, Ze0zx6, Hf0zx6, Pf0zx6, Xf0zx6, Fg0zx6, Ng0zx6;
wire Vg0zx6, Dh0zx6, Lh0zx6, Th0zx6, Bi0zx6, Ji0zx6, Ri0zx6, Zi0zx6, Hj0zx6, Pj0zx6;
wire Xj0zx6, Fk0zx6, Nk0zx6, Vk0zx6, Dl0zx6, Ll0zx6, Tl0zx6, Bm0zx6, Jm0zx6, Rm0zx6;
wire Zm0zx6, Hn0zx6, Pn0zx6, Xn0zx6, Fo0zx6, No0zx6, Vo0zx6, Dp0zx6, Lp0zx6, Tp0zx6;
wire Bq0zx6, Jq0zx6, Rq0zx6, Zq0zx6, Hr0zx6, Pr0zx6, Xr0zx6, Fs0zx6, Ns0zx6, Vs0zx6;
wire Dt0zx6, Lt0zx6, Tt0zx6, Bu0zx6, Ju0zx6, Ru0zx6, Zu0zx6, Hv0zx6, Pv0zx6, Xv0zx6;
wire Fw0zx6, Nw0zx6, Vw0zx6, Dx0zx6, Lx0zx6, Tx0zx6, By0zx6, Jy0zx6, Ry0zx6, Zy0zx6;
wire Hz0zx6, Pz0zx6, Xz0zx6, F01zx6, N01zx6, V01zx6, D11zx6, L11zx6, T11zx6, B21zx6;
wire J21zx6, R21zx6, Z21zx6, H31zx6, P31zx6, X31zx6, F41zx6, N41zx6, V41zx6, D51zx6;
wire L51zx6, T51zx6, B61zx6, J61zx6, R61zx6, Z61zx6, H71zx6, P71zx6, X71zx6, F81zx6;
wire N81zx6, V81zx6, D91zx6, L91zx6, T91zx6, Ba1zx6, Ja1zx6, Ra1zx6, Za1zx6, Hb1zx6;
wire Pb1zx6, Xb1zx6, Fc1zx6, Nc1zx6, Vc1zx6, Dd1zx6, Ld1zx6, Td1zx6, Be1zx6, Je1zx6;
wire Re1zx6, Ze1zx6, Hf1zx6, Pf1zx6, Xf1zx6, Fg1zx6, Ng1zx6, Vg1zx6, Y0jhy6, G1jhy6;
wire O1jhy6, W1jhy6, E2jhy6, M2jhy6, U2jhy6, C3jhy6, K3jhy6, S3jhy6, A4jhy6, I4jhy6;
wire Q4jhy6, Y4jhy6, G5jhy6, O5jhy6, W5jhy6, E6jhy6, M6jhy6, U6jhy6, C7jhy6, K7jhy6;
wire S7jhy6, A8jhy6, I8jhy6, Q8jhy6, Y8jhy6, G9jhy6, O9jhy6, W9jhy6, Eajhy6, Majhy6;
wire Uajhy6, Cbjhy6, Kbjhy6, Sbjhy6, Acjhy6, Icjhy6, Qcjhy6, Ycjhy6, Gdjhy6, Odjhy6;
wire Wdjhy6, Eejhy6, Mejhy6, Uejhy6, Cfjhy6, Kfjhy6, Sfjhy6, Agjhy6, Igjhy6, Qgjhy6;
wire Ygjhy6, Ghjhy6, Ohjhy6, Whjhy6, Eijhy6, Mijhy6, Uijhy6, Cjjhy6, Kjjhy6, Sjjhy6;
wire Akjhy6, Ikjhy6, Qkjhy6, Ykjhy6, Gljhy6, Oljhy6, Wljhy6, Emjhy6, Mmjhy6, Umjhy6;
wire Cnjhy6, Knjhy6, Snjhy6, Aojhy6, Iojhy6, Qojhy6, Yojhy6, Gpjhy6, Opjhy6, Wpjhy6;
wire Eqjhy6, Mqjhy6, Uqjhy6, Crjhy6, Krjhy6, Srjhy6, Asjhy6, Isjhy6, Qsjhy6, Ysjhy6;
wire Gtjhy6, Otjhy6, Wtjhy6, Eujhy6, Mujhy6, Uujhy6, Cvjhy6, Kvjhy6, Svjhy6, Awjhy6;
wire Iwjhy6, Qwjhy6, Ywjhy6, Gxjhy6, Oxjhy6, Wxjhy6, Eyjhy6, Myjhy6, Uyjhy6, Czjhy6;
wire Kzjhy6, Szjhy6, A0khy6, I0khy6, Q0khy6, Y0khy6, G1khy6, O1khy6, W1khy6, E2khy6;
wire M2khy6, U2khy6, C3khy6, K3khy6, S3khy6, A4khy6, I4khy6, Q4khy6, Y4khy6, G5khy6;
wire O5khy6, W5khy6, E6khy6, M6khy6, U6khy6, C7khy6, K7khy6, S7khy6, A8khy6, I8khy6;
wire Q8khy6, Y8khy6, G9khy6, O9khy6, W9khy6, Eakhy6, Makhy6, Uakhy6, Cbkhy6, Kbkhy6;
wire Sbkhy6, Ackhy6, Ickhy6, Qckhy6, Yckhy6, Gdkhy6, Odkhy6, Wdkhy6, Eekhy6, Mekhy6;
wire Uekhy6, Cfkhy6, Kfkhy6, Sfkhy6, Agkhy6, Igkhy6, Qgkhy6, Ygkhy6, Ghkhy6, Ohkhy6;
wire Whkhy6, Eikhy6, Mikhy6, Uikhy6, Cjkhy6, Kjkhy6, Sjkhy6, Akkhy6, Ikkhy6, Qkkhy6;
wire Ykkhy6, Glkhy6, Olkhy6, Wlkhy6, Emkhy6, Mmkhy6, Umkhy6, Cnkhy6, Knkhy6, Snkhy6;
wire Aokhy6, Iokhy6, Qokhy6, Yokhy6, Gpkhy6, Opkhy6, Wpkhy6, Eqkhy6, Mqkhy6, Uqkhy6;
wire Crkhy6, Krkhy6, Srkhy6, Askhy6, Iskhy6, Qskhy6, Yskhy6, Gtkhy6, Otkhy6, Wtkhy6;
wire Eukhy6, Mukhy6, Uukhy6, Cvkhy6, Kvkhy6, Svkhy6, Awkhy6, Iwkhy6, Qwkhy6, Ywkhy6;
wire Gxkhy6, Oxkhy6, Wxkhy6, Eykhy6, Mykhy6, Uykhy6, Czkhy6, Kzkhy6, Szkhy6, A0lhy6;
wire I0lhy6, Q0lhy6, Y0lhy6, G1lhy6, O1lhy6, W1lhy6, E2lhy6, M2lhy6, U2lhy6, C3lhy6;
wire K3lhy6, S3lhy6, A4lhy6, I4lhy6, Q4lhy6, Y4lhy6, G5lhy6, O5lhy6, W5lhy6, E6lhy6;
wire M6lhy6, U6lhy6, C7lhy6, K7lhy6, S7lhy6, A8lhy6, I8lhy6, Q8lhy6, Y8lhy6, G9lhy6;
wire O9lhy6, W9lhy6, Ealhy6, Malhy6, Ualhy6, Cblhy6, Kblhy6, Sblhy6, Aclhy6, Iclhy6;
wire Qclhy6, Yclhy6, Gdlhy6, Odlhy6, Wdlhy6, Eelhy6, Melhy6, Uelhy6, Cflhy6, Kflhy6;
wire Sflhy6, Aglhy6, Iglhy6, Qglhy6, Yglhy6, Ghlhy6, Ohlhy6, Whlhy6, Eilhy6, Milhy6;
wire Uilhy6, Cjlhy6, Kjlhy6, Sjlhy6, Aklhy6, Iklhy6, Qklhy6, Yklhy6, Gllhy6, Ollhy6;
wire Wllhy6, Emlhy6, Mmlhy6, Umlhy6, Cnlhy6, Knlhy6, Snlhy6, Aolhy6, Iolhy6, Qolhy6;
wire Yolhy6, Gplhy6, Oplhy6, Wplhy6, Eqlhy6, Mqlhy6, Uqlhy6, Crlhy6, Krlhy6, Srlhy6;
wire Aslhy6, Islhy6, Qslhy6, Yslhy6, Gtlhy6, Otlhy6, Wtlhy6, Eulhy6, Mulhy6, Uulhy6;
wire Cvlhy6, Kvlhy6, Svlhy6, Awlhy6, Iwlhy6, Qwlhy6, Ywlhy6, Gxlhy6, Oxlhy6, Wxlhy6;
wire Eylhy6, Mylhy6, Uylhy6, Czlhy6, Kzlhy6, Szlhy6, A0mhy6, I0mhy6, Q0mhy6, Y0mhy6;
wire G1mhy6, O1mhy6, W1mhy6, E2mhy6, M2mhy6, U2mhy6, C3mhy6, K3mhy6, S3mhy6, A4mhy6;
wire I4mhy6, Q4mhy6, Y4mhy6, G5mhy6, O5mhy6, W5mhy6, E6mhy6, M6mhy6, U6mhy6, C7mhy6;
wire K7mhy6, S7mhy6, A8mhy6, I8mhy6, Q8mhy6, Y8mhy6, G9mhy6, O9mhy6, W9mhy6, Eamhy6;
wire Mamhy6, Uamhy6, Cbmhy6, Kbmhy6, Sbmhy6, Acmhy6, Icmhy6, Qcmhy6, Ycmhy6, Gdmhy6;
wire Odmhy6, Wdmhy6, Eemhy6, Memhy6, Uemhy6, Cfmhy6, Kfmhy6, Sfmhy6, Agmhy6, Igmhy6;
wire Qgmhy6, Ygmhy6, Ghmhy6, Ohmhy6, Whmhy6, Eimhy6, Mimhy6, Uimhy6, Cjmhy6, Kjmhy6;
wire Sjmhy6, Akmhy6, Ikmhy6, Qkmhy6, Ykmhy6, Glmhy6, Olmhy6, Wlmhy6, Emmhy6, Mmmhy6;
wire Ummhy6, Cnmhy6, Knmhy6, Snmhy6, Aomhy6, Iomhy6, Qomhy6, Yomhy6, Gpmhy6, Opmhy6;
wire Wpmhy6, Eqmhy6, Mqmhy6, Uqmhy6, Crmhy6, Krmhy6, Srmhy6, Asmhy6, Ismhy6, Qsmhy6;
wire Ysmhy6, Gtmhy6, Otmhy6, Wtmhy6, Eumhy6, Mumhy6, Uumhy6, Cvmhy6, Kvmhy6, Svmhy6;
wire Awmhy6, Iwmhy6, Qwmhy6, Ywmhy6, Gxmhy6, Oxmhy6, Wxmhy6, Eymhy6, Mymhy6, Uymhy6;
wire Czmhy6, Kzmhy6, Szmhy6, A0nhy6, I0nhy6, Q0nhy6, Y0nhy6, G1nhy6, O1nhy6, W1nhy6;
wire E2nhy6, M2nhy6, U2nhy6, C3nhy6, K3nhy6, S3nhy6, A4nhy6, I4nhy6, Q4nhy6, Y4nhy6;
wire G5nhy6, O5nhy6, W5nhy6, E6nhy6, M6nhy6, U6nhy6, C7nhy6, K7nhy6, S7nhy6, A8nhy6;
wire I8nhy6, Q8nhy6, Y8nhy6, G9nhy6, O9nhy6, W9nhy6, Eanhy6, Manhy6, Uanhy6, Cbnhy6;
wire Kbnhy6, Sbnhy6, Acnhy6, Icnhy6, Qcnhy6, Ycnhy6, Gdnhy6, Odnhy6, Wdnhy6, Eenhy6;
wire Menhy6, Uenhy6, Cfnhy6, Kfnhy6, Sfnhy6, Agnhy6, Ignhy6, Qgnhy6, Ygnhy6, Ghnhy6;
wire Ohnhy6, Whnhy6, Einhy6, Minhy6, Uinhy6, Cjnhy6, Kjnhy6, Sjnhy6, Aknhy6, Iknhy6;
wire Qknhy6, Yknhy6, Glnhy6, Olnhy6, Wlnhy6, Emnhy6, Mmnhy6, Umnhy6, Cnnhy6, Knnhy6;
wire Snnhy6, Aonhy6, Ionhy6, Qonhy6, Yonhy6, Gpnhy6, Opnhy6, Wpnhy6, Eqnhy6, Mqnhy6;
wire Uqnhy6, Crnhy6, Krnhy6, Srnhy6, Asnhy6, Isnhy6, Qsnhy6, Ysnhy6, Gtnhy6, Otnhy6;
wire Wtnhy6, Eunhy6, Munhy6, Uunhy6, Cvnhy6, Kvnhy6, Svnhy6, Awnhy6, Iwnhy6, Qwnhy6;
wire Ywnhy6, Gxnhy6, Oxnhy6, Wxnhy6, Eynhy6, Mynhy6, Uynhy6, Cznhy6, Kznhy6, Sznhy6;
wire A0ohy6, I0ohy6, Q0ohy6, Y0ohy6, G1ohy6, O1ohy6, W1ohy6, E2ohy6, M2ohy6, U2ohy6;
wire C3ohy6, K3ohy6, S3ohy6, A4ohy6, I4ohy6, Q4ohy6, Y4ohy6, G5ohy6, O5ohy6, W5ohy6;
wire E6ohy6, M6ohy6, U6ohy6, C7ohy6, K7ohy6, S7ohy6, A8ohy6, I8ohy6, Q8ohy6, Y8ohy6;
wire G9ohy6, O9ohy6, W9ohy6, Eaohy6, Maohy6, Uaohy6, Cbohy6, Kbohy6, Sbohy6, Acohy6;
wire Icohy6, Qcohy6, Ycohy6, Gdohy6, Odohy6, Wdohy6, Eeohy6, Meohy6, Ueohy6, Cfohy6;
wire Kfohy6, Sfohy6, Agohy6, Igohy6, Qgohy6, Ygohy6, Ghohy6, Ohohy6, Whohy6, Eiohy6;
wire Miohy6, Uiohy6, Cjohy6, Kjohy6, Sjohy6, Akohy6, Ikohy6, Qkohy6, Ykohy6, Glohy6;
wire Olohy6, Wlohy6, Emohy6, Mmohy6, Umohy6, Cnohy6, Knohy6, Snohy6, Aoohy6, Ioohy6;
wire Qoohy6, Yoohy6, Gpohy6, Opohy6, Wpohy6, Eqohy6, Mqohy6, Uqohy6, Crohy6, Krohy6;
wire Srohy6, Asohy6, Isohy6, Qsohy6, Ysohy6, Gtohy6, Otohy6, Wtohy6, Euohy6, Muohy6;
wire Uuohy6, Cvohy6, Kvohy6, Svohy6, Awohy6, Iwohy6, Qwohy6, Ywohy6, Gxohy6, Oxohy6;
wire Wxohy6, Eyohy6, Myohy6, Uyohy6, Czohy6, Kzohy6, Szohy6, A0phy6, I0phy6, Q0phy6;
wire Y0phy6, G1phy6, O1phy6, W1phy6, E2phy6, M2phy6, U2phy6, C3phy6, K3phy6, S3phy6;
wire A4phy6, I4phy6, Q4phy6, Y4phy6, G5phy6, O5phy6, W5phy6, E6phy6, M6phy6, U6phy6;
wire C7phy6, K7phy6, S7phy6, A8phy6, I8phy6, Q8phy6, Y8phy6, G9phy6, O9phy6, W9phy6;
wire Eaphy6, Maphy6, Uaphy6, Cbphy6, Kbphy6, Sbphy6, Acphy6, Icphy6, Qcphy6, Ycphy6;
wire Gdphy6, Odphy6, Wdphy6, Eephy6, Mephy6, Uephy6, Cfphy6, Kfphy6, Sfphy6, Agphy6;
wire Igphy6, Qgphy6, Ygphy6, Ghphy6, Ohphy6, Whphy6, Eiphy6, Miphy6, Uiphy6, Cjphy6;
wire Kjphy6, Sjphy6, Akphy6, Ikphy6, Qkphy6, Ykphy6, Glphy6, Olphy6, Wlphy6, Emphy6;
wire Mmphy6, Umphy6, Cnphy6, Knphy6, Snphy6, Aophy6, Iophy6, Qophy6, Yophy6, Gpphy6;
wire Opphy6, Wpphy6, Eqphy6, Mqphy6, Uqphy6, Crphy6, Krphy6, Srphy6, Asphy6, Isphy6;
wire Qsphy6, Ysphy6, Gtphy6, Otphy6, Wtphy6, Euphy6, Muphy6, Uuphy6, Cvphy6, Kvphy6;
wire Svphy6, Awphy6, Iwphy6, Qwphy6, Ywphy6, Gxphy6, Oxphy6, Wxphy6, Eyphy6, Myphy6;
wire Uyphy6, Czphy6, Kzphy6, Szphy6, A0qhy6, I0qhy6, Q0qhy6, Y0qhy6, G1qhy6, O1qhy6;
wire W1qhy6, E2qhy6, M2qhy6, U2qhy6, C3qhy6, K3qhy6, S3qhy6, A4qhy6, I4qhy6, Q4qhy6;
wire Y4qhy6, G5qhy6, O5qhy6, W5qhy6, E6qhy6, M6qhy6, U6qhy6, C7qhy6, K7qhy6, S7qhy6;
wire A8qhy6, I8qhy6, Q8qhy6, Y8qhy6, G9qhy6, O9qhy6, W9qhy6, Eaqhy6, Maqhy6, Uaqhy6;
wire Cbqhy6, Kbqhy6, Sbqhy6, Acqhy6, Icqhy6, Qcqhy6, Ycqhy6, Gdqhy6, Odqhy6, Wdqhy6;
wire Eeqhy6, Meqhy6, Ueqhy6, Cfqhy6, Kfqhy6, Sfqhy6, Agqhy6, Igqhy6, Qgqhy6, Ygqhy6;
wire Ghqhy6, Ohqhy6, Whqhy6, Eiqhy6, Miqhy6, Uiqhy6, Cjqhy6, Kjqhy6, Sjqhy6, Akqhy6;
wire Ikqhy6, Qkqhy6, Ykqhy6, Glqhy6, Olqhy6, Wlqhy6, Emqhy6, Mmqhy6, Umqhy6, Cnqhy6;
wire Knqhy6, Snqhy6, Aoqhy6, Ioqhy6, Qoqhy6, Yoqhy6, Gpqhy6, Opqhy6, Wpqhy6, Eqqhy6;
wire Mqqhy6, Uqqhy6, Crqhy6, Krqhy6, Srqhy6, Asqhy6, Isqhy6, Qsqhy6, Ysqhy6, Gtqhy6;
wire Otqhy6, Wtqhy6, Euqhy6, Muqhy6, Uuqhy6, Cvqhy6, Kvqhy6, Svqhy6, Awqhy6, Iwqhy6;
wire Qwqhy6, Ywqhy6, Gxqhy6, Oxqhy6, Wxqhy6, Eyqhy6, Myqhy6, Uyqhy6, Czqhy6, Kzqhy6;
wire Szqhy6, A0rhy6, I0rhy6, Q0rhy6, Y0rhy6, G1rhy6, O1rhy6, W1rhy6, E2rhy6, M2rhy6;
wire U2rhy6, C3rhy6, K3rhy6, S3rhy6, A4rhy6, I4rhy6, Q4rhy6, Y4rhy6, G5rhy6, O5rhy6;
wire W5rhy6, E6rhy6, M6rhy6, U6rhy6, C7rhy6, K7rhy6, S7rhy6, A8rhy6, I8rhy6, Q8rhy6;
wire Y8rhy6, G9rhy6, O9rhy6, W9rhy6, Earhy6, Marhy6, Uarhy6, Cbrhy6, Kbrhy6, Sbrhy6;
wire Acrhy6, Icrhy6, Qcrhy6, Ycrhy6, Gdrhy6, Odrhy6, Wdrhy6, Eerhy6, Merhy6, Uerhy6;
wire Cfrhy6, Kfrhy6, Sfrhy6, Agrhy6, Igrhy6, Qgrhy6, Ygrhy6, Ghrhy6, Ohrhy6, Whrhy6;
wire Eirhy6, Mirhy6, Uirhy6, Cjrhy6, Kjrhy6, Sjrhy6, Akrhy6, Ikrhy6, Qkrhy6, Ykrhy6;
wire Glrhy6, Olrhy6, Wlrhy6, Emrhy6, Mmrhy6, Umrhy6, Cnrhy6, Knrhy6, Snrhy6, Aorhy6;
wire Iorhy6, Qorhy6, Yorhy6, Gprhy6, Oprhy6, Wprhy6, Eqrhy6, Mqrhy6, Uqrhy6, Crrhy6;
wire Krrhy6, Srrhy6, Asrhy6, Isrhy6, Qsrhy6, Ysrhy6, Gtrhy6, Otrhy6, Wtrhy6, Eurhy6;
wire Murhy6, Uurhy6, Cvrhy6, Kvrhy6, Svrhy6, Awrhy6, Iwrhy6, Qwrhy6, Ywrhy6, Gxrhy6;
wire Oxrhy6, Wxrhy6, Eyrhy6, Myrhy6, Uyrhy6, Czrhy6, Kzrhy6, Szrhy6, A0shy6, I0shy6;
wire Q0shy6, Y0shy6, G1shy6, O1shy6, W1shy6, E2shy6, M2shy6, U2shy6, C3shy6, K3shy6;
wire S3shy6, A4shy6, I4shy6, Q4shy6, Y4shy6, G5shy6, O5shy6, W5shy6, E6shy6, M6shy6;
wire U6shy6, C7shy6, K7shy6, S7shy6, A8shy6, I8shy6, Q8shy6, Y8shy6, G9shy6, O9shy6;
wire W9shy6, Eashy6, Mashy6, Uashy6, Cbshy6, Kbshy6, Sbshy6, Acshy6, Icshy6, Qcshy6;
wire Ycshy6, Gdshy6, Odshy6, Wdshy6, Eeshy6, Meshy6, Ueshy6, Cfshy6, Kfshy6, Sfshy6;
wire Agshy6, Igshy6, Qgshy6, Ygshy6, Ghshy6, Ohshy6, Whshy6, Eishy6, Mishy6, Uishy6;
wire Cjshy6, Kjshy6, Sjshy6, Akshy6, Ikshy6, Qkshy6, Ykshy6, Glshy6, Olshy6, Wlshy6;
wire Emshy6, Mmshy6, Umshy6, Cnshy6, Knshy6, Snshy6, Aoshy6, Ioshy6, Qoshy6, Yoshy6;
wire Gpshy6, Opshy6, Wpshy6, Eqshy6, Mqshy6, Uqshy6, Crshy6, Krshy6, Srshy6, Asshy6;
wire Isshy6, Qsshy6, Ysshy6, Gtshy6, Otshy6, Wtshy6, Eushy6, Mushy6, Uushy6, Cvshy6;
wire Kvshy6, Svshy6, Awshy6, Iwshy6, Qwshy6, Ywshy6, Gxshy6, Oxshy6, Wxshy6, Eyshy6;
wire Myshy6, Uyshy6, Czshy6, Kzshy6, Szshy6, A0thy6, I0thy6, Q0thy6, Y0thy6, G1thy6;
wire O1thy6, W1thy6, E2thy6, M2thy6, U2thy6, C3thy6, K3thy6, S3thy6, A4thy6, I4thy6;
wire Q4thy6, Y4thy6, G5thy6, O5thy6, W5thy6, E6thy6, M6thy6, U6thy6, C7thy6, K7thy6;
wire S7thy6, A8thy6, I8thy6, Q8thy6, Y8thy6, G9thy6, O9thy6, W9thy6, Eathy6, Mathy6;
wire Uathy6, Cbthy6, Kbthy6, Sbthy6, Acthy6, Icthy6, Qcthy6, Ycthy6, Gdthy6, Odthy6;
wire Wdthy6, Eethy6, Methy6, Uethy6, Cfthy6, Kfthy6, Sfthy6, Agthy6, Igthy6, Qgthy6;
wire Ygthy6, Ghthy6, Ohthy6, Whthy6, Eithy6, Mithy6, Uithy6, Cjthy6, Kjthy6, Sjthy6;
wire Akthy6, Ikthy6, Qkthy6, Ykthy6, Glthy6, Olthy6, Wlthy6, Emthy6, Mmthy6, Umthy6;
wire Cnthy6, Knthy6, Snthy6, Aothy6, Iothy6, Qothy6, Yothy6, Gpthy6, Opthy6, Wpthy6;
wire Eqthy6, Mqthy6, Uqthy6, Crthy6, Krthy6, Srthy6, Asthy6, Isthy6, Qsthy6, Ysthy6;
wire Gtthy6, Otthy6, Wtthy6, Euthy6, Muthy6, Uuthy6, Cvthy6, Kvthy6, Svthy6, Awthy6;
wire Iwthy6, Qwthy6, Ywthy6, Gxthy6, Oxthy6, Wxthy6, Eythy6, Mythy6, Uythy6, Czthy6;
wire Kzthy6, Szthy6, A0uhy6, I0uhy6, Q0uhy6, Y0uhy6, G1uhy6, O1uhy6, W1uhy6, E2uhy6;
wire M2uhy6, U2uhy6, C3uhy6, K3uhy6, S3uhy6, A4uhy6, I4uhy6, Q4uhy6, Y4uhy6, G5uhy6;
wire O5uhy6, W5uhy6, E6uhy6, M6uhy6, U6uhy6, C7uhy6, K7uhy6, S7uhy6, A8uhy6, I8uhy6;
wire Q8uhy6, Y8uhy6, G9uhy6, O9uhy6, W9uhy6, Eauhy6, Mauhy6, Uauhy6, Cbuhy6, Kbuhy6;
wire Sbuhy6, Acuhy6, Icuhy6, Qcuhy6, Ycuhy6, Gduhy6, Oduhy6, Wduhy6, Eeuhy6, Meuhy6;
wire Ueuhy6, Cfuhy6, Kfuhy6, Sfuhy6, Aguhy6, Iguhy6, Qguhy6, Yguhy6, Ghuhy6, Ohuhy6;
wire Whuhy6, Eiuhy6, Miuhy6, Uiuhy6, Cjuhy6, Kjuhy6, Sjuhy6, Akuhy6, Ikuhy6, Qkuhy6;
wire Ykuhy6, Gluhy6, Oluhy6, Wluhy6, Emuhy6, Mmuhy6, Umuhy6, Cnuhy6, Knuhy6, Snuhy6;
wire Aouhy6, Iouhy6, Qouhy6, Youhy6, Gpuhy6, Opuhy6, Wpuhy6, Equhy6, Mquhy6, Uquhy6;
wire Cruhy6, Kruhy6, Sruhy6, Asuhy6, Isuhy6, Qsuhy6, Ysuhy6, Gtuhy6, Otuhy6, Wtuhy6;
wire Euuhy6, Muuhy6, Uuuhy6, Cvuhy6, Kvuhy6, Svuhy6, Awuhy6, Iwuhy6, Qwuhy6, Ywuhy6;
wire Gxuhy6, Oxuhy6, Wxuhy6, Eyuhy6, Myuhy6, Uyuhy6, Czuhy6, Kzuhy6, Szuhy6, A0vhy6;
wire I0vhy6, Q0vhy6, Y0vhy6, G1vhy6, O1vhy6, W1vhy6, E2vhy6, M2vhy6, U2vhy6, C3vhy6;
wire K3vhy6, S3vhy6, A4vhy6, I4vhy6, Q4vhy6, Y4vhy6, G5vhy6, O5vhy6, W5vhy6, E6vhy6;
wire M6vhy6, U6vhy6, C7vhy6, K7vhy6, S7vhy6, A8vhy6, I8vhy6, Q8vhy6, Y8vhy6, G9vhy6;
wire O9vhy6, W9vhy6, Eavhy6, Mavhy6, Uavhy6, Cbvhy6, Kbvhy6, Sbvhy6, Acvhy6, Icvhy6;
wire Qcvhy6, Ycvhy6, Gdvhy6, Odvhy6, Wdvhy6, Eevhy6, Mevhy6, Uevhy6, Cfvhy6, Kfvhy6;
wire Sfvhy6, Agvhy6, Igvhy6, Qgvhy6, Ygvhy6, Ghvhy6, Ohvhy6, Whvhy6, Eivhy6, Mivhy6;
wire Uivhy6, Cjvhy6, Kjvhy6, Sjvhy6, Akvhy6, Ikvhy6, Qkvhy6, Ykvhy6, Glvhy6, Olvhy6;
wire Wlvhy6, Emvhy6, Mmvhy6, Umvhy6, Cnvhy6, Knvhy6, Snvhy6, Aovhy6, Iovhy6, Qovhy6;
wire Yovhy6, Gpvhy6, Opvhy6, Wpvhy6, Eqvhy6, Mqvhy6, Uqvhy6, Crvhy6, Krvhy6, Srvhy6;
wire Asvhy6, Isvhy6, Qsvhy6, Ysvhy6, Gtvhy6, Otvhy6, Wtvhy6, Euvhy6, Muvhy6, Uuvhy6;
wire Cvvhy6, Kvvhy6, Svvhy6, Awvhy6, Iwvhy6, Qwvhy6, Ywvhy6, Gxvhy6, Oxvhy6, Wxvhy6;
wire Eyvhy6, Myvhy6, Uyvhy6, Czvhy6, Kzvhy6, Szvhy6, A0why6, I0why6, Q0why6, Y0why6;
wire G1why6, O1why6, W1why6, E2why6, M2why6, U2why6, C3why6, K3why6, S3why6, A4why6;
wire I4why6, Q4why6, Y4why6, G5why6, O5why6, W5why6, E6why6, M6why6, U6why6, C7why6;
wire K7why6, S7why6, A8why6, I8why6, Q8why6, Y8why6, G9why6, O9why6, W9why6, Eawhy6;
wire Mawhy6, Uawhy6, Cbwhy6, Kbwhy6, Sbwhy6, Acwhy6, Icwhy6, Qcwhy6, Ycwhy6, Gdwhy6;
wire Odwhy6, Wdwhy6, Eewhy6, Mewhy6, Uewhy6, Cfwhy6, Kfwhy6, Sfwhy6, Agwhy6, Igwhy6;
wire Qgwhy6, Ygwhy6, Ghwhy6, Ohwhy6, Whwhy6, Eiwhy6, Miwhy6, Uiwhy6, Cjwhy6, Kjwhy6;
wire Sjwhy6, Akwhy6, Ikwhy6, Qkwhy6, Ykwhy6, Glwhy6, Olwhy6, Wlwhy6, Emwhy6, Mmwhy6;
wire Umwhy6, Cnwhy6, Knwhy6, Snwhy6, Aowhy6, Iowhy6, Qowhy6, Yowhy6, Gpwhy6, Opwhy6;
wire Wpwhy6, Eqwhy6, Mqwhy6, Uqwhy6, Crwhy6, Krwhy6, Srwhy6, Aswhy6, Iswhy6, Qswhy6;
wire Yswhy6, Gtwhy6, Otwhy6, Wtwhy6, Euwhy6, Muwhy6, Uuwhy6, Cvwhy6, Kvwhy6, Svwhy6;
wire Awwhy6, Iwwhy6, Qwwhy6, Ywwhy6, Gxwhy6, Oxwhy6, Wxwhy6, Eywhy6, Mywhy6, Uywhy6;
wire Czwhy6, Kzwhy6, Szwhy6, A0xhy6, I0xhy6, Q0xhy6, Y0xhy6, G1xhy6, O1xhy6, W1xhy6;
wire E2xhy6, M2xhy6, U2xhy6, C3xhy6, K3xhy6, S3xhy6, A4xhy6, I4xhy6, Q4xhy6, Y4xhy6;
wire G5xhy6, O5xhy6, W5xhy6, E6xhy6, M6xhy6, U6xhy6, C7xhy6, K7xhy6, S7xhy6, A8xhy6;
wire I8xhy6, Q8xhy6, Y8xhy6, G9xhy6, O9xhy6, W9xhy6, Eaxhy6, Maxhy6, Uaxhy6, Cbxhy6;
wire Kbxhy6, Sbxhy6, Acxhy6, Icxhy6, Qcxhy6, Ycxhy6, Gdxhy6, Odxhy6, Wdxhy6, Eexhy6;
wire Mexhy6, Uexhy6, Cfxhy6, Kfxhy6, Sfxhy6, Agxhy6, Igxhy6, Qgxhy6, Ygxhy6, Ghxhy6;
wire Ohxhy6, Whxhy6, Eixhy6, Mixhy6, Uixhy6, Cjxhy6, Kjxhy6, Sjxhy6, Akxhy6, Ikxhy6;
wire Qkxhy6, Ykxhy6, Glxhy6, Olxhy6, Wlxhy6, Emxhy6, Mmxhy6, Umxhy6, Cnxhy6, Knxhy6;
wire Snxhy6, Aoxhy6, Ioxhy6, Qoxhy6, Yoxhy6, Gpxhy6, Opxhy6, Wpxhy6, Eqxhy6, Mqxhy6;
wire Uqxhy6, Crxhy6, Krxhy6, Srxhy6, Asxhy6, Isxhy6, Qsxhy6, Ysxhy6, Gtxhy6, Otxhy6;
wire Wtxhy6, Euxhy6, Muxhy6, Uuxhy6, Cvxhy6, Kvxhy6, Svxhy6, Awxhy6, Iwxhy6, Qwxhy6;
wire Ywxhy6, Gxxhy6, Oxxhy6, Wxxhy6, Eyxhy6, Myxhy6, Uyxhy6, Czxhy6, Kzxhy6, Szxhy6;
wire A0yhy6, I0yhy6, Q0yhy6, Y0yhy6, G1yhy6, O1yhy6, W1yhy6, E2yhy6, M2yhy6, U2yhy6;
wire C3yhy6, K3yhy6, S3yhy6, A4yhy6, I4yhy6, Q4yhy6, Y4yhy6, G5yhy6, O5yhy6, W5yhy6;
wire E6yhy6, M6yhy6, U6yhy6, C7yhy6, K7yhy6, S7yhy6, A8yhy6, I8yhy6, Q8yhy6, Y8yhy6;
wire G9yhy6, O9yhy6, W9yhy6, Eayhy6, Mayhy6, Uayhy6, Cbyhy6, Kbyhy6, Sbyhy6, Acyhy6;
wire Icyhy6, Qcyhy6, Ycyhy6, Gdyhy6, Odyhy6, Wdyhy6, Eeyhy6, Meyhy6, Ueyhy6, Cfyhy6;
wire Kfyhy6, Sfyhy6, Agyhy6, Igyhy6, Qgyhy6, Ygyhy6, Ghyhy6, Ohyhy6, Whyhy6, Eiyhy6;
wire Miyhy6, Uiyhy6, Cjyhy6, Kjyhy6, Sjyhy6, Akyhy6, Ikyhy6, Qkyhy6, Ykyhy6, Glyhy6;
wire Olyhy6, Wlyhy6, Emyhy6, Mmyhy6, Umyhy6, Cnyhy6, Knyhy6, Snyhy6, Aoyhy6, Ioyhy6;
wire Qoyhy6, Yoyhy6, Gpyhy6, Opyhy6, Wpyhy6, Eqyhy6, Mqyhy6, Uqyhy6, Cryhy6, Kryhy6;
wire Sryhy6, Asyhy6, Isyhy6, Qsyhy6, Ysyhy6, Gtyhy6, Otyhy6, Wtyhy6, Euyhy6, Muyhy6;
wire Uuyhy6, Cvyhy6, Kvyhy6, Svyhy6, Awyhy6, Iwyhy6, Qwyhy6, Ywyhy6, Gxyhy6, Oxyhy6;
wire Wxyhy6, Eyyhy6, Myyhy6, Uyyhy6, Czyhy6, Kzyhy6, Szyhy6, A0zhy6, I0zhy6, Q0zhy6;
wire Y0zhy6, G1zhy6, O1zhy6, W1zhy6, E2zhy6, M2zhy6, U2zhy6, C3zhy6, K3zhy6, S3zhy6;
wire A4zhy6, I4zhy6, Q4zhy6, Y4zhy6, G5zhy6, O5zhy6, W5zhy6, E6zhy6, M6zhy6, U6zhy6;
wire C7zhy6, K7zhy6, S7zhy6, A8zhy6, I8zhy6, Q8zhy6, Y8zhy6, G9zhy6, O9zhy6, W9zhy6;
wire Eazhy6, Mazhy6, Uazhy6, Cbzhy6, Kbzhy6, Sbzhy6, Aczhy6, Iczhy6, Qczhy6, Yczhy6;
wire Gdzhy6, Odzhy6, Wdzhy6, Eezhy6, Mezhy6, Uezhy6, Cfzhy6, Kfzhy6, Sfzhy6, Agzhy6;
wire Igzhy6, Qgzhy6, Ygzhy6, Ghzhy6, Ohzhy6, Whzhy6, Eizhy6, Mizhy6, Uizhy6, Cjzhy6;
wire Kjzhy6, Sjzhy6, Akzhy6, Ikzhy6, Qkzhy6, Ykzhy6, Glzhy6, Olzhy6, Wlzhy6, Emzhy6;
wire Mmzhy6, Umzhy6, Cnzhy6, Knzhy6, Snzhy6, Aozhy6, Iozhy6, Qozhy6, Yozhy6, Gpzhy6;
wire Opzhy6, Wpzhy6, Eqzhy6, Mqzhy6, Uqzhy6, Crzhy6, Krzhy6, Srzhy6, Aszhy6, Iszhy6;
wire Qszhy6, Yszhy6, Gtzhy6, Otzhy6, Wtzhy6, Euzhy6, Muzhy6, Uuzhy6, Cvzhy6, Kvzhy6;
wire Svzhy6, Awzhy6, Iwzhy6, Qwzhy6, Ywzhy6, Gxzhy6, Oxzhy6, Wxzhy6, Eyzhy6, Myzhy6;
wire Uyzhy6, Czzhy6, Kzzhy6, Szzhy6, A00iy6, I00iy6, Q00iy6, Y00iy6, G10iy6, O10iy6;
wire W10iy6, E20iy6, M20iy6, U20iy6, C30iy6, K30iy6, S30iy6, A40iy6, I40iy6, Q40iy6;
wire Y40iy6, G50iy6, O50iy6, W50iy6, E60iy6, M60iy6, U60iy6, C70iy6, K70iy6, S70iy6;
wire A80iy6, I80iy6, Q80iy6, Y80iy6, G90iy6, O90iy6, W90iy6, Ea0iy6, Ma0iy6, Ua0iy6;
wire Cb0iy6, Kb0iy6, Sb0iy6, Ac0iy6, Ic0iy6, Qc0iy6, Yc0iy6, Gd0iy6, Od0iy6, Wd0iy6;
wire Ee0iy6, Me0iy6, Ue0iy6, Cf0iy6, Kf0iy6, Sf0iy6, Ag0iy6, Ig0iy6, Qg0iy6, Yg0iy6;
wire Gh0iy6, Oh0iy6, Wh0iy6, Ei0iy6, Mi0iy6, Ui0iy6, Cj0iy6, Kj0iy6, Sj0iy6, Ak0iy6;
wire Ik0iy6, Qk0iy6, Yk0iy6, Gl0iy6, Ol0iy6, Wl0iy6, Em0iy6, Mm0iy6, Um0iy6, Cn0iy6;
wire Kn0iy6, Sn0iy6, Ao0iy6, Io0iy6, Qo0iy6, Yo0iy6, Gp0iy6, Op0iy6, Wp0iy6, Eq0iy6;
wire Mq0iy6, Uq0iy6, Cr0iy6, Kr0iy6, Sr0iy6, As0iy6, Is0iy6, Qs0iy6, Ys0iy6, Gt0iy6;
wire Ot0iy6, Wt0iy6, Eu0iy6, Mu0iy6, Uu0iy6, Cv0iy6, Kv0iy6, Sv0iy6, Aw0iy6, Iw0iy6;
wire Qw0iy6, Yw0iy6, Gx0iy6, Ox0iy6, Wx0iy6, Ey0iy6, My0iy6, Uy0iy6, Cz0iy6, Kz0iy6;
wire Sz0iy6, A01iy6, I01iy6, Q01iy6, Y01iy6, G11iy6, O11iy6, W11iy6, E21iy6, M21iy6;
wire U21iy6, C31iy6, K31iy6, S31iy6, A41iy6, I41iy6, Q41iy6, Y41iy6, G51iy6, O51iy6;
wire W51iy6, E61iy6, M61iy6, U61iy6, C71iy6, K71iy6, S71iy6, A81iy6, I81iy6, Q81iy6;
wire Y81iy6, G91iy6, O91iy6, W91iy6, Ea1iy6, Ma1iy6, Ua1iy6, Cb1iy6, Kb1iy6, Sb1iy6;
wire Ac1iy6, Ic1iy6, Qc1iy6, Yc1iy6, Gd1iy6, Od1iy6, Wd1iy6, Ee1iy6, Me1iy6, Ue1iy6;
wire Cf1iy6, Kf1iy6, Sf1iy6, Ag1iy6, Ig1iy6, Qg1iy6, Yg1iy6, Gh1iy6, Oh1iy6, Wh1iy6;
wire Ei1iy6, Mi1iy6, Ui1iy6, Cj1iy6, Kj1iy6, Sj1iy6, Ak1iy6, Ik1iy6, Qk1iy6, Yk1iy6;
wire Gl1iy6, Ol1iy6, Wl1iy6, Em1iy6, Mm1iy6, Um1iy6, Cn1iy6, Kn1iy6, Sn1iy6, Ao1iy6;
wire Io1iy6, Qo1iy6, Yo1iy6, Gp1iy6, Op1iy6, Wp1iy6, Eq1iy6, Mq1iy6, Uq1iy6, Cr1iy6;
wire Kr1iy6, Sr1iy6, As1iy6, Is1iy6, Qs1iy6, Ys1iy6, Gt1iy6, Ot1iy6, Wt1iy6, Eu1iy6;
wire Mu1iy6, Uu1iy6, Cv1iy6, Kv1iy6, Sv1iy6, Aw1iy6, Iw1iy6, Qw1iy6, Yw1iy6, Gx1iy6;
wire Ox1iy6, Wx1iy6, Ey1iy6, My1iy6, Uy1iy6, Cz1iy6, Kz1iy6, Sz1iy6, A02iy6, I02iy6;
wire Q02iy6, Y02iy6, G12iy6, O12iy6, W12iy6, E22iy6, M22iy6, U22iy6, C32iy6, K32iy6;
wire S32iy6, A42iy6, I42iy6, Q42iy6, Y42iy6, G52iy6, O52iy6, W52iy6, E62iy6, M62iy6;
wire U62iy6, C72iy6, K72iy6, S72iy6, A82iy6, I82iy6, Q82iy6, Y82iy6, G92iy6, O92iy6;
wire W92iy6, Ea2iy6, Ma2iy6, Ua2iy6, Cb2iy6, Kb2iy6, Sb2iy6, Ac2iy6, Ic2iy6, Qc2iy6;
wire Yc2iy6, Gd2iy6, Od2iy6, Wd2iy6, Ee2iy6, Me2iy6, Ue2iy6, Cf2iy6, Kf2iy6, Sf2iy6;
wire Ag2iy6, Ig2iy6, Qg2iy6, Yg2iy6, Gh2iy6, Oh2iy6, Wh2iy6, Ei2iy6, Mi2iy6, Ui2iy6;
wire Cj2iy6, Kj2iy6, Sj2iy6, Ak2iy6, Ik2iy6, Qk2iy6, Yk2iy6, Gl2iy6, Ol2iy6, Wl2iy6;
wire Em2iy6, Mm2iy6, Um2iy6, Cn2iy6, Kn2iy6, Sn2iy6, Ao2iy6, Io2iy6, Qo2iy6, Yo2iy6;
wire Gp2iy6, Op2iy6, Wp2iy6, Eq2iy6, Mq2iy6, Uq2iy6, Cr2iy6, Kr2iy6, Sr2iy6, As2iy6;
wire Is2iy6, Qs2iy6, Ys2iy6, Gt2iy6, Ot2iy6, Wt2iy6, Eu2iy6, Mu2iy6, Uu2iy6, Cv2iy6;
wire Kv2iy6, Sv2iy6, Aw2iy6, Iw2iy6, Qw2iy6, Yw2iy6, Gx2iy6, Ox2iy6, Wx2iy6, Ey2iy6;
wire My2iy6, Uy2iy6, Cz2iy6, Kz2iy6, Sz2iy6, A03iy6, I03iy6, Q03iy6, Y03iy6, G13iy6;
wire O13iy6, W13iy6, E23iy6, M23iy6, U23iy6, C33iy6, K33iy6, S33iy6, A43iy6, I43iy6;
wire Q43iy6, Y43iy6, G53iy6, O53iy6, W53iy6, E63iy6, M63iy6, U63iy6, C73iy6, K73iy6;
wire S73iy6, A83iy6, I83iy6, Q83iy6, Y83iy6, G93iy6, O93iy6, W93iy6, Ea3iy6, Ma3iy6;
wire Ua3iy6, Cb3iy6, Kb3iy6, Sb3iy6, Ac3iy6, Ic3iy6, Qc3iy6, Yc3iy6, Gd3iy6, Od3iy6;
wire Wd3iy6, Ee3iy6, Me3iy6, Ue3iy6, Cf3iy6, Kf3iy6, Sf3iy6, Ag3iy6, Ig3iy6, Qg3iy6;
wire Yg3iy6, Gh3iy6, Oh3iy6, Wh3iy6, Ei3iy6, Mi3iy6, Ui3iy6, Cj3iy6, Kj3iy6, Sj3iy6;
wire Ak3iy6, Ik3iy6, Qk3iy6, Yk3iy6, Gl3iy6, Ol3iy6, Wl3iy6, Em3iy6, Mm3iy6, Um3iy6;
wire Cn3iy6, Kn3iy6, Sn3iy6, Ao3iy6, Io3iy6, Qo3iy6, Yo3iy6, Gp3iy6, Op3iy6, Wp3iy6;
wire Eq3iy6, Mq3iy6, Uq3iy6, Cr3iy6, Kr3iy6, Sr3iy6, As3iy6, Is3iy6, Qs3iy6, Ys3iy6;
wire Gt3iy6, Ot3iy6, Wt3iy6, Eu3iy6, Mu3iy6, Uu3iy6, Cv3iy6, Kv3iy6, Sv3iy6, Aw3iy6;
wire Iw3iy6, Qw3iy6, Yw3iy6, Gx3iy6, Ox3iy6, Wx3iy6, Ey3iy6, My3iy6, Uy3iy6, Cz3iy6;
wire Kz3iy6, Sz3iy6, A04iy6, I04iy6, Q04iy6, Y04iy6, G14iy6, O14iy6, W14iy6, E24iy6;
wire M24iy6, U24iy6, C34iy6, K34iy6, S34iy6, A44iy6, I44iy6, Q44iy6, Y44iy6, G54iy6;
wire O54iy6, W54iy6, E64iy6, M64iy6, U64iy6, C74iy6, K74iy6, S74iy6, A84iy6, I84iy6;
wire Q84iy6, Y84iy6, G94iy6, O94iy6, W94iy6, Ea4iy6, Ma4iy6, Ua4iy6, Cb4iy6, Kb4iy6;
wire Sb4iy6, Ac4iy6, Ic4iy6, Qc4iy6, Yc4iy6, Gd4iy6, Od4iy6, Wd4iy6, Ee4iy6, Me4iy6;
wire Ue4iy6, Cf4iy6, Kf4iy6, Sf4iy6, Ag4iy6, Ig4iy6, Qg4iy6, Yg4iy6, Gh4iy6, Oh4iy6;
wire Wh4iy6, Ei4iy6, Mi4iy6, Ui4iy6, Cj4iy6, Kj4iy6, Sj4iy6, Ak4iy6, Ik4iy6, Qk4iy6;
wire Yk4iy6, Gl4iy6, Ol4iy6, Wl4iy6, Em4iy6, Mm4iy6, Um4iy6, Cn4iy6, Kn4iy6, Sn4iy6;
wire Ao4iy6, Io4iy6, Qo4iy6, Yo4iy6, Gp4iy6, Op4iy6, Wp4iy6, Eq4iy6, Mq4iy6, Uq4iy6;
wire Cr4iy6, Kr4iy6, Sr4iy6, As4iy6, Is4iy6, Qs4iy6, Ys4iy6, Gt4iy6, Ot4iy6, Wt4iy6;
wire Eu4iy6, Mu4iy6, Uu4iy6, Cv4iy6, Kv4iy6, Sv4iy6, Aw4iy6, Iw4iy6, Qw4iy6, Yw4iy6;
wire Gx4iy6, Ox4iy6, Wx4iy6, Ey4iy6, My4iy6, Uy4iy6, Cz4iy6, Kz4iy6, Sz4iy6, A05iy6;
wire I05iy6, Q05iy6, Y05iy6, G15iy6, O15iy6, W15iy6, E25iy6, M25iy6, U25iy6, C35iy6;
wire K35iy6, S35iy6, A45iy6, I45iy6, Q45iy6, Y45iy6, G55iy6, O55iy6, W55iy6, E65iy6;
wire M65iy6, U65iy6, C75iy6, K75iy6, S75iy6, A85iy6, I85iy6, Q85iy6, Y85iy6, G95iy6;
wire O95iy6, W95iy6, Ea5iy6, Ma5iy6, Ua5iy6, Cb5iy6, Kb5iy6, Sb5iy6, Ac5iy6, Ic5iy6;
wire Qc5iy6, Yc5iy6, Gd5iy6, Od5iy6, Wd5iy6, Ee5iy6, Me5iy6, Ue5iy6, Cf5iy6, Kf5iy6;
wire Sf5iy6, Ag5iy6, Ig5iy6, Qg5iy6, Yg5iy6, Gh5iy6, Oh5iy6, Wh5iy6, Ei5iy6, Mi5iy6;
wire Ui5iy6, Cj5iy6, Kj5iy6, Sj5iy6, Ak5iy6, Ik5iy6, Qk5iy6, Yk5iy6, Gl5iy6, Ol5iy6;
wire Wl5iy6, Em5iy6, Mm5iy6, Um5iy6, Cn5iy6, Kn5iy6, Sn5iy6, Ao5iy6, Io5iy6, Qo5iy6;
wire Yo5iy6, Gp5iy6, Op5iy6, Wp5iy6, Eq5iy6, Mq5iy6, Uq5iy6, Cr5iy6, Kr5iy6, Sr5iy6;
wire As5iy6, Is5iy6, Qs5iy6, Ys5iy6, Gt5iy6, Ot5iy6, Wt5iy6, Eu5iy6, Mu5iy6, Uu5iy6;
wire Cv5iy6, Kv5iy6, Sv5iy6, Aw5iy6, Iw5iy6, Qw5iy6, Yw5iy6, Gx5iy6, Ox5iy6, Wx5iy6;
wire Ey5iy6, My5iy6, Uy5iy6, Cz5iy6, Kz5iy6, Sz5iy6, A06iy6, I06iy6, Q06iy6, Y06iy6;
wire G16iy6, O16iy6, W16iy6, E26iy6, M26iy6, U26iy6, C36iy6, K36iy6, S36iy6, A46iy6;
wire I46iy6, Q46iy6, Y46iy6, G56iy6, O56iy6, W56iy6, E66iy6, M66iy6, U66iy6, C76iy6;
wire K76iy6, S76iy6, A86iy6, I86iy6, Q86iy6, Y86iy6, G96iy6, O96iy6, W96iy6, Ea6iy6;
wire Ma6iy6, Ua6iy6, Cb6iy6, Kb6iy6, Sb6iy6, Ac6iy6, Ic6iy6, Qc6iy6, Yc6iy6, Gd6iy6;
wire Od6iy6, Wd6iy6, Ee6iy6, Me6iy6, Ue6iy6, Cf6iy6, Kf6iy6, Sf6iy6, Ag6iy6, Ig6iy6;
wire Qg6iy6, Yg6iy6, Gh6iy6, Oh6iy6, Wh6iy6, Ei6iy6, Mi6iy6, Ui6iy6, Cj6iy6, Kj6iy6;
wire Sj6iy6, Ak6iy6, Ik6iy6, Qk6iy6, Yk6iy6, Gl6iy6, Ol6iy6, Wl6iy6, Em6iy6, Mm6iy6;
wire Um6iy6, Cn6iy6, Kn6iy6, Sn6iy6, Ao6iy6, Io6iy6, Qo6iy6, Yo6iy6, Gp6iy6, Op6iy6;
wire Wp6iy6, Eq6iy6, Mq6iy6, Uq6iy6, Cr6iy6, Kr6iy6, Sr6iy6, As6iy6, Is6iy6, Qs6iy6;
wire Ys6iy6, Gt6iy6, Ot6iy6, Wt6iy6, Eu6iy6, Mu6iy6, Uu6iy6, Cv6iy6, Kv6iy6, Sv6iy6;
wire Aw6iy6, Iw6iy6, Qw6iy6, Yw6iy6, Gx6iy6, Ox6iy6, Wx6iy6, Ey6iy6, My6iy6, Uy6iy6;
wire Cz6iy6, Kz6iy6, Sz6iy6, A07iy6, I07iy6, Q07iy6, Y07iy6, G17iy6, O17iy6, W17iy6;
wire E27iy6, M27iy6, U27iy6, C37iy6, K37iy6, S37iy6, A47iy6, I47iy6, Q47iy6, Y47iy6;
wire G57iy6, O57iy6, W57iy6, E67iy6, M67iy6, U67iy6, C77iy6, K77iy6, S77iy6, A87iy6;
wire I87iy6, Q87iy6, Y87iy6, G97iy6, O97iy6, W97iy6, Ea7iy6, Ma7iy6, Ua7iy6, Cb7iy6;
wire Kb7iy6, Sb7iy6, Ac7iy6, Ic7iy6, Qc7iy6, Yc7iy6, Gd7iy6, Od7iy6, Wd7iy6, Ee7iy6;
wire Me7iy6, Ue7iy6, Cf7iy6, Kf7iy6, Sf7iy6, Ag7iy6, Ig7iy6, Qg7iy6, Yg7iy6, Gh7iy6;
wire Oh7iy6, Wh7iy6, Ei7iy6, Mi7iy6, Ui7iy6, Cj7iy6, Kj7iy6, Sj7iy6, Ak7iy6, Ik7iy6;
wire Qk7iy6, Yk7iy6, Gl7iy6, Ol7iy6, Wl7iy6, Em7iy6, Mm7iy6, Um7iy6, Cn7iy6, Kn7iy6;
wire Sn7iy6, Ao7iy6, Io7iy6, Qo7iy6, Yo7iy6, Gp7iy6, Op7iy6, Wp7iy6, Eq7iy6, Mq7iy6;
wire Uq7iy6, Cr7iy6, Kr7iy6, Sr7iy6, As7iy6, Is7iy6, Qs7iy6, Ys7iy6, Gt7iy6, Ot7iy6;
wire Wt7iy6, Eu7iy6, Mu7iy6, Uu7iy6, Cv7iy6, Kv7iy6, Sv7iy6, Aw7iy6, Iw7iy6, Qw7iy6;
wire Yw7iy6, Gx7iy6, Ox7iy6, Wx7iy6, Ey7iy6, My7iy6, Uy7iy6, Cz7iy6, Kz7iy6, Sz7iy6;
wire A08iy6, I08iy6, Q08iy6, Y08iy6, G18iy6, O18iy6, W18iy6, E28iy6, M28iy6, U28iy6;
wire C38iy6, K38iy6, S38iy6, A48iy6, I48iy6, Q48iy6, Y48iy6, G58iy6, O58iy6, W58iy6;
wire E68iy6, M68iy6, U68iy6, C78iy6, K78iy6, S78iy6, A88iy6, I88iy6, Q88iy6, Y88iy6;
wire G98iy6, O98iy6, W98iy6, Ea8iy6, Ma8iy6, Ua8iy6, Cb8iy6, Kb8iy6, Sb8iy6, Ac8iy6;
wire Ic8iy6, Qc8iy6, Yc8iy6, Gd8iy6, Od8iy6, Wd8iy6, Ee8iy6, Me8iy6, Ue8iy6, Cf8iy6;
wire Kf8iy6, Sf8iy6, Ag8iy6, Ig8iy6, Qg8iy6, Yg8iy6, Gh8iy6, Oh8iy6, Wh8iy6, Ei8iy6;
wire Mi8iy6, Ui8iy6, Cj8iy6, Kj8iy6, Sj8iy6, Ak8iy6, Ik8iy6, Qk8iy6, Yk8iy6, Gl8iy6;
wire Ol8iy6, Wl8iy6, Em8iy6, Mm8iy6, Um8iy6, Cn8iy6, Kn8iy6, Sn8iy6, Ao8iy6, Io8iy6;
wire Qo8iy6, Yo8iy6, Gp8iy6, Op8iy6, Wp8iy6, Eq8iy6, Mq8iy6, Uq8iy6, Cr8iy6, Kr8iy6;
wire Sr8iy6, As8iy6, Is8iy6, Qs8iy6, Ys8iy6, Gt8iy6, Ot8iy6, Wt8iy6, Eu8iy6, Mu8iy6;
wire Uu8iy6, Cv8iy6, Kv8iy6, Sv8iy6, Aw8iy6, Iw8iy6, Qw8iy6, Yw8iy6, Gx8iy6, Ox8iy6;
wire Wx8iy6, Ey8iy6, My8iy6, Uy8iy6, Cz8iy6, Kz8iy6, Sz8iy6, A09iy6, I09iy6, Q09iy6;
wire Y09iy6, G19iy6, O19iy6, W19iy6, E29iy6, M29iy6, U29iy6, C39iy6, K39iy6, S39iy6;
wire A49iy6, I49iy6, Q49iy6, Y49iy6, G59iy6, O59iy6, W59iy6, E69iy6, M69iy6, U69iy6;
wire C79iy6, K79iy6, S79iy6, A89iy6, I89iy6, Q89iy6, Y89iy6, G99iy6, O99iy6, W99iy6;
wire Ea9iy6, Ma9iy6, Ua9iy6, Cb9iy6, Kb9iy6, Sb9iy6, Ac9iy6, Ic9iy6, Qc9iy6, Yc9iy6;
wire Gd9iy6, Od9iy6, Wd9iy6, Ee9iy6, Me9iy6, Ue9iy6, Cf9iy6, Kf9iy6, Sf9iy6, Ag9iy6;
wire Ig9iy6, Qg9iy6, Yg9iy6, Gh9iy6, Oh9iy6, Wh9iy6, Ei9iy6, Mi9iy6, Ui9iy6, Cj9iy6;
wire Kj9iy6, Sj9iy6, Ak9iy6, Ik9iy6, Qk9iy6, Yk9iy6, Gl9iy6, Ol9iy6, Wl9iy6, Em9iy6;
wire Mm9iy6, Um9iy6, Cn9iy6, Kn9iy6, Sn9iy6, Ao9iy6, Io9iy6, Qo9iy6, Yo9iy6, Gp9iy6;
wire Op9iy6, Wp9iy6, Eq9iy6, Mq9iy6, Uq9iy6, Cr9iy6, Kr9iy6, Sr9iy6, As9iy6, Is9iy6;
wire Qs9iy6, Ys9iy6, Gt9iy6, Ot9iy6, Wt9iy6, Eu9iy6, Mu9iy6, Uu9iy6, Cv9iy6, Kv9iy6;
wire Sv9iy6, Aw9iy6, Iw9iy6, Qw9iy6, Yw9iy6, Gx9iy6, Ox9iy6, Wx9iy6, Ey9iy6, My9iy6;
wire Uy9iy6, Cz9iy6, Kz9iy6, Sz9iy6, A0aiy6, I0aiy6, Q0aiy6, Y0aiy6, G1aiy6, O1aiy6;
wire W1aiy6, E2aiy6, M2aiy6, U2aiy6, C3aiy6, K3aiy6, S3aiy6, A4aiy6, I4aiy6, Q4aiy6;
wire Y4aiy6, G5aiy6, O5aiy6, W5aiy6, E6aiy6, M6aiy6, U6aiy6, C7aiy6, K7aiy6, S7aiy6;
wire A8aiy6, I8aiy6, Q8aiy6, Y8aiy6, G9aiy6, O9aiy6, W9aiy6, Eaaiy6, Maaiy6, Uaaiy6;
wire Cbaiy6, Kbaiy6, Sbaiy6, Acaiy6, Icaiy6, Qcaiy6, Ycaiy6, Gdaiy6, Odaiy6, Wdaiy6;
wire Eeaiy6, Meaiy6, Ueaiy6, Cfaiy6, Kfaiy6, Sfaiy6, Agaiy6, Igaiy6, Qgaiy6, Ygaiy6;
wire Ghaiy6, Ohaiy6, Whaiy6, Eiaiy6, Miaiy6, Uiaiy6, Cjaiy6, Kjaiy6, Sjaiy6, Akaiy6;
wire Ikaiy6, Qkaiy6, Ykaiy6, Glaiy6, Olaiy6, Wlaiy6, Emaiy6, Mmaiy6, Umaiy6, Cnaiy6;
wire Knaiy6, Snaiy6, Aoaiy6, Ioaiy6, Qoaiy6, Yoaiy6, Gpaiy6, Opaiy6, Wpaiy6, Eqaiy6;
wire Mqaiy6, Uqaiy6, Craiy6, Kraiy6, Sraiy6, Asaiy6, Isaiy6, Qsaiy6, Ysaiy6, Gtaiy6;
wire Otaiy6, Wtaiy6, Euaiy6, Muaiy6, Uuaiy6, Cvaiy6, Kvaiy6, Svaiy6, Awaiy6, Iwaiy6;
wire Qwaiy6, Ywaiy6, Gxaiy6, Oxaiy6, Wxaiy6, Eyaiy6, Myaiy6, Uyaiy6, Czaiy6, Kzaiy6;
wire Szaiy6, A0biy6, I0biy6, Q0biy6, Y0biy6, G1biy6, O1biy6, W1biy6, E2biy6, M2biy6;
wire U2biy6, C3biy6, K3biy6, S3biy6, A4biy6, I4biy6, Q4biy6, Y4biy6, G5biy6, O5biy6;
wire W5biy6, E6biy6, M6biy6, U6biy6, C7biy6, K7biy6, S7biy6, A8biy6, I8biy6, Q8biy6;
wire Y8biy6, G9biy6, O9biy6, W9biy6, Eabiy6, Mabiy6, Uabiy6, Cbbiy6, Kbbiy6, Sbbiy6;
wire Acbiy6, Icbiy6, Qcbiy6, Ycbiy6, Gdbiy6, Odbiy6, Wdbiy6, Eebiy6, Mebiy6, Uebiy6;
wire Cfbiy6, Kfbiy6, Sfbiy6, Agbiy6, Igbiy6, Qgbiy6, Ygbiy6, Ghbiy6, Ohbiy6, Whbiy6;
wire Eibiy6, Mibiy6, Uibiy6, Cjbiy6, Kjbiy6, Sjbiy6, Akbiy6, Ikbiy6, Qkbiy6, Ykbiy6;
wire Glbiy6, Olbiy6, Wlbiy6, Embiy6, Mmbiy6, Umbiy6, Cnbiy6, Knbiy6, Snbiy6, Aobiy6;
wire Iobiy6, Qobiy6, Yobiy6, Gpbiy6, Opbiy6, Wpbiy6, Eqbiy6, Mqbiy6, Uqbiy6, Crbiy6;
wire Krbiy6, Srbiy6, Asbiy6, Isbiy6, Qsbiy6, Ysbiy6, Gtbiy6, Otbiy6, Wtbiy6, Eubiy6;
wire Mubiy6, Uubiy6, Cvbiy6, Kvbiy6, Svbiy6, Awbiy6, Iwbiy6, Qwbiy6, Ywbiy6, Gxbiy6;
wire Oxbiy6, Wxbiy6, Eybiy6, Mybiy6, Uybiy6, Czbiy6, Kzbiy6, Szbiy6, A0ciy6, I0ciy6;
wire Q0ciy6, Y0ciy6, G1ciy6, O1ciy6, W1ciy6, E2ciy6, M2ciy6, U2ciy6, C3ciy6, K3ciy6;
wire S3ciy6, A4ciy6, I4ciy6, Q4ciy6, Y4ciy6, G5ciy6, O5ciy6, W5ciy6, E6ciy6, M6ciy6;
wire U6ciy6, C7ciy6, K7ciy6, S7ciy6, A8ciy6, I8ciy6, Q8ciy6, Y8ciy6, G9ciy6, O9ciy6;
wire W9ciy6, Eaciy6, Maciy6, Uaciy6, Cbciy6, Kbciy6, Sbciy6, Acciy6, Icciy6, Qcciy6;
wire Ycciy6, Gdciy6, Odciy6, Wdciy6, Eeciy6, Meciy6, Ueciy6, Cfciy6, Kfciy6, Sfciy6;
wire Agciy6, Igciy6, Qgciy6, Ygciy6, Ghciy6, Ohciy6, Whciy6, Eiciy6, Miciy6, Uiciy6;
wire Cjciy6, Kjciy6, Sjciy6, Akciy6, Ikciy6, Qkciy6, Ykciy6, Glciy6, Olciy6, Wlciy6;
wire Emciy6, Mmciy6, Umciy6, Cnciy6, Knciy6, Snciy6, Aociy6, Iociy6, Qociy6, Yociy6;
wire Gpciy6, Opciy6, Wpciy6, Eqciy6, Mqciy6, Uqciy6, Crciy6, Krciy6, Srciy6, Asciy6;
wire Isciy6, Qsciy6, Ysciy6, Gtciy6, Otciy6, Wtciy6, Euciy6, Muciy6, Uuciy6, Cvciy6;
wire Kvciy6, Svciy6, Awciy6, Iwciy6, Qwciy6, Ywciy6, Gxciy6, Oxciy6, Wxciy6, Eyciy6;
wire Myciy6, Uyciy6, Czciy6, Kzciy6, Szciy6, A0diy6, I0diy6, Q0diy6, Y0diy6, G1diy6;
wire O1diy6, W1diy6, E2diy6, M2diy6, U2diy6, C3diy6, K3diy6, S3diy6, A4diy6, I4diy6;
wire Q4diy6, Y4diy6, G5diy6, O5diy6, W5diy6, E6diy6, M6diy6, U6diy6, C7diy6, K7diy6;
wire S7diy6, A8diy6, I8diy6, Q8diy6, Y8diy6, G9diy6, O9diy6, W9diy6, Eadiy6, Madiy6;
wire Uadiy6, Cbdiy6, Kbdiy6, Sbdiy6, Acdiy6, Icdiy6, Qcdiy6, Ycdiy6, Gddiy6, Oddiy6;
wire Wddiy6, Eediy6, Mediy6, Uediy6, Cfdiy6, Kfdiy6, Sfdiy6, Agdiy6, Igdiy6, Qgdiy6;
wire Ygdiy6, Ghdiy6, Ohdiy6, Whdiy6, Eidiy6, Midiy6, Uidiy6, Cjdiy6, Kjdiy6, Sjdiy6;
wire Akdiy6, Ikdiy6, Qkdiy6, Ykdiy6, Gldiy6, Oldiy6, Wldiy6, Emdiy6, Mmdiy6, Umdiy6;
wire Cndiy6, Kndiy6, Sndiy6, Aodiy6, Iodiy6, Qodiy6, Yodiy6, Gpdiy6, Opdiy6, Wpdiy6;
wire Eqdiy6, Mqdiy6, Uqdiy6, Crdiy6, Krdiy6, Srdiy6, Asdiy6, Isdiy6, Qsdiy6, Ysdiy6;
wire Gtdiy6, Otdiy6, Wtdiy6, Eudiy6, Mudiy6, Uudiy6, Cvdiy6, Kvdiy6, Svdiy6, Awdiy6;
wire Iwdiy6, Qwdiy6, Ywdiy6, Gxdiy6, Oxdiy6, Wxdiy6, Eydiy6, Mydiy6, Uydiy6, Czdiy6;
wire Kzdiy6, Szdiy6, A0eiy6, I0eiy6, Q0eiy6, Y0eiy6, G1eiy6, O1eiy6, W1eiy6, E2eiy6;
wire M2eiy6, U2eiy6, C3eiy6, K3eiy6, S3eiy6, A4eiy6, I4eiy6, Q4eiy6, Y4eiy6, G5eiy6;
wire O5eiy6, W5eiy6, E6eiy6, M6eiy6, U6eiy6, C7eiy6, K7eiy6, S7eiy6, A8eiy6, I8eiy6;
wire Q8eiy6, Y8eiy6, G9eiy6, O9eiy6, W9eiy6, Eaeiy6, Maeiy6, Uaeiy6, Cbeiy6, Kbeiy6;
wire Sbeiy6, Aceiy6, Iceiy6, Qceiy6, Yceiy6, Gdeiy6, Odeiy6, Wdeiy6, Eeeiy6, Meeiy6;
wire Ueeiy6, Cfeiy6, Kfeiy6, Sfeiy6, Ageiy6, Igeiy6, Qgeiy6, Ygeiy6, Gheiy6, Oheiy6;
wire Wheiy6, Eieiy6, Mieiy6, Uieiy6, Cjeiy6, Kjeiy6, Sjeiy6, Akeiy6, Ikeiy6, Qkeiy6;
wire Ykeiy6, Gleiy6, Oleiy6, Wleiy6, Emeiy6, Mmeiy6, Umeiy6, Cneiy6, Kneiy6, Sneiy6;
wire Aoeiy6, Ioeiy6, Qoeiy6, Yoeiy6, Gpeiy6, Opeiy6, Wpeiy6, Eqeiy6, Mqeiy6, Uqeiy6;
wire Creiy6, Kreiy6, Sreiy6, Aseiy6, Iseiy6, Qseiy6, Yseiy6, Gteiy6, Oteiy6, Wteiy6;
wire Eueiy6, Mueiy6, Uueiy6, Cveiy6, Kveiy6, Sveiy6, Aweiy6, Iweiy6, Qweiy6, Yweiy6;
wire Gxeiy6, Oxeiy6, Wxeiy6, Eyeiy6, Myeiy6, Uyeiy6, Czeiy6, Kzeiy6, Szeiy6, A0fiy6;
wire I0fiy6, Q0fiy6, Y0fiy6, G1fiy6, O1fiy6, W1fiy6, E2fiy6, M2fiy6, U2fiy6, C3fiy6;
wire K3fiy6, S3fiy6, A4fiy6, I4fiy6, Q4fiy6, Y4fiy6, G5fiy6, O5fiy6, W5fiy6, E6fiy6;
wire M6fiy6, U6fiy6, C7fiy6, K7fiy6, S7fiy6, A8fiy6, I8fiy6, Q8fiy6, Y8fiy6, G9fiy6;
wire O9fiy6, W9fiy6, Eafiy6, Mafiy6, Uafiy6, Cbfiy6, Kbfiy6, Sbfiy6, Acfiy6, Icfiy6;
wire Qcfiy6, Ycfiy6, Gdfiy6, Odfiy6, Wdfiy6, Eefiy6, Mefiy6, Uefiy6, Cffiy6, Kffiy6;
wire Sffiy6, Agfiy6, Igfiy6, Qgfiy6, Ygfiy6, Ghfiy6, Ohfiy6, Whfiy6, Eifiy6, Mifiy6;
wire Uifiy6, Cjfiy6, Kjfiy6, Sjfiy6, Akfiy6, Ikfiy6, Qkfiy6, Ykfiy6, Glfiy6, Olfiy6;
wire Wlfiy6, Emfiy6, Mmfiy6, Umfiy6, Cnfiy6, Knfiy6, Snfiy6, Aofiy6, Iofiy6, Qofiy6;
wire Yofiy6, Gpfiy6, Opfiy6, Wpfiy6, Eqfiy6, Mqfiy6, Uqfiy6, Crfiy6, Krfiy6, Srfiy6;
wire Asfiy6, Isfiy6, Qsfiy6, Ysfiy6, Gtfiy6, Otfiy6, Wtfiy6, Eufiy6, Mufiy6, Uufiy6;
wire Cvfiy6, Kvfiy6, Svfiy6, Awfiy6, Iwfiy6, Qwfiy6, Ywfiy6, Gxfiy6, Oxfiy6, Wxfiy6;
wire Eyfiy6, Myfiy6, Uyfiy6, Czfiy6, Kzfiy6, Szfiy6, A0giy6, I0giy6, Q0giy6, Y0giy6;
wire G1giy6, O1giy6, W1giy6, E2giy6, M2giy6, U2giy6, C3giy6, K3giy6, S3giy6, A4giy6;
wire I4giy6, Q4giy6, Y4giy6, G5giy6, O5giy6, W5giy6, E6giy6, M6giy6, U6giy6, C7giy6;
wire K7giy6, S7giy6, A8giy6, I8giy6, Q8giy6, Y8giy6, G9giy6, O9giy6, W9giy6, Eagiy6;
wire Magiy6, Uagiy6, Cbgiy6, Kbgiy6, Sbgiy6, Acgiy6, Icgiy6, Qcgiy6, Ycgiy6, Gdgiy6;
wire Odgiy6, Wdgiy6, Eegiy6, Megiy6, Uegiy6, Cfgiy6, Kfgiy6, Sfgiy6, Aggiy6, Iggiy6;
wire Qggiy6, Yggiy6, Ghgiy6, Ohgiy6, Whgiy6, Eigiy6, Migiy6, Uigiy6, Cjgiy6, Kjgiy6;
wire Sjgiy6, Akgiy6, Ikgiy6, Qkgiy6, Ykgiy6, Glgiy6, Olgiy6, Wlgiy6, Emgiy6, Mmgiy6;
wire Umgiy6, Cngiy6, Kngiy6, Sngiy6, Aogiy6, Iogiy6, Qogiy6, Yogiy6, Gpgiy6, Opgiy6;
wire Wpgiy6, Eqgiy6, Mqgiy6, Uqgiy6, Crgiy6, Krgiy6, Srgiy6, Asgiy6, Isgiy6, Qsgiy6;
wire Ysgiy6, Gtgiy6, Otgiy6, Wtgiy6, Eugiy6, Mugiy6, Uugiy6, Cvgiy6, Kvgiy6, Svgiy6;
wire Awgiy6, Iwgiy6, Qwgiy6, Ywgiy6, Gxgiy6, Oxgiy6, Wxgiy6, Eygiy6, Mygiy6, Uygiy6;
wire Czgiy6, Kzgiy6, Szgiy6, A0hiy6, I0hiy6, Q0hiy6, Y0hiy6, G1hiy6, O1hiy6, W1hiy6;
wire E2hiy6, M2hiy6, U2hiy6, C3hiy6, K3hiy6, S3hiy6, A4hiy6, I4hiy6, Q4hiy6, Y4hiy6;
wire G5hiy6, O5hiy6, W5hiy6, E6hiy6, M6hiy6, U6hiy6, C7hiy6, K7hiy6, S7hiy6, A8hiy6;
wire I8hiy6, Q8hiy6, Y8hiy6, G9hiy6, O9hiy6, W9hiy6, Eahiy6, Mahiy6, Uahiy6, Cbhiy6;
wire Kbhiy6, Sbhiy6, Achiy6, Ichiy6, Qchiy6, Ychiy6, Gdhiy6, Odhiy6, Wdhiy6, Eehiy6;
wire Mehiy6, Uehiy6, Cfhiy6, Kfhiy6, Sfhiy6, Aghiy6, Ighiy6, Qghiy6, Yghiy6, Ghhiy6;
wire Ohhiy6, Whhiy6, Eihiy6, Mihiy6, Uihiy6, Cjhiy6, Kjhiy6, Sjhiy6, Akhiy6, Ikhiy6;
wire Qkhiy6, Ykhiy6, Glhiy6, Olhiy6, Wlhiy6, Emhiy6, Mmhiy6, Umhiy6, Cnhiy6, Knhiy6;
wire Snhiy6, Aohiy6, Iohiy6, Qohiy6, Yohiy6, Gphiy6, Ophiy6, Wphiy6, Eqhiy6, Mqhiy6;
wire Uqhiy6, Crhiy6, Krhiy6, Srhiy6, Ashiy6, Ishiy6, Qshiy6, Yshiy6, Gthiy6, Othiy6;
wire Wthiy6, Euhiy6, Muhiy6, Uuhiy6, Cvhiy6, Kvhiy6, Svhiy6, Awhiy6, Iwhiy6, Qwhiy6;
wire Ywhiy6, Gxhiy6, Oxhiy6, Wxhiy6, Eyhiy6, Myhiy6, Uyhiy6, Czhiy6, Kzhiy6, Szhiy6;
wire A0iiy6, I0iiy6, Q0iiy6, Y0iiy6, G1iiy6, O1iiy6, W1iiy6, E2iiy6, M2iiy6, U2iiy6;
wire C3iiy6, K3iiy6, S3iiy6, A4iiy6, I4iiy6, Q4iiy6, Y4iiy6, G5iiy6, O5iiy6, W5iiy6;
wire E6iiy6, M6iiy6, U6iiy6, C7iiy6, K7iiy6, S7iiy6, A8iiy6, I8iiy6, Q8iiy6, Y8iiy6;
wire G9iiy6, O9iiy6, W9iiy6, Eaiiy6, Maiiy6, Uaiiy6, Cbiiy6, Kbiiy6, Sbiiy6, Aciiy6;
wire Iciiy6, Qciiy6, Yciiy6, Gdiiy6, Odiiy6, Wdiiy6, Eeiiy6, Meiiy6, Ueiiy6, Cfiiy6;
wire Kfiiy6, Sfiiy6, Agiiy6, Igiiy6, Qgiiy6, Ygiiy6, Ghiiy6, Ohiiy6, Whiiy6, Eiiiy6;
wire Miiiy6, Uiiiy6, Cjiiy6, Kjiiy6, Sjiiy6, Akiiy6, Ikiiy6, Qkiiy6, Ykiiy6, Gliiy6;
wire Oliiy6, Wliiy6, Emiiy6, Mmiiy6, Umiiy6, Cniiy6, Kniiy6, Sniiy6, Aoiiy6, Ioiiy6;
wire Qoiiy6, Yoiiy6, Gpiiy6, Opiiy6, Wpiiy6, Eqiiy6, Mqiiy6, Uqiiy6, Criiy6, Kriiy6;
wire Sriiy6, Asiiy6, Isiiy6, Qsiiy6, Ysiiy6, Gtiiy6, Otiiy6, Wtiiy6, Euiiy6, Muiiy6;
wire Uuiiy6, Cviiy6, Kviiy6, Sviiy6, Awiiy6, Iwiiy6, Qwiiy6, Ywiiy6, Gxiiy6, Oxiiy6;
wire Wxiiy6, Eyiiy6, Myiiy6, Uyiiy6, Cziiy6, Kziiy6, Sziiy6, A0jiy6, I0jiy6, Q0jiy6;
wire Y0jiy6, G1jiy6, O1jiy6, W1jiy6, E2jiy6, M2jiy6, U2jiy6, C3jiy6, K3jiy6, S3jiy6;
wire A4jiy6, I4jiy6, Q4jiy6, Y4jiy6, G5jiy6, O5jiy6, W5jiy6, E6jiy6, M6jiy6, U6jiy6;
wire C7jiy6, K7jiy6, S7jiy6, A8jiy6, I8jiy6, Q8jiy6, Y8jiy6, G9jiy6, O9jiy6, W9jiy6;
wire Eajiy6, Majiy6, Uajiy6, Cbjiy6, Kbjiy6, Sbjiy6, Acjiy6, Icjiy6, Qcjiy6, Ycjiy6;
wire Gdjiy6, Odjiy6, Wdjiy6, Eejiy6, Mejiy6, Uejiy6, Cfjiy6, Kfjiy6, Sfjiy6, Agjiy6;
wire Igjiy6, Qgjiy6, Ygjiy6, Ghjiy6, Ohjiy6, Whjiy6, Eijiy6, Mijiy6, Uijiy6, Cjjiy6;
wire Kjjiy6, Sjjiy6, Akjiy6, Ikjiy6, Qkjiy6, Ykjiy6, Gljiy6, Oljiy6, Wljiy6, Emjiy6;
wire Mmjiy6, Umjiy6, Cnjiy6, Knjiy6, Snjiy6, Aojiy6, Iojiy6, Qojiy6, Yojiy6, Gpjiy6;
wire Opjiy6, Wpjiy6, Eqjiy6, Mqjiy6, Uqjiy6, Crjiy6, Krjiy6, Srjiy6, Asjiy6, Isjiy6;
wire Qsjiy6, Ysjiy6, Gtjiy6, Otjiy6, Wtjiy6, Eujiy6, Mujiy6, Uujiy6, Cvjiy6, Kvjiy6;
wire Svjiy6, Awjiy6, Iwjiy6, Qwjiy6, Ywjiy6, Gxjiy6, Oxjiy6, Wxjiy6, Eyjiy6, Myjiy6;
wire Uyjiy6, Czjiy6, Kzjiy6, Szjiy6, A0kiy6, I0kiy6, Q0kiy6, Y0kiy6, G1kiy6, O1kiy6;
wire W1kiy6, E2kiy6, M2kiy6, U2kiy6, C3kiy6, K3kiy6, S3kiy6, A4kiy6, I4kiy6, Q4kiy6;
wire Y4kiy6, G5kiy6, O5kiy6, W5kiy6, E6kiy6, M6kiy6, U6kiy6, C7kiy6, K7kiy6, S7kiy6;
wire A8kiy6, I8kiy6, Q8kiy6, Y8kiy6, G9kiy6, O9kiy6, W9kiy6, Eakiy6, Makiy6, Uakiy6;
wire Cbkiy6, Kbkiy6, Sbkiy6, Ackiy6, Ickiy6, Qckiy6, Yckiy6, Gdkiy6, Odkiy6, Wdkiy6;
wire Eekiy6, Mekiy6, Uekiy6, Cfkiy6, Kfkiy6, Sfkiy6, Agkiy6, Igkiy6, Qgkiy6, Ygkiy6;
wire Ghkiy6, Ohkiy6, Whkiy6, Eikiy6, Mikiy6, Uikiy6, Cjkiy6, Kjkiy6, Sjkiy6, Akkiy6;
wire Ikkiy6, Qkkiy6, Ykkiy6, Glkiy6, Olkiy6, Wlkiy6, Emkiy6, Mmkiy6, Umkiy6, Cnkiy6;
wire Knkiy6, Snkiy6, Aokiy6, Iokiy6, Qokiy6, Yokiy6, Gpkiy6, Opkiy6, Wpkiy6, Eqkiy6;
wire Mqkiy6, Uqkiy6, Crkiy6, Krkiy6, Srkiy6, Askiy6, Iskiy6, Qskiy6, Yskiy6, Gtkiy6;
wire Otkiy6, Wtkiy6, Eukiy6, Mukiy6, Uukiy6, Cvkiy6, Kvkiy6, Svkiy6, Awkiy6, Iwkiy6;
wire Qwkiy6, Ywkiy6, Gxkiy6, Oxkiy6, Wxkiy6, Eykiy6, Mykiy6, Uykiy6, Czkiy6, Kzkiy6;
wire Szkiy6, A0liy6, I0liy6, Q0liy6, Y0liy6, G1liy6, O1liy6, W1liy6, E2liy6, M2liy6;
wire U2liy6, C3liy6, K3liy6, S3liy6, A4liy6, I4liy6, Q4liy6, Y4liy6, G5liy6, O5liy6;
wire W5liy6, E6liy6, M6liy6, U6liy6, C7liy6, K7liy6, S7liy6, A8liy6, I8liy6, Q8liy6;
wire Y8liy6, G9liy6, O9liy6, W9liy6, Ealiy6, Maliy6, Ualiy6, Cbliy6, Kbliy6, Sbliy6;
wire Acliy6, Icliy6, Qcliy6, Ycliy6, Gdliy6, Odliy6, Wdliy6, Eeliy6, Meliy6, Ueliy6;
wire Cfliy6, Kfliy6, Sfliy6, Agliy6, Igliy6, Qgliy6, Ygliy6, Ghliy6, Ohliy6, Whliy6;
wire Eiliy6, Miliy6, Uiliy6, Cjliy6, Kjliy6, Sjliy6, Akliy6, Ikliy6, Qkliy6, Ykliy6;
wire Glliy6, Olliy6, Wlliy6, Emliy6, Mmliy6, Umliy6, Cnliy6, Knliy6, Snliy6, Aoliy6;
wire Ioliy6, Qoliy6, Yoliy6, Gpliy6, Opliy6, Wpliy6, Eqliy6, Mqliy6, Uqliy6, Crliy6;
wire Krliy6, Srliy6, Asliy6, Isliy6, Qsliy6, Ysliy6, Gtliy6, Otliy6, Wtliy6, Euliy6;
wire Muliy6, Uuliy6, Cvliy6, Kvliy6, Svliy6, Awliy6, Iwliy6, Qwliy6, Ywliy6, Gxliy6;
wire Oxliy6, Wxliy6, Eyliy6, Myliy6, Uyliy6, Czliy6, Kzliy6, Szliy6, A0miy6, I0miy6;
wire Q0miy6, Y0miy6, G1miy6, O1miy6, W1miy6, E2miy6, M2miy6, U2miy6, C3miy6, K3miy6;
wire S3miy6, A4miy6, I4miy6, Q4miy6, Y4miy6, G5miy6, O5miy6, W5miy6, E6miy6, M6miy6;
wire U6miy6, C7miy6, K7miy6, S7miy6, A8miy6, I8miy6, Q8miy6, Y8miy6, G9miy6, O9miy6;
wire W9miy6, Eamiy6, Mamiy6, Uamiy6, Cbmiy6, Kbmiy6, Sbmiy6, Acmiy6, Icmiy6, Qcmiy6;
wire Ycmiy6, Gdmiy6, Odmiy6, Wdmiy6, Eemiy6, Memiy6, Uemiy6, Cfmiy6, Kfmiy6, Sfmiy6;
wire Agmiy6, Igmiy6, Qgmiy6, Ygmiy6, Ghmiy6, Ohmiy6, Whmiy6, Eimiy6, Mimiy6, Uimiy6;
wire Cjmiy6, Kjmiy6, Sjmiy6, Akmiy6, Ikmiy6, Qkmiy6, Ykmiy6, Glmiy6, Olmiy6, Wlmiy6;
wire Emmiy6, Mmmiy6, Ummiy6, Cnmiy6, Knmiy6, Snmiy6, Aomiy6, Iomiy6, Qomiy6, Yomiy6;
wire Gpmiy6, Opmiy6, Wpmiy6, Eqmiy6, Mqmiy6, Uqmiy6, Crmiy6, Krmiy6, Srmiy6, Asmiy6;
wire Ismiy6, Qsmiy6, Ysmiy6, Gtmiy6, Otmiy6, Wtmiy6, Eumiy6, Mumiy6, Uumiy6, Cvmiy6;
wire Kvmiy6, Svmiy6, Awmiy6, Iwmiy6, Qwmiy6, Ywmiy6, Gxmiy6, Oxmiy6, Wxmiy6, Eymiy6;
wire Mymiy6, Uymiy6, Czmiy6, Kzmiy6, Szmiy6, A0niy6, I0niy6, Q0niy6, Y0niy6, G1niy6;
wire O1niy6, W1niy6, E2niy6, M2niy6, U2niy6, C3niy6, K3niy6, S3niy6, A4niy6, I4niy6;
wire Q4niy6, Y4niy6, G5niy6, O5niy6, W5niy6, E6niy6, M6niy6, U6niy6, C7niy6, K7niy6;
wire S7niy6, A8niy6, I8niy6, Q8niy6, Y8niy6, G9niy6, O9niy6, W9niy6, Eaniy6, Maniy6;
wire Uaniy6, Cbniy6, Kbniy6, Sbniy6, Acniy6, Icniy6, Qcniy6, Ycniy6, Gdniy6, Odniy6;
wire Wdniy6, Eeniy6, Meniy6, Ueniy6, Cfniy6, Kfniy6, Sfniy6, Agniy6, Igniy6, Qgniy6;
wire Ygniy6, Ghniy6, Ohniy6, Whniy6, Einiy6, Miniy6, Uiniy6, Cjniy6, Kjniy6, Sjniy6;
wire Akniy6, Ikniy6, Qkniy6, Ykniy6, Glniy6, Olniy6, Wlniy6, Emniy6, Mmniy6, Umniy6;
wire Cnniy6, Knniy6, Snniy6, Aoniy6, Ioniy6, Qoniy6, Yoniy6, Gpniy6, Opniy6, Wpniy6;
wire Eqniy6, Mqniy6, Uqniy6, Crniy6, Krniy6, Srniy6, Asniy6, Isniy6, Qsniy6, Ysniy6;
wire Gtniy6, Otniy6, Wtniy6, Euniy6, Muniy6, Uuniy6, Cvniy6, Kvniy6, Svniy6, Awniy6;
wire Iwniy6, Qwniy6, Ywniy6, Gxniy6, Oxniy6, Wxniy6, Eyniy6, Myniy6, Uyniy6, Czniy6;
wire Kzniy6, Szniy6, A0oiy6, I0oiy6, Q0oiy6, Y0oiy6, G1oiy6, O1oiy6, W1oiy6, E2oiy6;
wire M2oiy6, U2oiy6, C3oiy6, K3oiy6, S3oiy6, A4oiy6, I4oiy6, Q4oiy6, Y4oiy6, G5oiy6;
wire O5oiy6, W5oiy6, E6oiy6, M6oiy6, U6oiy6, C7oiy6, K7oiy6, S7oiy6, A8oiy6, I8oiy6;
wire Q8oiy6, Y8oiy6, G9oiy6, O9oiy6, W9oiy6, Eaoiy6, Maoiy6, Uaoiy6, Cboiy6, Kboiy6;
wire Sboiy6, Acoiy6, Icoiy6, Qcoiy6, Ycoiy6, Gdoiy6, Odoiy6, Wdoiy6, Eeoiy6, Meoiy6;
wire Ueoiy6, Cfoiy6, Kfoiy6, Sfoiy6, Agoiy6, Igoiy6, Qgoiy6, Ygoiy6, Ghoiy6, Ohoiy6;
wire Whoiy6, Eioiy6, Mioiy6, Uioiy6, Cjoiy6, Kjoiy6, Sjoiy6, Akoiy6, Ikoiy6, Qkoiy6;
wire Ykoiy6, Gloiy6, Oloiy6, Wloiy6, Emoiy6, Mmoiy6, Umoiy6, Cnoiy6, Knoiy6, Snoiy6;
wire Aooiy6, Iooiy6, Qooiy6, Yooiy6, Gpoiy6, Opoiy6, Wpoiy6, Eqoiy6, Mqoiy6, Uqoiy6;
wire Croiy6, Kroiy6, Sroiy6, Asoiy6, Isoiy6, Qsoiy6, Ysoiy6, Gtoiy6, Otoiy6, Wtoiy6;
wire Euoiy6, Muoiy6, Uuoiy6, Cvoiy6, Kvoiy6, Svoiy6, Awoiy6, Iwoiy6, Qwoiy6, Ywoiy6;
wire Gxoiy6, Oxoiy6, Wxoiy6, Eyoiy6, Myoiy6, Uyoiy6, Czoiy6, Kzoiy6, Szoiy6, A0piy6;
wire I0piy6, Q0piy6, Y0piy6, G1piy6, O1piy6, W1piy6, E2piy6, M2piy6, U2piy6, C3piy6;
wire K3piy6, S3piy6, A4piy6, I4piy6, Q4piy6, Y4piy6, G5piy6, O5piy6, W5piy6, E6piy6;
wire M6piy6, U6piy6, C7piy6, K7piy6, S7piy6, A8piy6, I8piy6, Q8piy6, Y8piy6, G9piy6;
wire O9piy6, W9piy6, Eapiy6, Mapiy6, Uapiy6, Cbpiy6, Kbpiy6, Sbpiy6, Acpiy6, Icpiy6;
wire Qcpiy6, Ycpiy6, Gdpiy6, Odpiy6, Wdpiy6, Eepiy6, Mepiy6, Uepiy6, Cfpiy6, Kfpiy6;
wire Sfpiy6, Agpiy6, Igpiy6, Qgpiy6, Ygpiy6, Ghpiy6, Ohpiy6, Whpiy6, Eipiy6, Mipiy6;
wire Uipiy6, Cjpiy6, Kjpiy6, Sjpiy6, Akpiy6, Ikpiy6, Qkpiy6, Ykpiy6, Glpiy6, Olpiy6;
wire Wlpiy6, Empiy6, Mmpiy6, Umpiy6, Cnpiy6, Knpiy6, Snpiy6, Aopiy6, Iopiy6, Qopiy6;
wire Yopiy6, Gppiy6, Oppiy6, Wppiy6, Eqpiy6, Mqpiy6, Uqpiy6, Crpiy6, Krpiy6, Srpiy6;
wire Aspiy6, Ispiy6, Qspiy6, Yspiy6, Gtpiy6, Otpiy6, Wtpiy6, Eupiy6, Mupiy6, Uupiy6;
wire Cvpiy6, Kvpiy6, Svpiy6, Awpiy6, Iwpiy6, Qwpiy6, Ywpiy6, Gxpiy6, Oxpiy6, Wxpiy6;
wire Eypiy6, Mypiy6, Uypiy6, Czpiy6, Kzpiy6, Szpiy6, A0qiy6, I0qiy6, Q0qiy6, Y0qiy6;
wire G1qiy6, O1qiy6, W1qiy6, E2qiy6, M2qiy6, U2qiy6, C3qiy6, K3qiy6, S3qiy6, A4qiy6;
wire I4qiy6, Q4qiy6, Y4qiy6, G5qiy6, O5qiy6, W5qiy6, E6qiy6, M6qiy6, U6qiy6, C7qiy6;
wire K7qiy6, S7qiy6, A8qiy6, I8qiy6, Q8qiy6, Y8qiy6, G9qiy6, O9qiy6, W9qiy6, Eaqiy6;
wire Maqiy6, Uaqiy6, Cbqiy6, Kbqiy6, Sbqiy6, Acqiy6, Icqiy6, Qcqiy6, Ycqiy6, Gdqiy6;
wire Odqiy6, Wdqiy6, Eeqiy6, Meqiy6, Ueqiy6, Cfqiy6, Kfqiy6, Sfqiy6, Agqiy6, Igqiy6;
wire Qgqiy6, Ygqiy6, Ghqiy6, Ohqiy6, Whqiy6, Eiqiy6, Miqiy6, Uiqiy6, Cjqiy6, Kjqiy6;
wire Sjqiy6, Akqiy6, Ikqiy6, Qkqiy6, Ykqiy6, Glqiy6, Olqiy6, Wlqiy6, Emqiy6, Mmqiy6;
wire Umqiy6, Cnqiy6, Knqiy6, Snqiy6, Aoqiy6, Ioqiy6, Qoqiy6, Yoqiy6, Gpqiy6, Opqiy6;
wire Wpqiy6, Eqqiy6, Mqqiy6, Uqqiy6, Crqiy6, Krqiy6, Srqiy6, Asqiy6, Isqiy6, Qsqiy6;
wire Ysqiy6, Gtqiy6, Otqiy6, Wtqiy6, Euqiy6, Muqiy6, Uuqiy6, Cvqiy6, Kvqiy6, Svqiy6;
wire Awqiy6, Iwqiy6, Qwqiy6, Ywqiy6, Gxqiy6, Oxqiy6, Wxqiy6, Eyqiy6, Myqiy6, Uyqiy6;
wire Czqiy6, Kzqiy6, Szqiy6, A0riy6, I0riy6, Q0riy6, Y0riy6, G1riy6, O1riy6, W1riy6;
wire E2riy6, M2riy6, U2riy6, C3riy6, K3riy6, S3riy6, A4riy6, I4riy6, Q4riy6, Y4riy6;
wire G5riy6, O5riy6, W5riy6, E6riy6, M6riy6, U6riy6, C7riy6, K7riy6, S7riy6, A8riy6;
wire I8riy6, Q8riy6, Y8riy6, G9riy6, O9riy6, W9riy6, Eariy6, Mariy6, Uariy6, Cbriy6;
wire Kbriy6, Sbriy6, Acriy6, Icriy6, Qcriy6, Ycriy6, Gdriy6, Odriy6, Wdriy6, Eeriy6;
wire Meriy6, Ueriy6, Cfriy6, Kfriy6, Sfriy6, Agriy6, Igriy6, Qgriy6, Ygriy6, Ghriy6;
wire Ohriy6, Whriy6, Eiriy6, Miriy6, Uiriy6, Cjriy6, Kjriy6, Sjriy6, Akriy6, Ikriy6;
wire Qkriy6, Ykriy6, Glriy6, Olriy6, Wlriy6, Emriy6, Mmriy6, Umriy6, Cnriy6, Knriy6;
wire Snriy6, Aoriy6, Ioriy6, Qoriy6, Yoriy6, Gpriy6, Opriy6, Wpriy6, Eqriy6, Mqriy6;
wire Uqriy6, Crriy6, Krriy6, Srriy6, Asriy6, Isriy6, Qsriy6, Ysriy6, Gtriy6, Otriy6;
wire Wtriy6, Euriy6, Muriy6, Uuriy6, Cvriy6, Kvriy6, Svriy6, Awriy6, Iwriy6, Qwriy6;
wire Ywriy6, Gxriy6, Oxriy6, Wxriy6, Eyriy6, Myriy6, Uyriy6, Czriy6, Kzriy6, Szriy6;
wire A0siy6, I0siy6, Q0siy6, Y0siy6, G1siy6, O1siy6, W1siy6, E2siy6, M2siy6, U2siy6;
wire C3siy6, K3siy6, S3siy6, A4siy6, I4siy6, Q4siy6, Y4siy6, G5siy6, O5siy6, W5siy6;
wire E6siy6, M6siy6, U6siy6, C7siy6, K7siy6, S7siy6, A8siy6, I8siy6, Q8siy6, Y8siy6;
wire G9siy6, O9siy6, W9siy6, Easiy6, Masiy6, Uasiy6, Cbsiy6, Kbsiy6, Sbsiy6, Acsiy6;
wire Icsiy6, Qcsiy6, Ycsiy6, Gdsiy6, Odsiy6, Wdsiy6, Eesiy6, Mesiy6, Uesiy6, Cfsiy6;
wire Kfsiy6, Sfsiy6, Agsiy6, Igsiy6, Qgsiy6, Ygsiy6, Ghsiy6, Ohsiy6, Whsiy6, Eisiy6;
wire Misiy6, Uisiy6, Cjsiy6, Kjsiy6, Sjsiy6, Aksiy6, Iksiy6, Qksiy6, Yksiy6, Glsiy6;
wire Olsiy6, Wlsiy6, Emsiy6, Mmsiy6, Umsiy6, Cnsiy6, Knsiy6, Snsiy6, Aosiy6, Iosiy6;
wire Qosiy6, Yosiy6, Gpsiy6, Opsiy6, Wpsiy6, Eqsiy6, Mqsiy6, Uqsiy6, Crsiy6, Krsiy6;
wire Srsiy6, Assiy6, Issiy6, Qssiy6, Yssiy6, Gtsiy6, Otsiy6, Wtsiy6, Eusiy6, Musiy6;
wire Uusiy6, Cvsiy6, Kvsiy6, Svsiy6, Awsiy6, Iwsiy6, Qwsiy6, Ywsiy6, Gxsiy6, Oxsiy6;
wire Wxsiy6, Eysiy6, Mysiy6, Uysiy6, Czsiy6, Kzsiy6, Szsiy6, A0tiy6, I0tiy6, Q0tiy6;
wire Y0tiy6, G1tiy6, O1tiy6, W1tiy6, E2tiy6, M2tiy6, U2tiy6, C3tiy6, K3tiy6, S3tiy6;
wire A4tiy6, I4tiy6, Q4tiy6, Y4tiy6, G5tiy6, O5tiy6, W5tiy6, E6tiy6, M6tiy6, U6tiy6;
wire C7tiy6, K7tiy6, S7tiy6, A8tiy6, I8tiy6, Q8tiy6, Y8tiy6, G9tiy6, O9tiy6, W9tiy6;
wire Eatiy6, Matiy6, Uatiy6, Cbtiy6, Kbtiy6, Sbtiy6, Actiy6, Ictiy6, Qctiy6, Yctiy6;
wire Gdtiy6, Odtiy6, Wdtiy6, Eetiy6, Metiy6, Uetiy6, Cftiy6, Kftiy6, Sftiy6, Agtiy6;
wire Igtiy6, Qgtiy6, Ygtiy6, Ghtiy6, Ohtiy6, Whtiy6, Eitiy6, Mitiy6, Uitiy6, Cjtiy6;
wire Kjtiy6, Sjtiy6, Aktiy6, Iktiy6, Qktiy6, Yktiy6, Gltiy6, Oltiy6, Wltiy6, Emtiy6;
wire Mmtiy6, Umtiy6, Cntiy6, Kntiy6, Sntiy6, Aotiy6, Iotiy6, Qotiy6, Yotiy6, Gptiy6;
wire Optiy6, Wptiy6, Eqtiy6, Mqtiy6, Uqtiy6, Crtiy6, Krtiy6, Srtiy6, Astiy6, Istiy6;
wire Qstiy6, Ystiy6, Gttiy6, Ottiy6, Wttiy6, Eutiy6, Mutiy6, Uutiy6, Cvtiy6, Kvtiy6;
wire Svtiy6, Awtiy6, Iwtiy6, Qwtiy6, Ywtiy6, Gxtiy6, Oxtiy6, Wxtiy6, Eytiy6, Mytiy6;
wire Uytiy6, Cztiy6, Kztiy6, Sztiy6, A0uiy6, I0uiy6, Q0uiy6, Y0uiy6, G1uiy6, O1uiy6;
wire W1uiy6, E2uiy6, M2uiy6, U2uiy6, C3uiy6, K3uiy6, S3uiy6, A4uiy6, I4uiy6, Q4uiy6;
wire Y4uiy6, G5uiy6, O5uiy6, W5uiy6, E6uiy6, M6uiy6, U6uiy6, C7uiy6, K7uiy6, S7uiy6;
wire A8uiy6, I8uiy6, Q8uiy6, Y8uiy6, G9uiy6, O9uiy6, W9uiy6, Eauiy6, Mauiy6, Uauiy6;
wire Cbuiy6, Kbuiy6, Sbuiy6, Acuiy6, Icuiy6, Qcuiy6, Ycuiy6, Gduiy6, Oduiy6, Wduiy6;
wire Eeuiy6, Meuiy6, Ueuiy6, Cfuiy6, Kfuiy6, Sfuiy6, Aguiy6, Iguiy6, Qguiy6, Yguiy6;
wire Ghuiy6, Ohuiy6, Whuiy6, Eiuiy6, Miuiy6, Uiuiy6, Cjuiy6, Kjuiy6, Sjuiy6, Akuiy6;
wire Ikuiy6, Qkuiy6, Ykuiy6, Gluiy6, Oluiy6, Wluiy6, Emuiy6, Mmuiy6, Umuiy6, Cnuiy6;
wire Knuiy6, Snuiy6, Aouiy6, Iouiy6, Qouiy6, Youiy6, Gpuiy6, Opuiy6, Wpuiy6, Equiy6;
wire Mquiy6, Uquiy6, Cruiy6, Kruiy6, Sruiy6, Asuiy6, Isuiy6, Qsuiy6, Ysuiy6, Gtuiy6;
wire Otuiy6, Wtuiy6, Euuiy6, Muuiy6, Uuuiy6, Cvuiy6, Kvuiy6, Svuiy6, Awuiy6, Iwuiy6;
wire Qwuiy6, Ywuiy6, Gxuiy6, Oxuiy6, Wxuiy6, Eyuiy6, Myuiy6, Uyuiy6, Czuiy6, Kzuiy6;
wire Szuiy6, A0viy6, I0viy6, Q0viy6, Y0viy6, G1viy6, O1viy6, W1viy6, E2viy6, M2viy6;
wire U2viy6, C3viy6, K3viy6, S3viy6, A4viy6, I4viy6, Q4viy6, Y4viy6, G5viy6, O5viy6;
wire W5viy6, E6viy6, M6viy6, U6viy6, C7viy6, K7viy6, S7viy6, A8viy6, I8viy6, Q8viy6;
wire Y8viy6, G9viy6, O9viy6, W9viy6, Eaviy6, Maviy6, Uaviy6, Cbviy6, Kbviy6, Sbviy6;
wire Acviy6, Icviy6, Qcviy6, Ycviy6, Gdviy6, Odviy6, Wdviy6, Eeviy6, Meviy6, Ueviy6;
wire Cfviy6, Kfviy6, Sfviy6, Agviy6, Igviy6, Qgviy6, Ygviy6, Ghviy6, Ohviy6, Whviy6;
wire Eiviy6, Miviy6, Uiviy6, Cjviy6, Kjviy6, Sjviy6, Akviy6, Ikviy6, Qkviy6, Ykviy6;
wire Glviy6, Olviy6, Wlviy6, Emviy6, Mmviy6, Umviy6, Cnviy6, Knviy6, Snviy6, Aoviy6;
wire Ioviy6, Qoviy6, Yoviy6, Gpviy6, Opviy6, Wpviy6, Eqviy6, Mqviy6, Uqviy6, Crviy6;
wire Krviy6, Srviy6, Asviy6, Isviy6, Qsviy6, Ysviy6, Gtviy6, Otviy6, Wtviy6, Euviy6;
wire Muviy6, Uuviy6, Cvviy6, Kvviy6, Svviy6, Awviy6, Iwviy6, Qwviy6, Ywviy6, Gxviy6;
wire Oxviy6, Wxviy6, Eyviy6, Myviy6, Uyviy6, Czviy6, Kzviy6, Szviy6, A0wiy6, I0wiy6;
wire Q0wiy6, Y0wiy6, G1wiy6, O1wiy6, W1wiy6, E2wiy6, M2wiy6, U2wiy6, C3wiy6, K3wiy6;
wire S3wiy6, A4wiy6, I4wiy6, Q4wiy6, Y4wiy6, G5wiy6, O5wiy6, W5wiy6, E6wiy6, M6wiy6;
wire U6wiy6, C7wiy6, K7wiy6, S7wiy6, A8wiy6, I8wiy6, Q8wiy6, Y8wiy6, G9wiy6, O9wiy6;
wire W9wiy6, Eawiy6, Mawiy6, Uawiy6, Cbwiy6, Kbwiy6, Sbwiy6, Acwiy6, Icwiy6, Qcwiy6;
wire Ycwiy6, Gdwiy6, Odwiy6, Wdwiy6, Eewiy6, Mewiy6, Uewiy6, Cfwiy6, Kfwiy6, Sfwiy6;
wire Agwiy6, Igwiy6, Qgwiy6, Ygwiy6, Ghwiy6, Ohwiy6, Whwiy6, Eiwiy6, Miwiy6, Uiwiy6;
wire Cjwiy6, Kjwiy6, Sjwiy6, Akwiy6, Ikwiy6, Qkwiy6, Ykwiy6, Glwiy6, Olwiy6, Wlwiy6;
wire Emwiy6, Mmwiy6, Umwiy6, Cnwiy6, Knwiy6, Snwiy6, Aowiy6, Iowiy6, Qowiy6, Yowiy6;
wire Gpwiy6, Opwiy6, Wpwiy6, Eqwiy6, Mqwiy6, Uqwiy6, Crwiy6, Krwiy6, Srwiy6, Aswiy6;
wire Iswiy6, Qswiy6, Yswiy6, Gtwiy6, Otwiy6, Wtwiy6, Euwiy6, Muwiy6, Uuwiy6, Cvwiy6;
wire Kvwiy6, Svwiy6, Awwiy6, Iwwiy6, Qwwiy6, Ywwiy6, Gxwiy6, Oxwiy6, Wxwiy6, Eywiy6;
wire Mywiy6, Uywiy6, Czwiy6, Kzwiy6, Szwiy6, A0xiy6, I0xiy6, Q0xiy6, Y0xiy6, G1xiy6;
wire O1xiy6, W1xiy6, E2xiy6, M2xiy6, U2xiy6, C3xiy6, K3xiy6, S3xiy6, A4xiy6, I4xiy6;
wire Q4xiy6, Y4xiy6, G5xiy6, O5xiy6, W5xiy6, E6xiy6, M6xiy6, U6xiy6, C7xiy6, K7xiy6;
wire S7xiy6, A8xiy6, I8xiy6, Q8xiy6, Y8xiy6, G9xiy6, O9xiy6, W9xiy6, Eaxiy6, Maxiy6;
wire Uaxiy6, Cbxiy6, Kbxiy6, Sbxiy6, Acxiy6, Icxiy6, Qcxiy6, Ycxiy6, Gdxiy6, Odxiy6;
wire Wdxiy6, Eexiy6, Mexiy6, Uexiy6, Cfxiy6, Kfxiy6, Sfxiy6, Agxiy6, Igxiy6, Qgxiy6;
wire Ygxiy6, Ghxiy6, Ohxiy6, Whxiy6, Eixiy6, Mixiy6, Uixiy6, Cjxiy6, Kjxiy6, Sjxiy6;
wire Akxiy6, Ikxiy6, Qkxiy6, Ykxiy6, Glxiy6, Olxiy6, Wlxiy6, Emxiy6, Mmxiy6, Umxiy6;
wire Cnxiy6, Knxiy6, Snxiy6, Aoxiy6, Ioxiy6, Qoxiy6, Yoxiy6, Gpxiy6, Opxiy6, Wpxiy6;
wire Eqxiy6, Mqxiy6, Uqxiy6, Crxiy6, Krxiy6, Srxiy6, Asxiy6, Isxiy6, Qsxiy6, Ysxiy6;
wire Gtxiy6, Otxiy6, Wtxiy6, Euxiy6, Muxiy6, Uuxiy6, Cvxiy6, Kvxiy6, Svxiy6, Awxiy6;
wire Iwxiy6, Qwxiy6, Ywxiy6, Gxxiy6, Oxxiy6, Wxxiy6, Eyxiy6, Myxiy6, Uyxiy6, Czxiy6;
wire Kzxiy6, Szxiy6, A0yiy6, I0yiy6, Q0yiy6, Y0yiy6, G1yiy6, O1yiy6, W1yiy6, E2yiy6;
wire M2yiy6, U2yiy6, C3yiy6, K3yiy6, S3yiy6, A4yiy6, I4yiy6, Q4yiy6, Y4yiy6, G5yiy6;
wire O5yiy6, W5yiy6, E6yiy6, M6yiy6, U6yiy6, C7yiy6, K7yiy6, S7yiy6, A8yiy6, I8yiy6;
wire Q8yiy6, Y8yiy6, G9yiy6, O9yiy6, W9yiy6, Eayiy6, Mayiy6, Uayiy6, Cbyiy6, Kbyiy6;
wire Sbyiy6, Acyiy6, Icyiy6, Qcyiy6, Ycyiy6, Gdyiy6, Odyiy6, Wdyiy6, Eeyiy6, Meyiy6;
wire Ueyiy6, Cfyiy6, Kfyiy6, Sfyiy6, Agyiy6, Igyiy6, Qgyiy6, Ygyiy6, Ghyiy6, Ohyiy6;
wire Whyiy6, Eiyiy6, Miyiy6, Uiyiy6, Cjyiy6, Kjyiy6, Sjyiy6, Akyiy6, Ikyiy6, Qkyiy6;
wire Ykyiy6, Glyiy6, Olyiy6, Wlyiy6, Emyiy6, Mmyiy6, Umyiy6, Cnyiy6, Knyiy6, Snyiy6;
wire Aoyiy6, Ioyiy6, Qoyiy6, Yoyiy6, Gpyiy6, Opyiy6, Wpyiy6, Eqyiy6, Mqyiy6, Uqyiy6;
wire Cryiy6, Kryiy6, Sryiy6, Asyiy6, Isyiy6, Qsyiy6, Ysyiy6, Gtyiy6, Otyiy6, Wtyiy6;
wire Euyiy6, Muyiy6, Uuyiy6, Cvyiy6, Kvyiy6, Svyiy6, Awyiy6, Iwyiy6, Qwyiy6, Ywyiy6;
wire Gxyiy6, Oxyiy6, Wxyiy6, Eyyiy6, Myyiy6, Uyyiy6, Czyiy6, Kzyiy6, Szyiy6, A0ziy6;
wire I0ziy6, Q0ziy6, Y0ziy6, G1ziy6, O1ziy6, W1ziy6, E2ziy6, M2ziy6, U2ziy6, C3ziy6;
wire K3ziy6, S3ziy6, A4ziy6, I4ziy6, Q4ziy6, Y4ziy6, G5ziy6, O5ziy6, W5ziy6, E6ziy6;
wire M6ziy6, U6ziy6, C7ziy6, K7ziy6, S7ziy6, A8ziy6, I8ziy6, Q8ziy6, Y8ziy6, G9ziy6;
wire O9ziy6, W9ziy6, Eaziy6, Maziy6, Uaziy6, Cbziy6, Kbziy6, Sbziy6, Acziy6, Icziy6;
wire Qcziy6, Ycziy6, Gdziy6, Odziy6, Wdziy6, Eeziy6, Meziy6, Ueziy6, Cfziy6, Kfziy6;
wire Sfziy6, Agziy6, Igziy6, Qgziy6, Ygziy6, Ghziy6, Ohziy6, Whziy6, Eiziy6, Miziy6;
wire Uiziy6, Cjziy6, Kjziy6, Sjziy6, Akziy6, Ikziy6, Qkziy6, Ykziy6, Glziy6, Olziy6;
wire Wlziy6, Emziy6, Mmziy6, Umziy6, Cnziy6, Knziy6, Snziy6, Aoziy6, Ioziy6, Qoziy6;
wire Yoziy6, Gpziy6, Opziy6, Wpziy6, Eqziy6, Mqziy6, Uqziy6, Crziy6, Krziy6, Srziy6;
wire Asziy6, Isziy6, Qsziy6, Ysziy6, Gtziy6, Otziy6, Wtziy6, Euziy6, Muziy6, Uuziy6;
wire Cvziy6, Kvziy6, Svziy6, Awziy6, Iwziy6, Qwziy6, Ywziy6, Gxziy6, Oxziy6, Wxziy6;
wire Eyziy6, Myziy6, Uyziy6, Czziy6, Kzziy6, Szziy6, A00jy6, I00jy6, Q00jy6, Y00jy6;
wire G10jy6, O10jy6, W10jy6, E20jy6, M20jy6, U20jy6, C30jy6, K30jy6, S30jy6, A40jy6;
wire I40jy6, Q40jy6, Y40jy6, G50jy6, O50jy6, W50jy6, E60jy6, M60jy6, U60jy6, C70jy6;
wire K70jy6, S70jy6, A80jy6, I80jy6, Q80jy6, Y80jy6, G90jy6, O90jy6, W90jy6, Ea0jy6;
wire Ma0jy6, Ua0jy6, Cb0jy6, Kb0jy6, Sb0jy6, Ac0jy6, Ic0jy6, Qc0jy6, Yc0jy6, Gd0jy6;
wire Od0jy6, Wd0jy6, Ee0jy6, Me0jy6, Ue0jy6, Cf0jy6, Kf0jy6, Sf0jy6, Ag0jy6, Ig0jy6;
wire Qg0jy6, Yg0jy6, Gh0jy6, Oh0jy6, Wh0jy6, Ei0jy6, Mi0jy6, Ui0jy6, Cj0jy6, Kj0jy6;
wire Sj0jy6, Ak0jy6, Ik0jy6, Qk0jy6, Yk0jy6, Gl0jy6, Ol0jy6, Wl0jy6, Em0jy6, Mm0jy6;
wire Um0jy6, Cn0jy6, Kn0jy6, Sn0jy6, Ao0jy6, Io0jy6, Qo0jy6, Yo0jy6, Gp0jy6, Op0jy6;
wire Wp0jy6, Eq0jy6, Mq0jy6, Uq0jy6, Cr0jy6, Kr0jy6, Sr0jy6, As0jy6, Is0jy6, Qs0jy6;
wire Ys0jy6, Gt0jy6, Ot0jy6, Wt0jy6, Eu0jy6, Mu0jy6, Uu0jy6, Cv0jy6, Kv0jy6, Sv0jy6;
wire Aw0jy6, Iw0jy6, Qw0jy6, Yw0jy6, Gx0jy6, Ox0jy6, Wx0jy6, Ey0jy6, My0jy6, Uy0jy6;
wire Cz0jy6, Kz0jy6, Sz0jy6, A01jy6, I01jy6, Q01jy6, Y01jy6, G11jy6, O11jy6, W11jy6;
wire E21jy6, M21jy6, U21jy6, C31jy6, K31jy6, S31jy6, A41jy6, I41jy6, Q41jy6, Y41jy6;
wire G51jy6, O51jy6, W51jy6, E61jy6, M61jy6, U61jy6, C71jy6, K71jy6, S71jy6, A81jy6;
wire I81jy6, Q81jy6, Y81jy6, G91jy6, O91jy6, W91jy6, Ea1jy6, Ma1jy6, Ua1jy6, Cb1jy6;
wire Kb1jy6, Sb1jy6, Ac1jy6, Ic1jy6, Qc1jy6, Yc1jy6, Gd1jy6, Od1jy6, Wd1jy6, Ee1jy6;
wire Me1jy6, Ue1jy6, Cf1jy6, Kf1jy6, Sf1jy6, Ag1jy6, Ig1jy6, Qg1jy6, Yg1jy6, Gh1jy6;
wire Oh1jy6, Wh1jy6, Ei1jy6, Mi1jy6, Ui1jy6, Cj1jy6, Kj1jy6, Sj1jy6, Ak1jy6, Ik1jy6;
wire Qk1jy6, Yk1jy6, Gl1jy6, Ol1jy6, Wl1jy6, Em1jy6, Mm1jy6, Um1jy6, Cn1jy6, Kn1jy6;
wire Sn1jy6, Ao1jy6, Io1jy6, Qo1jy6, Yo1jy6, Gp1jy6, Op1jy6, Wp1jy6, Eq1jy6, Mq1jy6;
wire Uq1jy6, Cr1jy6, Kr1jy6, Sr1jy6, As1jy6, Is1jy6, Qs1jy6, Ys1jy6, Gt1jy6, Ot1jy6;
wire Wt1jy6, Eu1jy6, Mu1jy6, Uu1jy6, Cv1jy6, Kv1jy6, Sv1jy6, Aw1jy6, Iw1jy6, Qw1jy6;
wire Yw1jy6, Gx1jy6, Ox1jy6, Wx1jy6, Ey1jy6, My1jy6, Uy1jy6, Cz1jy6, Kz1jy6, Sz1jy6;
wire A02jy6, I02jy6, Q02jy6, Y02jy6, G12jy6, O12jy6, W12jy6, E22jy6, M22jy6, U22jy6;
wire C32jy6, K32jy6, S32jy6, A42jy6, I42jy6, Q42jy6, Y42jy6, G52jy6, O52jy6, W52jy6;
wire E62jy6, M62jy6, U62jy6, C72jy6, K72jy6, S72jy6, A82jy6, I82jy6, Q82jy6, Y82jy6;
wire G92jy6, O92jy6, W92jy6, Ea2jy6, Ma2jy6, Ua2jy6, Cb2jy6, Kb2jy6, Sb2jy6, Ac2jy6;
wire Ic2jy6, Qc2jy6, Yc2jy6, Gd2jy6, Od2jy6, Wd2jy6, Ee2jy6, Me2jy6, Ue2jy6, Cf2jy6;
wire Kf2jy6, Sf2jy6, Ag2jy6, Ig2jy6, Qg2jy6, Yg2jy6, Gh2jy6, Oh2jy6, Wh2jy6, Ei2jy6;
wire Mi2jy6, Ui2jy6, Cj2jy6, Kj2jy6, Sj2jy6, Ak2jy6, Ik2jy6, Qk2jy6, Yk2jy6, Gl2jy6;
wire Ol2jy6, Wl2jy6, Em2jy6, Mm2jy6, Um2jy6, Cn2jy6, Kn2jy6, Sn2jy6, Ao2jy6, Io2jy6;
wire Qo2jy6, Yo2jy6, Gp2jy6, Op2jy6, Wp2jy6, Eq2jy6, Mq2jy6, Uq2jy6, Cr2jy6, Kr2jy6;
wire Sr2jy6, As2jy6, Is2jy6, Qs2jy6, Ys2jy6, Gt2jy6, Ot2jy6, Wt2jy6, Eu2jy6, Mu2jy6;
wire Uu2jy6, Cv2jy6, Kv2jy6, Sv2jy6, Aw2jy6, Iw2jy6, Qw2jy6, Yw2jy6, Gx2jy6, Ox2jy6;
wire Wx2jy6, Ey2jy6, My2jy6, Uy2jy6, Cz2jy6, Kz2jy6, Sz2jy6, A03jy6, I03jy6, Q03jy6;
wire Y03jy6, G13jy6, O13jy6, W13jy6, E23jy6, M23jy6, U23jy6, C33jy6, K33jy6, S33jy6;
wire A43jy6, I43jy6, Q43jy6, Y43jy6, G53jy6, O53jy6, W53jy6, E63jy6, M63jy6, U63jy6;
wire C73jy6, K73jy6, S73jy6, A83jy6, I83jy6, Q83jy6, Y83jy6, G93jy6, O93jy6, W93jy6;
wire Ea3jy6, Ma3jy6, Ua3jy6, Cb3jy6, Kb3jy6, Sb3jy6, Ac3jy6, Ic3jy6, Qc3jy6, Yc3jy6;
wire Gd3jy6, Od3jy6, Wd3jy6, Ee3jy6, Me3jy6, Ue3jy6, Cf3jy6, Kf3jy6, Sf3jy6, Ag3jy6;
wire Ig3jy6, Qg3jy6, Yg3jy6, Gh3jy6, Oh3jy6, Wh3jy6, Ei3jy6, Mi3jy6, Ui3jy6, Cj3jy6;
wire Kj3jy6, Sj3jy6, Ak3jy6, Ik3jy6, Qk3jy6, Yk3jy6, Gl3jy6, Ol3jy6, Wl3jy6, Em3jy6;
wire Mm3jy6, Um3jy6, Cn3jy6, Kn3jy6, Sn3jy6, Ao3jy6, Io3jy6, Qo3jy6, Yo3jy6, Gp3jy6;
wire Op3jy6, Wp3jy6, Eq3jy6, Mq3jy6, Uq3jy6, Cr3jy6, Kr3jy6, Sr3jy6, As3jy6, Is3jy6;
wire Qs3jy6, Ys3jy6, Gt3jy6, Ot3jy6, Wt3jy6, Eu3jy6, Mu3jy6, Uu3jy6, Cv3jy6, Kv3jy6;
wire Sv3jy6, Aw3jy6, Iw3jy6, Qw3jy6, Yw3jy6, Gx3jy6, Ox3jy6, Wx3jy6, Ey3jy6, My3jy6;
wire Uy3jy6, Cz3jy6, Kz3jy6, Sz3jy6, A04jy6, I04jy6, Q04jy6, Y04jy6, G14jy6, O14jy6;
wire W14jy6, E24jy6, M24jy6, U24jy6, C34jy6, K34jy6, S34jy6, A44jy6, I44jy6, Q44jy6;
wire Y44jy6, G54jy6, O54jy6, W54jy6, E64jy6, M64jy6, U64jy6, C74jy6, K74jy6, S74jy6;
wire A84jy6, I84jy6, Q84jy6, Y84jy6, G94jy6, O94jy6, W94jy6, Ea4jy6, Ma4jy6, Ua4jy6;
wire Cb4jy6, Kb4jy6, Sb4jy6, Ac4jy6, Ic4jy6, Qc4jy6, Yc4jy6, Gd4jy6, Od4jy6, Wd4jy6;
wire Ee4jy6, Me4jy6, Ue4jy6, Cf4jy6, Kf4jy6, Sf4jy6, Ag4jy6, Ig4jy6, Qg4jy6, Yg4jy6;
wire Gh4jy6, Oh4jy6, Wh4jy6, Ei4jy6, Mi4jy6, Ui4jy6, Cj4jy6, Kj4jy6, Sj4jy6, Ak4jy6;
wire Ik4jy6, Qk4jy6, Yk4jy6, Gl4jy6, Ol4jy6, Wl4jy6, Em4jy6, Mm4jy6, Um4jy6, Cn4jy6;
wire Kn4jy6, Sn4jy6, Ao4jy6, Io4jy6, Qo4jy6, Yo4jy6, Gp4jy6, Op4jy6, Wp4jy6, Eq4jy6;
wire Mq4jy6, Uq4jy6, Cr4jy6, Kr4jy6, Sr4jy6, As4jy6, Is4jy6, Qs4jy6, Ys4jy6, Gt4jy6;
wire Ot4jy6, Wt4jy6, Eu4jy6, Mu4jy6, Uu4jy6, Cv4jy6, Kv4jy6, Sv4jy6, Aw4jy6, Iw4jy6;
wire Qw4jy6, Yw4jy6, Gx4jy6, Ox4jy6, Wx4jy6, Ey4jy6, My4jy6, Uy4jy6, Cz4jy6, Kz4jy6;
wire Sz4jy6, A05jy6, I05jy6, Q05jy6, Y05jy6, G15jy6, O15jy6, W15jy6, E25jy6, M25jy6;
wire U25jy6, C35jy6, K35jy6, S35jy6, A45jy6, I45jy6, Q45jy6, Y45jy6, G55jy6, O55jy6;
wire W55jy6, E65jy6, M65jy6, U65jy6, C75jy6, K75jy6, S75jy6, A85jy6, I85jy6, Q85jy6;
wire Y85jy6, G95jy6, O95jy6, W95jy6, Ea5jy6, Ma5jy6, Ua5jy6, Cb5jy6, Kb5jy6, Sb5jy6;
wire Ac5jy6, Ic5jy6, Qc5jy6, Yc5jy6, Gd5jy6, Od5jy6, Wd5jy6, Ee5jy6, Me5jy6, Ue5jy6;
wire Cf5jy6, Kf5jy6, Sf5jy6, Ag5jy6, Ig5jy6, Qg5jy6, Yg5jy6, Gh5jy6, Oh5jy6, Wh5jy6;
wire Ei5jy6, Mi5jy6, Ui5jy6, Cj5jy6, Kj5jy6, Sj5jy6, Ak5jy6, Ik5jy6, Qk5jy6, Yk5jy6;
wire Gl5jy6, Ol5jy6, Wl5jy6, Em5jy6, Mm5jy6, Um5jy6, Cn5jy6, Kn5jy6, Sn5jy6, Ao5jy6;
wire Io5jy6, Qo5jy6, Yo5jy6, Gp5jy6, Op5jy6, Wp5jy6, Eq5jy6, Mq5jy6, Uq5jy6, Cr5jy6;
wire Kr5jy6, Sr5jy6, As5jy6, Is5jy6, Qs5jy6, Ys5jy6, Gt5jy6, Ot5jy6, Wt5jy6, Eu5jy6;
wire Mu5jy6, Uu5jy6, Cv5jy6, Kv5jy6, Sv5jy6, Aw5jy6, Iw5jy6, Qw5jy6, Yw5jy6, Gx5jy6;
wire Ox5jy6, Wx5jy6, Ey5jy6, My5jy6, Uy5jy6, Cz5jy6, Kz5jy6, Sz5jy6, A06jy6, I06jy6;
wire Q06jy6, Y06jy6, G16jy6, O16jy6, W16jy6, E26jy6, M26jy6, U26jy6, C36jy6, K36jy6;
wire S36jy6, A46jy6, I46jy6, Q46jy6, Y46jy6, G56jy6, O56jy6, W56jy6, E66jy6, M66jy6;
wire U66jy6, C76jy6, K76jy6, S76jy6, A86jy6, I86jy6, Q86jy6, Y86jy6, G96jy6, O96jy6;
wire W96jy6, Ea6jy6, Ma6jy6, Ua6jy6, Cb6jy6, Kb6jy6, Sb6jy6, Ac6jy6, Ic6jy6, Qc6jy6;
wire Yc6jy6, Gd6jy6, Od6jy6, Wd6jy6, Ee6jy6, Me6jy6, Ue6jy6, Cf6jy6, Kf6jy6, Sf6jy6;
wire Ag6jy6, Ig6jy6, Qg6jy6, Yg6jy6, Gh6jy6, Oh6jy6, Wh6jy6, Ei6jy6, Mi6jy6, Ui6jy6;
wire Cj6jy6, Kj6jy6, Sj6jy6, Ak6jy6, Ik6jy6, Qk6jy6, Yk6jy6, Gl6jy6, Ol6jy6, Wl6jy6;
wire Em6jy6, Mm6jy6, Um6jy6, Cn6jy6, Kn6jy6, Sn6jy6, Ao6jy6, Io6jy6, Qo6jy6, Yo6jy6;
wire Gp6jy6, Op6jy6, Wp6jy6, Eq6jy6, Mq6jy6, Uq6jy6, Cr6jy6, Kr6jy6, Sr6jy6, As6jy6;
wire Is6jy6, Qs6jy6, Ys6jy6, Gt6jy6, Ot6jy6, Wt6jy6, Eu6jy6, Mu6jy6, Uu6jy6, Cv6jy6;
wire Kv6jy6, Sv6jy6, Aw6jy6, Iw6jy6, Qw6jy6, Yw6jy6, Gx6jy6, Ox6jy6, Wx6jy6, Ey6jy6;
wire My6jy6, Uy6jy6, Cz6jy6, Kz6jy6, Sz6jy6, A07jy6, I07jy6, Q07jy6, Y07jy6, G17jy6;
wire O17jy6, W17jy6, E27jy6, M27jy6, U27jy6, C37jy6, K37jy6, S37jy6, A47jy6, I47jy6;
wire Q47jy6, Y47jy6, G57jy6, O57jy6, W57jy6, E67jy6, M67jy6, U67jy6, C77jy6, K77jy6;
wire S77jy6, A87jy6, I87jy6, Q87jy6, Y87jy6, G97jy6, O97jy6, W97jy6, Ea7jy6, Ma7jy6;
wire Ua7jy6, Cb7jy6, Kb7jy6, Sb7jy6, Ac7jy6, Ic7jy6, Qc7jy6, Yc7jy6, Gd7jy6, Od7jy6;
wire Wd7jy6, Ee7jy6, Me7jy6, Ue7jy6, Cf7jy6, Kf7jy6, Sf7jy6, Ag7jy6, Ig7jy6, Qg7jy6;
wire Yg7jy6, Gh7jy6, Oh7jy6, Wh7jy6, Ei7jy6, Mi7jy6, Ui7jy6, Cj7jy6, Kj7jy6, Sj7jy6;
wire Ak7jy6, Ik7jy6, Qk7jy6, Yk7jy6, Gl7jy6, Ol7jy6, Wl7jy6, Em7jy6, Mm7jy6, Um7jy6;
wire Cn7jy6, Kn7jy6, Sn7jy6, Ao7jy6, Io7jy6, Qo7jy6, Yo7jy6, Gp7jy6, Op7jy6, Wp7jy6;
wire Eq7jy6, Mq7jy6, Uq7jy6, Cr7jy6, Kr7jy6, Sr7jy6, As7jy6, Is7jy6, Qs7jy6, Ys7jy6;
wire Gt7jy6, Ot7jy6, Wt7jy6, Eu7jy6, Mu7jy6, Uu7jy6, Cv7jy6, Kv7jy6, Sv7jy6, Aw7jy6;
wire Iw7jy6, Qw7jy6, Yw7jy6, Gx7jy6, Ox7jy6, Wx7jy6, Ey7jy6, My7jy6, Uy7jy6, Cz7jy6;
wire Kz7jy6, Sz7jy6, A08jy6, I08jy6, Q08jy6, Y08jy6, G18jy6, O18jy6, W18jy6, E28jy6;
wire M28jy6, U28jy6, C38jy6, K38jy6, S38jy6, A48jy6, I48jy6, Q48jy6, Y48jy6, G58jy6;
wire O58jy6, W58jy6, E68jy6, M68jy6, U68jy6, C78jy6, K78jy6, S78jy6, A88jy6, I88jy6;
wire Q88jy6, Y88jy6, G98jy6, O98jy6, W98jy6, Ea8jy6, Ma8jy6, Ua8jy6, Cb8jy6, Kb8jy6;
wire Sb8jy6, Ac8jy6, Ic8jy6, Qc8jy6, Yc8jy6, Gd8jy6, Od8jy6, Wd8jy6, Ee8jy6, Me8jy6;
wire Ue8jy6, Cf8jy6, Kf8jy6, Sf8jy6, Ag8jy6, Ig8jy6, Qg8jy6, Yg8jy6, Gh8jy6, Oh8jy6;
wire Wh8jy6, Ei8jy6, Mi8jy6, Ui8jy6, Cj8jy6, Kj8jy6, Sj8jy6, Ak8jy6, Ik8jy6, Qk8jy6;
wire Yk8jy6, Gl8jy6, Ol8jy6, Wl8jy6, Em8jy6, Mm8jy6, Um8jy6, Cn8jy6, Kn8jy6, Sn8jy6;
wire Ao8jy6, Io8jy6, Qo8jy6, Yo8jy6, Gp8jy6, Op8jy6, Wp8jy6, Eq8jy6, Mq8jy6, Uq8jy6;
wire Cr8jy6, Kr8jy6, Sr8jy6, As8jy6, Is8jy6, Qs8jy6, Ys8jy6, Gt8jy6, Ot8jy6, Wt8jy6;
wire Eu8jy6, Mu8jy6, Uu8jy6, Cv8jy6, Kv8jy6, Sv8jy6, Aw8jy6, Iw8jy6, Qw8jy6, Yw8jy6;
wire Gx8jy6, Ox8jy6, Wx8jy6, Ey8jy6, My8jy6, Uy8jy6, Cz8jy6, Kz8jy6, Sz8jy6, A09jy6;
wire I09jy6, Q09jy6, Y09jy6, G19jy6, O19jy6, W19jy6, E29jy6, M29jy6, U29jy6, C39jy6;
wire K39jy6, S39jy6, A49jy6, I49jy6, Q49jy6, Y49jy6, G59jy6, O59jy6, W59jy6, E69jy6;
wire M69jy6, U69jy6, C79jy6, K79jy6, S79jy6, A89jy6, I89jy6, Q89jy6, Y89jy6, G99jy6;
wire O99jy6, W99jy6, Ea9jy6, Ma9jy6, Ua9jy6, Cb9jy6, Kb9jy6, Sb9jy6, Ac9jy6, Ic9jy6;
wire Qc9jy6, Yc9jy6, Gd9jy6, Od9jy6, Wd9jy6, Ee9jy6, Me9jy6, Ue9jy6, Cf9jy6, Kf9jy6;
wire Sf9jy6, Ag9jy6, Ig9jy6, Qg9jy6, Yg9jy6, Gh9jy6, Oh9jy6, Wh9jy6, Ei9jy6, Mi9jy6;
wire Ui9jy6, Cj9jy6, Kj9jy6, Sj9jy6, Ak9jy6, Ik9jy6, Qk9jy6, Yk9jy6, Gl9jy6, Ol9jy6;
wire Wl9jy6, Em9jy6, Mm9jy6, Um9jy6, Cn9jy6, Kn9jy6, Sn9jy6, Ao9jy6, Io9jy6, Qo9jy6;
wire Yo9jy6, Gp9jy6, Op9jy6, Wp9jy6, Eq9jy6, Mq9jy6, Uq9jy6, Cr9jy6, Kr9jy6, Sr9jy6;
wire As9jy6, Is9jy6, Qs9jy6, Ys9jy6, Gt9jy6, Ot9jy6, Wt9jy6, Eu9jy6, Mu9jy6, Uu9jy6;
wire Cv9jy6, Kv9jy6, Sv9jy6, Aw9jy6, Iw9jy6, Qw9jy6, Yw9jy6, Gx9jy6, Ox9jy6, Wx9jy6;
wire Ey9jy6, My9jy6, Uy9jy6, Cz9jy6, Kz9jy6, Sz9jy6, A0ajy6, I0ajy6, Q0ajy6, Y0ajy6;
wire G1ajy6, O1ajy6, W1ajy6, E2ajy6, M2ajy6, U2ajy6, C3ajy6, K3ajy6, S3ajy6, A4ajy6;
wire I4ajy6, Q4ajy6, Y4ajy6, G5ajy6, O5ajy6, W5ajy6, E6ajy6, M6ajy6, U6ajy6, C7ajy6;
wire K7ajy6, S7ajy6, A8ajy6, I8ajy6, Q8ajy6, Y8ajy6, G9ajy6, O9ajy6, W9ajy6, Eaajy6;
wire Maajy6, Uaajy6, Cbajy6, Kbajy6, Sbajy6, Acajy6, Icajy6, Qcajy6, Ycajy6, Gdajy6;
wire Odajy6, Wdajy6, Eeajy6, Meajy6, Ueajy6, Cfajy6, Kfajy6, Sfajy6, Agajy6, Igajy6;
wire Qgajy6, Ygajy6, Ghajy6, Ohajy6, Whajy6, Eiajy6, Miajy6, Uiajy6, Cjajy6, Kjajy6;
wire Sjajy6, Akajy6, Ikajy6, Qkajy6, Ykajy6, Glajy6, Olajy6, Wlajy6, Emajy6, Mmajy6;
wire Umajy6, Cnajy6, Knajy6, Snajy6, Aoajy6, Ioajy6, Qoajy6, Yoajy6, Gpajy6, Opajy6;
wire Wpajy6, Eqajy6, Mqajy6, Uqajy6, Crajy6, Krajy6, Srajy6, Asajy6, Isajy6, Qsajy6;
wire Ysajy6, Gtajy6, Otajy6, Wtajy6, Euajy6, Muajy6, Uuajy6, Cvajy6, Kvajy6, Svajy6;
wire Awajy6, Iwajy6, Qwajy6, Ywajy6, Gxajy6, Oxajy6, Wxajy6, Eyajy6, Myajy6, Uyajy6;
wire Czajy6, Kzajy6, Szajy6, A0bjy6, I0bjy6, Q0bjy6, Y0bjy6, G1bjy6, O1bjy6, W1bjy6;
wire E2bjy6, M2bjy6, U2bjy6, C3bjy6, K3bjy6, S3bjy6, A4bjy6, I4bjy6, Q4bjy6, Y4bjy6;
wire G5bjy6, O5bjy6, W5bjy6, E6bjy6, M6bjy6, U6bjy6, C7bjy6, K7bjy6, S7bjy6, A8bjy6;
wire I8bjy6, Q8bjy6, Y8bjy6, G9bjy6, O9bjy6, W9bjy6, Eabjy6, Mabjy6, Uabjy6, Cbbjy6;
wire Kbbjy6, Sbbjy6, Acbjy6, Icbjy6, Qcbjy6, Ycbjy6, Gdbjy6, Odbjy6, Wdbjy6, Eebjy6;
wire Mebjy6, Uebjy6, Cfbjy6, Kfbjy6, Sfbjy6, Agbjy6, Igbjy6, Qgbjy6, Ygbjy6, Ghbjy6;
wire Ohbjy6, Whbjy6, Eibjy6, Mibjy6, Uibjy6, Cjbjy6, Kjbjy6, Sjbjy6, Akbjy6, Ikbjy6;
wire Qkbjy6, Ykbjy6, Glbjy6, Olbjy6, Wlbjy6, Embjy6, Mmbjy6, Umbjy6, Cnbjy6, Knbjy6;
wire Snbjy6, Aobjy6, Iobjy6, Qobjy6, Yobjy6, Gpbjy6, Opbjy6, Wpbjy6, Eqbjy6, Mqbjy6;
wire Uqbjy6, Crbjy6, Krbjy6, Srbjy6, Asbjy6, Isbjy6, Qsbjy6, Ysbjy6, Gtbjy6, Otbjy6;
wire Wtbjy6, Eubjy6, Mubjy6, Uubjy6, Cvbjy6, Kvbjy6, Svbjy6, Awbjy6, Iwbjy6, Qwbjy6;
wire Ywbjy6, Gxbjy6, Oxbjy6, Wxbjy6, Eybjy6, Mybjy6, Uybjy6, Czbjy6, Kzbjy6, Szbjy6;
wire A0cjy6, I0cjy6, Q0cjy6, Y0cjy6, G1cjy6, O1cjy6, W1cjy6, E2cjy6, M2cjy6, U2cjy6;
wire C3cjy6, K3cjy6, S3cjy6, A4cjy6, I4cjy6, Q4cjy6, Y4cjy6, G5cjy6, O5cjy6, W5cjy6;
wire E6cjy6, M6cjy6, U6cjy6, C7cjy6, K7cjy6, S7cjy6, A8cjy6, I8cjy6, Q8cjy6, Y8cjy6;
wire G9cjy6, O9cjy6, W9cjy6, Eacjy6, Macjy6, Uacjy6, Cbcjy6, Kbcjy6, Sbcjy6, Accjy6;
wire Iccjy6, Qccjy6, Yccjy6, Gdcjy6, Odcjy6, Wdcjy6, Eecjy6, Mecjy6, Uecjy6, Cfcjy6;
wire Kfcjy6, Sfcjy6, Agcjy6, Igcjy6, Qgcjy6, Ygcjy6, Ghcjy6, Ohcjy6, Whcjy6, Eicjy6;
wire Micjy6, Uicjy6, Cjcjy6, Kjcjy6, Sjcjy6, Akcjy6, Ikcjy6, Qkcjy6, Ykcjy6, Glcjy6;
wire Olcjy6, Wlcjy6, Emcjy6, Mmcjy6, Umcjy6, Cncjy6, Kncjy6, Sncjy6, Aocjy6, Iocjy6;
wire Qocjy6, Yocjy6, Gpcjy6, Opcjy6, Wpcjy6, Eqcjy6, Mqcjy6, Uqcjy6, Crcjy6, Krcjy6;
wire Srcjy6, Ascjy6, Iscjy6, Qscjy6, Yscjy6, Gtcjy6, Otcjy6, Wtcjy6, Eucjy6, Mucjy6;
wire Uucjy6, Cvcjy6, Kvcjy6, Svcjy6, Awcjy6, Iwcjy6, Qwcjy6, Ywcjy6, Gxcjy6, Oxcjy6;
wire Wxcjy6, Eycjy6, Mycjy6, Uycjy6, Czcjy6, Kzcjy6, Szcjy6, A0djy6, I0djy6, Q0djy6;
wire Y0djy6, G1djy6, O1djy6, W1djy6, E2djy6, M2djy6, U2djy6, C3djy6, K3djy6, S3djy6;
wire A4djy6, I4djy6, Q4djy6, Y4djy6, G5djy6, O5djy6, W5djy6, E6djy6, M6djy6, U6djy6;
wire C7djy6, K7djy6, S7djy6, A8djy6, I8djy6, Q8djy6, Y8djy6, G9djy6, O9djy6, W9djy6;
wire Eadjy6, Madjy6, Uadjy6, Cbdjy6, Kbdjy6, Sbdjy6, Acdjy6, Icdjy6, Qcdjy6, Ycdjy6;
wire Gddjy6, Oddjy6, Wddjy6, Eedjy6, Medjy6, Uedjy6, Cfdjy6, Kfdjy6, Sfdjy6, Agdjy6;
wire Igdjy6, Qgdjy6, Ygdjy6, Ghdjy6, Ohdjy6, Whdjy6, Eidjy6, Midjy6, Uidjy6, Cjdjy6;
wire Kjdjy6, Sjdjy6, Akdjy6, Ikdjy6, Qkdjy6, Ykdjy6, Gldjy6, Oldjy6, Wldjy6, Emdjy6;
wire Mmdjy6, Umdjy6, Cndjy6, Kndjy6, Sndjy6, Aodjy6, Iodjy6, Qodjy6, Yodjy6, Gpdjy6;
wire Opdjy6, Wpdjy6, Eqdjy6, Mqdjy6, Uqdjy6, Crdjy6, Krdjy6, Srdjy6, Asdjy6, Isdjy6;
wire Qsdjy6, Ysdjy6, Gtdjy6, Otdjy6, Wtdjy6, Eudjy6, Mudjy6, Uudjy6, Cvdjy6, Kvdjy6;
wire Svdjy6, Awdjy6, Iwdjy6, Qwdjy6, Ywdjy6, Gxdjy6, Oxdjy6, Wxdjy6, Eydjy6, Mydjy6;
wire Uydjy6, Czdjy6, Kzdjy6, Szdjy6, A0ejy6, I0ejy6, Q0ejy6, Y0ejy6, G1ejy6, O1ejy6;
wire W1ejy6, E2ejy6, M2ejy6, U2ejy6, C3ejy6, K3ejy6, S3ejy6, A4ejy6, I4ejy6, Q4ejy6;
wire Y4ejy6, G5ejy6, O5ejy6, W5ejy6, E6ejy6, M6ejy6, U6ejy6, C7ejy6, K7ejy6, S7ejy6;
wire A8ejy6, I8ejy6, Q8ejy6, Y8ejy6, G9ejy6, O9ejy6, W9ejy6, Eaejy6, Maejy6, Uaejy6;
wire Cbejy6, Kbejy6, Sbejy6, Acejy6, Icejy6, Qcejy6, Ycejy6, Gdejy6, Odejy6, Wdejy6;
wire Eeejy6, Meejy6, Ueejy6, Cfejy6, Kfejy6, Sfejy6, Agejy6, Igejy6, Qgejy6, Ygejy6;
wire Ghejy6, Ohejy6, Whejy6, Eiejy6, Miejy6, Uiejy6, Cjejy6, Kjejy6, Sjejy6, Akejy6;
wire Ikejy6, Qkejy6, Ykejy6, Glejy6, Olejy6, Wlejy6, Emejy6, Mmejy6, Umejy6, Cnejy6;
wire Knejy6, Snejy6, Aoejy6, Ioejy6, Qoejy6, Yoejy6, Gpejy6, Opejy6, Wpejy6, Eqejy6;
wire Mqejy6, Uqejy6, Crejy6, Krejy6, Srejy6, Asejy6, Isejy6, Qsejy6, Ysejy6, Gtejy6;
wire Otejy6, Wtejy6, Euejy6, Muejy6, Uuejy6, Cvejy6, Kvejy6, Svejy6, Awejy6, Iwejy6;
wire Qwejy6, Ywejy6, Gxejy6, Oxejy6, Wxejy6, Eyejy6, Myejy6, Uyejy6, Czejy6, Kzejy6;
wire Szejy6, A0fjy6, I0fjy6, Q0fjy6, Y0fjy6, G1fjy6, O1fjy6, W1fjy6, E2fjy6, M2fjy6;
wire U2fjy6, C3fjy6, K3fjy6, S3fjy6, A4fjy6, I4fjy6, Q4fjy6, Y4fjy6, G5fjy6, O5fjy6;
wire W5fjy6, E6fjy6, M6fjy6, U6fjy6, C7fjy6, K7fjy6, S7fjy6, A8fjy6, I8fjy6, Q8fjy6;
wire Y8fjy6, G9fjy6, O9fjy6, W9fjy6, Eafjy6, Mafjy6, Uafjy6, Cbfjy6, Kbfjy6, Sbfjy6;
wire Acfjy6, Icfjy6, Qcfjy6, Ycfjy6, Gdfjy6, Odfjy6, Wdfjy6, Eefjy6, Mefjy6, Uefjy6;
wire Cffjy6, Kffjy6, Sffjy6, Agfjy6, Igfjy6, Qgfjy6, Ygfjy6, Ghfjy6, Ohfjy6, Whfjy6;
wire Eifjy6, Mifjy6, Uifjy6, Cjfjy6, Kjfjy6, Sjfjy6, Akfjy6, Ikfjy6, Qkfjy6, Ykfjy6;
wire Glfjy6, Olfjy6, Wlfjy6, Emfjy6, Mmfjy6, Umfjy6, Cnfjy6, Knfjy6, Snfjy6, Aofjy6;
wire Iofjy6, Qofjy6, Yofjy6, Gpfjy6, Opfjy6, Wpfjy6, Eqfjy6, Mqfjy6, Uqfjy6, Crfjy6;
wire Krfjy6, Srfjy6, Asfjy6, Isfjy6, Qsfjy6, Ysfjy6, Gtfjy6, Otfjy6, Wtfjy6, Eufjy6;
wire Mufjy6, Uufjy6, Cvfjy6, Kvfjy6, Svfjy6, Awfjy6, Iwfjy6, Qwfjy6, Ywfjy6, Gxfjy6;
wire Oxfjy6, Wxfjy6, Eyfjy6, Myfjy6, Uyfjy6, Czfjy6, Kzfjy6, Szfjy6, A0gjy6, I0gjy6;
wire Q0gjy6, Y0gjy6, G1gjy6, O1gjy6, W1gjy6, E2gjy6, M2gjy6, U2gjy6, C3gjy6, K3gjy6;
wire S3gjy6, A4gjy6, I4gjy6, Q4gjy6, Y4gjy6, G5gjy6, O5gjy6, W5gjy6, E6gjy6, M6gjy6;
wire U6gjy6, C7gjy6, K7gjy6, S7gjy6, A8gjy6, I8gjy6, Q8gjy6, Y8gjy6, G9gjy6, O9gjy6;
wire W9gjy6, Eagjy6, Magjy6, Uagjy6, Cbgjy6, Kbgjy6, Sbgjy6, Acgjy6, Icgjy6, Qcgjy6;
wire Ycgjy6, Gdgjy6, Odgjy6, Wdgjy6, Eegjy6, Megjy6, Uegjy6, Cfgjy6, Kfgjy6, Sfgjy6;
wire Aggjy6, Iggjy6, Qggjy6, Yggjy6, Ghgjy6, Ohgjy6, Whgjy6, Eigjy6, Migjy6, Uigjy6;
wire Cjgjy6, Kjgjy6, Sjgjy6, Akgjy6, Ikgjy6, Qkgjy6, Ykgjy6, Glgjy6, Olgjy6, Wlgjy6;
wire Emgjy6, Mmgjy6, Umgjy6, Cngjy6, Kngjy6, Sngjy6, Aogjy6, Iogjy6, Qogjy6, Yogjy6;
wire Gpgjy6, Opgjy6, Wpgjy6, Eqgjy6, Mqgjy6, Uqgjy6, Crgjy6, Krgjy6, Srgjy6, Asgjy6;
wire Isgjy6, Qsgjy6, Ysgjy6, Gtgjy6, Otgjy6, Wtgjy6, Eugjy6, Mugjy6, Uugjy6, Cvgjy6;
wire Kvgjy6, Svgjy6, Awgjy6, Iwgjy6, Qwgjy6, Ywgjy6, Gxgjy6, Oxgjy6, Wxgjy6, Eygjy6;
wire Mygjy6, Uygjy6, Czgjy6, Kzgjy6, Szgjy6, A0hjy6, I0hjy6, Q0hjy6, Y0hjy6, Gpu5z6;
wire Opu5z6, Wpu5z6, Equ5z6, Mqu5z6, Uqu5z6, Cru5z6, Kru5z6, Sru5z6, Asu5z6, Isu5z6;
wire Qsu5z6, Ysu5z6, Gtu5z6, Otu5z6, Wtu5z6, Euu5z6, Muu5z6, Uuu5z6, Cvu5z6, Kvu5z6;
wire Svu5z6, Awu5z6, Iwu5z6, Qwu5z6, Ywu5z6, Gxu5z6, Oxu5z6, Wxu5z6, Eyu5z6, Myu5z6;
wire Uyu5z6, Czu5z6, Kzu5z6, Szu5z6, A0v5z6, I0v5z6, Q0v5z6, Y0v5z6, G1v5z6, O1v5z6;
wire W1v5z6, E2v5z6, M2v5z6, U2v5z6, C3v5z6, K3v5z6, S3v5z6, A4v5z6, I4v5z6, Q4v5z6;
wire Y4v5z6, G5v5z6, O5v5z6, W5v5z6, E6v5z6, M6v5z6, U6v5z6, C7v5z6, K7v5z6, S7v5z6;
wire A8v5z6, I8v5z6, Q8v5z6, Y8v5z6, G9v5z6, O9v5z6, W9v5z6, Eav5z6, Mav5z6, Uav5z6;
wire Cbv5z6, Kbv5z6, Sbv5z6, Acv5z6, Icv5z6, Qcv5z6, Ycv5z6, Gdv5z6, Odv5z6, Wdv5z6;
wire Eev5z6, Mev5z6, Uev5z6, Cfv5z6, Kfv5z6, Sfv5z6, Agv5z6, Igv5z6, Qgv5z6, Ygv5z6;
wire Ghv5z6, Ohv5z6, Whv5z6, Eiv5z6, Miv5z6, Uiv5z6, Cjv5z6, Kjv5z6, Sjv5z6, Akv5z6;
wire Ikv5z6, Qkv5z6, Ykv5z6, Glv5z6, Olv5z6, Wlv5z6, Emv5z6, Mmv5z6, Umv5z6, Cnv5z6;
wire Knv5z6, Snv5z6, Aov5z6, Iov5z6, Qov5z6, Yov5z6, Gpv5z6, Opv5z6, Wpv5z6, Eqv5z6;
wire Mqv5z6, Uqv5z6, Crv5z6, Krv5z6, Srv5z6, Asv5z6, Isv5z6, Qsv5z6, Ysv5z6, Gtv5z6;
wire Otv5z6, Wtv5z6, Euv5z6, Muv5z6, Uuv5z6, Cvv5z6, Kvv5z6, Svv5z6, Awv5z6, Iwv5z6;
wire Qwv5z6, Ywv5z6, Gxv5z6, Oxv5z6, Wxv5z6, Eyv5z6, Myv5z6, Uyv5z6, Czv5z6, Kzv5z6;
wire Szv5z6, A0w5z6, I0w5z6, Q0w5z6, Y0w5z6, G1w5z6, O1w5z6, W1w5z6, E2w5z6, M2w5z6;
wire U2w5z6, C3w5z6, K3w5z6, S3w5z6, A4w5z6, I4w5z6, Q4w5z6, Y4w5z6, G5w5z6, O5w5z6;
wire W5w5z6, E6w5z6, M6w5z6, U6w5z6, C7w5z6, K7w5z6, S7w5z6, A8w5z6, I8w5z6, Q8w5z6;
wire Y8w5z6, G9w5z6, O9w5z6, W9w5z6, Eaw5z6, Maw5z6, Uaw5z6, Cbw5z6, Kbw5z6, Sbw5z6;
wire Acw5z6, Icw5z6, Qcw5z6, Ycw5z6, Gdw5z6, Odw5z6, Wdw5z6, Eew5z6, Mew5z6, Uew5z6;
wire Cfw5z6, Kfw5z6, Sfw5z6, Agw5z6, Igw5z6, Qgw5z6, Ygw5z6, Ghw5z6, Ohw5z6, Whw5z6;
wire Eiw5z6, Miw5z6, Uiw5z6, Cjw5z6, Kjw5z6, Sjw5z6, Akw5z6, Ikw5z6, Qkw5z6, Ykw5z6;
wire Glw5z6, Olw5z6, Wlw5z6, Emw5z6, Mmw5z6, Umw5z6, Cnw5z6, Knw5z6, Snw5z6, Aow5z6;
wire Iow5z6, Qow5z6, Yow5z6, Gpw5z6, Opw5z6, Wpw5z6, Eqw5z6, Mqw5z6, Uqw5z6, Crw5z6;
wire Krw5z6, Srw5z6, Asw5z6, Isw5z6, Qsw5z6, Ysw5z6, Gtw5z6, Otw5z6, Wtw5z6, Euw5z6;
wire Muw5z6, Uuw5z6, Cvw5z6, Kvw5z6, Svw5z6, Aww5z6, Iww5z6, Qww5z6, Yww5z6, Gxw5z6;
wire Oxw5z6, Wxw5z6, Eyw5z6, Myw5z6, Uyw5z6, Czw5z6, Kzw5z6, Szw5z6, A0x5z6, I0x5z6;
wire Q0x5z6, Y0x5z6, G1x5z6, O1x5z6, W1x5z6, E2x5z6, M2x5z6, U2x5z6, C3x5z6, K3x5z6;
wire S3x5z6, A4x5z6, I4x5z6, Q4x5z6, Y4x5z6, G5x5z6, O5x5z6, W5x5z6, E6x5z6, M6x5z6;
wire U6x5z6, C7x5z6, K7x5z6, S7x5z6, A8x5z6, I8x5z6, Q8x5z6, Y8x5z6, G9x5z6, O9x5z6;
wire W9x5z6, Eax5z6, Max5z6, Uax5z6, Cbx5z6, Kbx5z6, Sbx5z6, Acx5z6, Icx5z6, Qcx5z6;
wire Ycx5z6, Gdx5z6, Odx5z6, Wdx5z6, Eex5z6, Mex5z6, Uex5z6, Cfx5z6, Kfx5z6, Sfx5z6;
wire Agx5z6, Igx5z6, Qgx5z6, Ygx5z6, Ghx5z6, Ohx5z6, Whx5z6, Eix5z6, Mix5z6, Uix5z6;
wire Cjx5z6, Kjx5z6, Sjx5z6, Akx5z6, Ikx5z6, Qkx5z6, Ykx5z6, Glx5z6, Olx5z6, Wlx5z6;
wire Emx5z6, Mmx5z6, Umx5z6, Cnx5z6, Knx5z6, Snx5z6, Aox5z6, Iox5z6, Qox5z6, Yox5z6;
wire Gpx5z6, Opx5z6, Wpx5z6, Eqx5z6, Mqx5z6, Uqx5z6, Crx5z6, Krx5z6, Srx5z6, Asx5z6;
wire Isx5z6, Qsx5z6, Ysx5z6, Gtx5z6, Otx5z6, Wtx5z6, Eux5z6, Mux5z6, Uux5z6, Cvx5z6;
wire Kvx5z6, Svx5z6, Awx5z6, Iwx5z6, Qwx5z6, Ywx5z6, Gxx5z6, Oxx5z6, Wxx5z6, Eyx5z6;
wire Myx5z6, Uyx5z6, Czx5z6, Kzx5z6, Szx5z6, A0y5z6, I0y5z6, Q0y5z6, Y0y5z6, G1y5z6;
wire O1y5z6, W1y5z6, E2y5z6, M2y5z6, U2y5z6, C3y5z6, K3y5z6, S3y5z6, A4y5z6, I4y5z6;
wire Q4y5z6, Y4y5z6, G5y5z6, O5y5z6, W5y5z6, E6y5z6, M6y5z6, U6y5z6, C7y5z6, K7y5z6;
wire S7y5z6, A8y5z6, I8y5z6, Q8y5z6, Y8y5z6, G9y5z6, O9y5z6, W9y5z6, Eay5z6, May5z6;
wire Uay5z6, Cby5z6, Kby5z6, Sby5z6, Acy5z6, Icy5z6, Qcy5z6, Ycy5z6, Gdy5z6, Ody5z6;
wire Wdy5z6, Eey5z6, Mey5z6, Uey5z6, Cfy5z6, Kfy5z6, Sfy5z6, Agy5z6, Igy5z6, Qgy5z6;
wire Ygy5z6, Ghy5z6, Ohy5z6, Why5z6, Eiy5z6, Miy5z6, Uiy5z6, Cjy5z6, Kjy5z6, Sjy5z6;
wire Aky5z6, Iky5z6, Qky5z6, Yky5z6, Gly5z6, Oly5z6, Wly5z6, Emy5z6, Mmy5z6, Umy5z6;
wire Cny5z6, Kny5z6, Sny5z6, Aoy5z6, Ioy5z6, Qoy5z6, Yoy5z6, Gpy5z6, Opy5z6, Wpy5z6;
wire Eqy5z6, Mqy5z6, Uqy5z6, Cry5z6, Kry5z6, Sry5z6, Asy5z6, Isy5z6, Qsy5z6, Ysy5z6;
wire Gty5z6, Oty5z6, Wty5z6, Euy5z6, Muy5z6, Uuy5z6, Cvy5z6, Kvy5z6, Svy5z6, Awy5z6;
wire Iwy5z6, Qwy5z6, Ywy5z6, Gxy5z6, Oxy5z6, Wxy5z6, Eyy5z6, Myy5z6, Uyy5z6, Czy5z6;
wire Kzy5z6, Szy5z6, A0z5z6, I0z5z6, Q0z5z6, Y0z5z6, G1z5z6, O1z5z6, W1z5z6, E2z5z6;
wire M2z5z6, U2z5z6, C3z5z6, K3z5z6, S3z5z6, A4z5z6, I4z5z6, Q4z5z6, Y4z5z6, G5z5z6;
wire O5z5z6, W5z5z6, E6z5z6, M6z5z6, U6z5z6, C7z5z6, K7z5z6, S7z5z6, A8z5z6, I8z5z6;
wire Q8z5z6, Y8z5z6, G9z5z6, O9z5z6, W9z5z6, Eaz5z6, Maz5z6, Uaz5z6, Cbz5z6, Kbz5z6;
wire Sbz5z6, Acz5z6, Icz5z6, Qcz5z6, Ycz5z6, Gdz5z6, Odz5z6, Wdz5z6, Eez5z6, Mez5z6;
wire Uez5z6, Cfz5z6, Kfz5z6, Sfz5z6, Agz5z6, Igz5z6, Qgz5z6, Ygz5z6, Ghz5z6, Ohz5z6;
wire Whz5z6, Eiz5z6, Miz5z6, Uiz5z6, Cjz5z6, Kjz5z6, Sjz5z6, Akz5z6, Ikz5z6, Qkz5z6;
wire Ykz5z6, Glz5z6, Olz5z6, Wlz5z6, Emz5z6, Mmz5z6, Umz5z6, Cnz5z6, Knz5z6, Snz5z6;
wire Aoz5z6, Ioz5z6, Qoz5z6, Yoz5z6, Gpz5z6, Opz5z6, Wpz5z6, Eqz5z6, Mqz5z6, Uqz5z6;
wire Crz5z6, Krz5z6, Srz5z6, Asz5z6, Isz5z6, Qsz5z6, Ysz5z6, Gtz5z6, Otz5z6, Wtz5z6;
wire Euz5z6, Muz5z6, Uuz5z6, Cvz5z6, Kvz5z6, Svz5z6, Awz5z6, Iwz5z6, Qwz5z6, Ywz5z6;
wire Gxz5z6, Oxz5z6, Wxz5z6, Eyz5z6, Myz5z6, Uyz5z6, Czz5z6, Kzz5z6, Szz5z6, A006z6;
wire I006z6, Q006z6, Y006z6, G106z6, O106z6, W106z6, E206z6, M206z6, U206z6, C306z6;
wire K306z6, S306z6, A406z6, I406z6, Q406z6, Y406z6, G506z6, O506z6, W506z6, E606z6;
wire M606z6, U606z6, C706z6, K706z6, S706z6, A806z6, I806z6, Q806z6, Y806z6, G906z6;
wire O906z6, W906z6, Ea06z6, Ma06z6, Ua06z6, Cb06z6, Kb06z6, Sb06z6, Ac06z6, Ic06z6;
wire Qc06z6, Yc06z6, Gd06z6, Od06z6, Wd06z6, Ee06z6, Me06z6, Ue06z6, Cf06z6, Kf06z6;
wire Sf06z6, Ag06z6, Ig06z6, Qg06z6, Yg06z6, Gh06z6, Oh06z6, Wh06z6, Ei06z6, Mi06z6;
wire Ui06z6, Cj06z6, Kj06z6, Sj06z6, Ak06z6, Ik06z6, Qk06z6, Yk06z6, Gl06z6, Ol06z6;
wire Wl06z6, Em06z6, Mm06z6, Um06z6, Cn06z6, Kn06z6, Sn06z6, Ao06z6, Io06z6, Qo06z6;
wire Yo06z6, Gp06z6, Op06z6, Wp06z6, Eq06z6, Mq06z6, Uq06z6, Cr06z6, Kr06z6, Sr06z6;
wire As06z6, Is06z6, Qs06z6, Ys06z6, Gt06z6, Ot06z6, Wt06z6, Eu06z6, Mu06z6, Uu06z6;
wire Cv06z6, Kv06z6, Sv06z6, Aw06z6, Iw06z6, Qw06z6, Yw06z6, Gx06z6, Ox06z6, Wx06z6;
wire Ey06z6, My06z6, Uy06z6, Cz06z6, Kz06z6, Sz06z6, A016z6, I016z6, Q016z6, Y016z6;
wire G116z6, O116z6, W116z6, E216z6, M216z6, U216z6, C316z6, K316z6, S316z6, A416z6;
wire I416z6, Q416z6, Y416z6, G516z6, O516z6, W516z6, E616z6, M616z6, U616z6, C716z6;
wire K716z6, S716z6, A816z6, I816z6, Q816z6, Y816z6, G916z6, O916z6, W916z6, Ea16z6;
wire Ma16z6, Ua16z6, Cb16z6, Kb16z6, Sb16z6, Ac16z6, Ic16z6, Qc16z6, Yc16z6, Gd16z6;
wire Od16z6, Wd16z6, Ee16z6, Me16z6, Ue16z6, Cf16z6, Kf16z6, Sf16z6, Ag16z6, Ig16z6;
wire Qg16z6, Yg16z6, Gh16z6, Oh16z6, Wh16z6, Ei16z6, Mi16z6, Ui16z6, Cj16z6, Kj16z6;
wire Sj16z6, Ak16z6, Ik16z6, Qk16z6, Yk16z6, Gl16z6, Ol16z6, Wl16z6, Em16z6, Mm16z6;
wire Um16z6, Cn16z6, Kn16z6, Sn16z6, Ao16z6, Io16z6, Qo16z6, Yo16z6, Gp16z6, Op16z6;
wire Wp16z6, Eq16z6, Mq16z6, Uq16z6, Cr16z6, Kr16z6, Sr16z6, As16z6, Is16z6, Qs16z6;
wire Ys16z6, Gt16z6, Ot16z6, Wt16z6, Eu16z6, Mu16z6, Uu16z6, Cv16z6, Kv16z6, Sv16z6;
wire Aw16z6, Iw16z6, Qw16z6, Yw16z6, Gx16z6, Ox16z6, Wx16z6, Ey16z6, My16z6, Uy16z6;
wire Cz16z6, Kz16z6, Sz16z6, A026z6, I026z6, Q026z6, Y026z6, G126z6, O126z6, W126z6;
wire E226z6, M226z6, U226z6, C326z6, K326z6, S326z6, A426z6, I426z6, Q426z6, Y426z6;
wire G526z6, O526z6, W526z6, E626z6, M626z6, U626z6, C726z6, K726z6, S726z6, A826z6;
wire I826z6, Q826z6, Y826z6, G926z6, O926z6, W926z6, Ea26z6, Ma26z6, Ua26z6, Cb26z6;
wire Kb26z6, Sb26z6, Ac26z6, Ic26z6, Qc26z6, Yc26z6, Gd26z6, Od26z6, Wd26z6, Ee26z6;
wire Me26z6, Ue26z6, Cf26z6, Kf26z6, Sf26z6, Ag26z6, Ig26z6, Qg26z6, Yg26z6, Gh26z6;
wire Oh26z6, Wh26z6, Ei26z6, Mi26z6, Ui26z6, Cj26z6, Kj26z6, Sj26z6, Ak26z6, Ik26z6;
wire Qk26z6, Yk26z6, Gl26z6, Ol26z6, Wl26z6, Em26z6, Mm26z6, Um26z6, Cn26z6, Kn26z6;
wire Sn26z6, Ao26z6, Io26z6, Qo26z6, Yo26z6, Gp26z6, Op26z6, Wp26z6, Eq26z6, Mq26z6;
wire Uq26z6, Cr26z6, Kr26z6, Sr26z6, As26z6, Is26z6, Qs26z6, Ys26z6, Gt26z6, Ot26z6;
wire Wt26z6, Eu26z6, Mu26z6, Uu26z6, Cv26z6, Kv26z6, Sv26z6, Aw26z6, Iw26z6, Qw26z6;
wire Yw26z6, Gx26z6, Ox26z6, Wx26z6, Ey26z6, My26z6, Uy26z6, Cz26z6, Kz26z6, Sz26z6;
wire A036z6, I036z6, Q036z6, Y036z6, G136z6, O136z6, W136z6, E236z6, M236z6, U236z6;
wire C336z6, K336z6, S336z6, A436z6, I436z6, Q436z6, Y436z6, G536z6, O536z6, W536z6;
wire E636z6, M636z6, U636z6, C736z6, K736z6, S736z6, A836z6, I836z6, Q836z6, Y836z6;
wire G936z6, O936z6, W936z6, Ea36z6, Ma36z6, Ua36z6, Cb36z6, Kb36z6, Sb36z6, Ac36z6;
wire Ic36z6, Qc36z6, Yc36z6, Gd36z6, Od36z6, Wd36z6, Ee36z6, Me36z6, Ue36z6, Cf36z6;
wire Kf36z6, Sf36z6, Ag36z6, Ig36z6, Qg36z6, Yg36z6, Gh36z6, Oh36z6, Wh36z6, Ei36z6;
wire Mi36z6, Ui36z6, Cj36z6, Kj36z6, Sj36z6, Ak36z6, Ik36z6, Qk36z6, Yk36z6, Gl36z6;
wire Ol36z6, Wl36z6, Em36z6, Mm36z6, Um36z6, Cn36z6, Kn36z6, Sn36z6, Ao36z6, Io36z6;
wire Qo36z6, Yo36z6, Gp36z6, Op36z6, Wp36z6, Eq36z6, Mq36z6, Uq36z6, Cr36z6, Kr36z6;
wire Sr36z6, As36z6, Is36z6, Qs36z6, Ys36z6, Gt36z6, Ot36z6, Wt36z6, Eu36z6, Mu36z6;
wire Uu36z6, Cv36z6, Kv36z6, Sv36z6, Aw36z6, Iw36z6, Qw36z6, Yw36z6, Gx36z6, Ox36z6;
wire Wx36z6, Ey36z6, My36z6, Uy36z6, Cz36z6, Kz36z6, Sz36z6, A046z6, I046z6, Q046z6;
wire Y046z6, G146z6, O146z6, W146z6, E246z6, M246z6, U246z6, C346z6, K346z6, S346z6;
wire A446z6, I446z6, Q446z6, Y446z6, G546z6, O546z6, W546z6, E646z6, M646z6, U646z6;
wire C746z6, K746z6, S746z6, A846z6, I846z6, Q846z6, Y846z6, G946z6, O946z6, W946z6;
wire Ea46z6, Ma46z6, Ua46z6, Cb46z6, Kb46z6, Sb46z6, Ac46z6, Ic46z6, Qc46z6, Yc46z6;
wire Gd46z6, Od46z6, Wd46z6, Ee46z6, Me46z6, Ue46z6, Cf46z6, Kf46z6, Sf46z6, Ag46z6;
wire Ig46z6, Qg46z6, Yg46z6, Gh46z6, Oh46z6, Wh46z6, Ei46z6, Mi46z6, Ui46z6, Cj46z6;
wire Kj46z6, Sj46z6, Ak46z6, Ik46z6, Qk46z6, Yk46z6, Gl46z6, Ol46z6, Wl46z6, Em46z6;
wire Mm46z6, Um46z6, Cn46z6, Kn46z6, Sn46z6, Ao46z6, Io46z6, Qo46z6, Yo46z6, Gp46z6;
wire Op46z6, Wp46z6, Eq46z6, Mq46z6, Uq46z6, Cr46z6, Kr46z6, Sr46z6, As46z6, Is46z6;
wire Qs46z6, Ys46z6, Gt46z6, Ot46z6, Wt46z6, Eu46z6, Mu46z6, Uu46z6, Cv46z6, Kv46z6;
wire Sv46z6, Aw46z6, Iw46z6, Qw46z6, Yw46z6, Gx46z6, Ox46z6, Wx46z6, Ey46z6, My46z6;
wire Uy46z6, Cz46z6, Kz46z6, Sz46z6, A056z6, I056z6, Q056z6, Y056z6, G156z6, O156z6;
wire W156z6, E256z6, M256z6, U256z6, C356z6, K356z6, S356z6, A456z6, I456z6, Q456z6;
wire Y456z6, G556z6, O556z6, W556z6, E656z6, M656z6, U656z6, C756z6, K756z6, S756z6;
wire A856z6, I856z6, Q856z6, Y856z6, G956z6, O956z6, W956z6, Ea56z6, Ma56z6, Ua56z6;
wire Cb56z6, Kb56z6, Sb56z6, Ac56z6, Ic56z6, Qc56z6, Yc56z6, Gd56z6, Od56z6, Wd56z6;
wire Ee56z6, Me56z6, Ue56z6, Cf56z6, Kf56z6, Sf56z6, Ag56z6, Ig56z6, Qg56z6, Yg56z6;
wire Gh56z6, Oh56z6, Wh56z6, Ei56z6, Mi56z6, Ui56z6, Cj56z6, Kj56z6, Sj56z6, Ak56z6;
wire Ik56z6, Qk56z6, Yk56z6, Gl56z6, Ol56z6, Wl56z6, Em56z6, Mm56z6, Um56z6, Cn56z6;
wire Kn56z6, Sn56z6, Ao56z6, Io56z6, Qo56z6, Yo56z6, Gp56z6, Op56z6, Wp56z6, Eq56z6;
wire Mq56z6, Uq56z6, Cr56z6, Kr56z6, Sr56z6, As56z6, Is56z6, Qs56z6, Ys56z6, Gt56z6;
wire Ot56z6, Wt56z6, Eu56z6, Mu56z6, Uu56z6, Cv56z6, Kv56z6, Sv56z6, Aw56z6, Iw56z6;
wire Qw56z6, Yw56z6, Gx56z6, Ox56z6, Wx56z6, Ey56z6, My56z6, Uy56z6, Cz56z6, Kz56z6;
wire Sz56z6, A066z6, I066z6, Q066z6, Y066z6, G166z6, O166z6, W166z6, E266z6, M266z6;
wire U266z6, C366z6, K366z6, S366z6, A466z6, I466z6, Q466z6, Y466z6, G566z6, O566z6;
wire W566z6, E666z6, M666z6, U666z6, C766z6, K766z6, S766z6, A866z6, I866z6, Q866z6;
wire Y866z6, G966z6, O966z6, W966z6, Ea66z6, Ma66z6, Ua66z6, Cb66z6, Kb66z6, Sb66z6;
wire Ac66z6, Ic66z6, Qc66z6, Yc66z6, Gd66z6, Od66z6, Wd66z6, Ee66z6, Me66z6, Ue66z6;
wire Cf66z6, Kf66z6, Sf66z6, Ag66z6, Ig66z6, Qg66z6, Yg66z6, Gh66z6, Oh66z6, Wh66z6;
wire Ei66z6, Mi66z6, Ui66z6, Cj66z6, Kj66z6, Sj66z6, Ak66z6, Ik66z6, Qk66z6, Yk66z6;
wire Gl66z6, Ol66z6, Wl66z6, Em66z6, Mm66z6, Um66z6, Cn66z6, Kn66z6, Sn66z6, Ao66z6;
wire Io66z6, Qo66z6, Yo66z6, Gp66z6, Op66z6, Wp66z6, Eq66z6, Mq66z6, Uq66z6, Cr66z6;
wire Kr66z6, Sr66z6, As66z6, Is66z6, Qs66z6, Ys66z6, Gt66z6, Ot66z6, Wt66z6, Eu66z6;
wire Mu66z6, Uu66z6, Cv66z6, Kv66z6, Sv66z6, Aw66z6, Iw66z6, Qw66z6, Yw66z6, Gx66z6;
wire Ox66z6, Wx66z6, Ey66z6, My66z6, Uy66z6, Cz66z6, Kz66z6, Sz66z6, A076z6, I076z6;
wire Q076z6, Y076z6, G176z6, O176z6, W176z6, E276z6, M276z6, U276z6, C376z6, K376z6;
wire S376z6, A476z6, I476z6, Q476z6, Y476z6, G576z6, O576z6, W576z6, E676z6, M676z6;
wire U676z6, C776z6, K776z6, S776z6, A876z6, I876z6, Q876z6, Y876z6, G976z6, O976z6;
wire W976z6, Ea76z6, Ma76z6, Ua76z6, Cb76z6, Kb76z6, Sb76z6, Ac76z6, Ic76z6, Qc76z6;
wire Yc76z6, Gd76z6, Od76z6, Wd76z6, Ee76z6, Me76z6, Ue76z6, Cf76z6, Kf76z6, Sf76z6;
wire Ag76z6, Ig76z6, Qg76z6, Yg76z6, Gh76z6, Oh76z6, Wh76z6, Ei76z6, Mi76z6, Ui76z6;
wire Cj76z6, Kj76z6, Sj76z6, Ak76z6, Ik76z6, Qk76z6, Yk76z6, Gl76z6, Ol76z6, Wl76z6;
wire Em76z6, Mm76z6, Um76z6, Cn76z6, Kn76z6, Sn76z6, Ao76z6, Io76z6, Qo76z6, Yo76z6;
wire Gp76z6, Op76z6, Wp76z6, Eq76z6, Mq76z6, Uq76z6, Cr76z6, Kr76z6, Sr76z6, As76z6;
wire Is76z6, Qs76z6, Ys76z6, Gt76z6, Ot76z6, Wt76z6, Eu76z6, Mu76z6, Uu76z6, Cv76z6;
wire Kv76z6, Sv76z6, Aw76z6, Iw76z6, Qw76z6, Yw76z6, Gx76z6, Ox76z6, Wx76z6, Ey76z6;
wire My76z6, Uy76z6, Cz76z6, Kz76z6, Sz76z6, A086z6, I086z6, Q086z6, Y086z6, G186z6;
wire O186z6, W186z6, E286z6, M286z6, U286z6, C386z6, K386z6, S386z6, A486z6, I486z6;
wire Q486z6, Y486z6, G586z6, O586z6, W586z6, E686z6, M686z6, U686z6, C786z6, K786z6;
wire S786z6, A886z6, I886z6, Q886z6, Y886z6, G986z6, O986z6, W986z6, Ea86z6, Ma86z6;
wire Ua86z6, Cb86z6, Kb86z6, Sb86z6, Ac86z6, Ic86z6, Qc86z6, Yc86z6, Gd86z6, Od86z6;
wire Wd86z6, Ee86z6, Me86z6, Ue86z6, Cf86z6, Kf86z6, Sf86z6, Ag86z6, Ig86z6, Qg86z6;
wire Yg86z6, Gh86z6, Oh86z6, Wh86z6, Ei86z6, Mi86z6, Ui86z6, Cj86z6, Kj86z6, Sj86z6;
wire Ak86z6, Ik86z6, Qk86z6, Yk86z6, Gl86z6, Ol86z6, Wl86z6, Em86z6, Mm86z6, Um86z6;
wire Cn86z6, Kn86z6, Sn86z6, Ao86z6, Io86z6, Qo86z6, Yo86z6, Gp86z6, Op86z6, Wp86z6;
wire Eq86z6, Mq86z6, Uq86z6, Cr86z6, Kr86z6, Sr86z6, As86z6, Is86z6, Qs86z6, Ys86z6;
wire Gt86z6, Ot86z6, Wt86z6, Eu86z6, Mu86z6, Uu86z6, Cv86z6, Kv86z6, Sv86z6, Aw86z6;
wire Iw86z6, Qw86z6, Yw86z6, Gx86z6, Ox86z6, Wx86z6, Ey86z6, My86z6, Uy86z6, Cz86z6;
wire Kz86z6, Sz86z6, A096z6, I096z6, Q096z6, Y096z6, G196z6, O196z6, W196z6, E296z6;
wire M296z6, U296z6, C396z6, K396z6, S396z6, A496z6, I496z6, Q496z6, Y496z6, G596z6;
wire O596z6, W596z6, E696z6, M696z6, U696z6, C796z6, K796z6, S796z6, A896z6, I896z6;
wire Q896z6, Y896z6, G996z6, O996z6, W996z6, Ea96z6, Ma96z6, Ua96z6, Cb96z6, Kb96z6;
wire Sb96z6, Ac96z6, Ic96z6, Qc96z6, Yc96z6, Gd96z6, Od96z6, Wd96z6, Ee96z6, Me96z6;
wire Ue96z6, Cf96z6, Kf96z6, Sf96z6, Ag96z6, Ig96z6, Qg96z6, Yg96z6, Gh96z6, Oh96z6;
wire Wh96z6, Ei96z6, Mi96z6, Ui96z6, Cj96z6, Kj96z6, Sj96z6, Ak96z6, Ik96z6, Qk96z6;
wire Yk96z6, Gl96z6, Ol96z6, Wl96z6, Em96z6, Mm96z6, Um96z6, Cn96z6, Kn96z6, Sn96z6;
wire Ao96z6, Io96z6, Qo96z6, Yo96z6, Gp96z6, Op96z6, Wp96z6, Eq96z6, Mq96z6, Uq96z6;
wire Cr96z6, Kr96z6, Sr96z6, As96z6, Is96z6, Qs96z6, Ys96z6, Gt96z6, Ot96z6, Wt96z6;
wire Eu96z6, Mu96z6, Uu96z6, Cv96z6, Kv96z6, Sv96z6, Aw96z6, Iw96z6, Qw96z6, Yw96z6;
wire Gx96z6, Ox96z6, Wx96z6, Ey96z6, My96z6, Uy96z6, Cz96z6, Kz96z6, Sz96z6, A0a6z6;
wire I0a6z6, Q0a6z6, Y0a6z6, G1a6z6, O1a6z6, W1a6z6, E2a6z6, M2a6z6, U2a6z6, C3a6z6;
wire K3a6z6, S3a6z6, A4a6z6, I4a6z6, Q4a6z6, Y4a6z6, G5a6z6, O5a6z6, W5a6z6, E6a6z6;
wire M6a6z6, U6a6z6, C7a6z6, K7a6z6, S7a6z6, A8a6z6, I8a6z6, Q8a6z6, Y8a6z6, G9a6z6;
wire O9a6z6, W9a6z6, Eaa6z6, Maa6z6, Uaa6z6, Cba6z6, Kba6z6, Sba6z6, Aca6z6, Ica6z6;
wire Qca6z6, Yca6z6, Gda6z6, Oda6z6, Wda6z6, Eea6z6, Mea6z6, Uea6z6, Cfa6z6, Kfa6z6;
wire Sfa6z6, Aga6z6, Iga6z6, Qga6z6, Yga6z6, Gha6z6, Oha6z6, Wha6z6, Eia6z6, Mia6z6;
wire Uia6z6, Cja6z6, Kja6z6, Sja6z6, Aka6z6, Ika6z6, Qka6z6, Yka6z6, Gla6z6, Ola6z6;
wire Wla6z6, Ema6z6, Mma6z6, Uma6z6, Cna6z6, Kna6z6, Sna6z6, Aoa6z6, Ioa6z6, Qoa6z6;
wire Yoa6z6, Gpa6z6, Opa6z6, Wpa6z6, Eqa6z6, Mqa6z6, Uqa6z6, Cra6z6, Kra6z6, Sra6z6;
wire Asa6z6, Isa6z6, Qsa6z6, Ysa6z6, Gta6z6, Ota6z6, Wta6z6, Eua6z6, Mua6z6, Uua6z6;
wire Cva6z6, Kva6z6, Sva6z6, Awa6z6, Iwa6z6, Qwa6z6, Ywa6z6, Gxa6z6, Oxa6z6, Wxa6z6;
wire Eya6z6, Mya6z6, Uya6z6, Cza6z6, Kza6z6, Sza6z6, A0b6z6, I0b6z6, Q0b6z6, Y0b6z6;
wire G1b6z6, O1b6z6, W1b6z6, E2b6z6, M2b6z6, U2b6z6, C3b6z6, K3b6z6, S3b6z6, A4b6z6;
wire I4b6z6, Q4b6z6, Y4b6z6, G5b6z6, O5b6z6, W5b6z6, E6b6z6, M6b6z6, U6b6z6, C7b6z6;
wire K7b6z6, S7b6z6, A8b6z6, I8b6z6, Q8b6z6, Y8b6z6, G9b6z6, O9b6z6, W9b6z6, Eab6z6;
wire Mab6z6, Uab6z6, Cbb6z6, Kbb6z6, Sbb6z6, Acb6z6, Icb6z6, Qcb6z6, Ycb6z6, Gdb6z6;
wire Odb6z6, Wdb6z6, Eeb6z6, Meb6z6, Ueb6z6, Cfb6z6, Kfb6z6, Sfb6z6, Agb6z6, Igb6z6;
wire Qgb6z6, Ygb6z6, Ghb6z6, Ohb6z6, Whb6z6, Eib6z6, Mib6z6, Uib6z6, Cjb6z6, Kjb6z6;
wire Sjb6z6, Akb6z6, Ikb6z6, Qkb6z6, Ykb6z6, Glb6z6, Olb6z6, Wlb6z6, Emb6z6, Mmb6z6;
wire Umb6z6, Cnb6z6, Knb6z6, Snb6z6, Aob6z6, Iob6z6, Qob6z6, Yob6z6, Gpb6z6, Opb6z6;
wire Wpb6z6, Eqb6z6, Mqb6z6, Uqb6z6, Crb6z6, Krb6z6, Srb6z6, Asb6z6, Isb6z6, Qsb6z6;
wire Ysb6z6, Gtb6z6, Otb6z6, Wtb6z6, Eub6z6, Mub6z6, Uub6z6, Cvb6z6, Kvb6z6, Svb6z6;
wire Awb6z6, Iwb6z6, Qwb6z6, Ywb6z6, Gxb6z6, Oxb6z6, Wxb6z6, Eyb6z6, Myb6z6, Uyb6z6;
wire Czb6z6, Kzb6z6, Szb6z6, A0c6z6, I0c6z6, Q0c6z6, Y0c6z6, G1c6z6, O1c6z6, W1c6z6;
wire E2c6z6, M2c6z6, U2c6z6, C3c6z6, K3c6z6, S3c6z6, A4c6z6, I4c6z6, Q4c6z6, Y4c6z6;
wire G5c6z6, O5c6z6, W5c6z6, E6c6z6, M6c6z6, U6c6z6, C7c6z6, K7c6z6, S7c6z6, A8c6z6;
wire I8c6z6, Q8c6z6, Y8c6z6, G9c6z6, O9c6z6, W9c6z6, Eac6z6, Mac6z6, Uac6z6, Cbc6z6;
wire Kbc6z6, Sbc6z6, Acc6z6, Icc6z6, Qcc6z6, Ycc6z6, Gdc6z6, Odc6z6, Wdc6z6, Eec6z6;
wire Mec6z6, Uec6z6, Cfc6z6, Kfc6z6, Sfc6z6, Agc6z6, Igc6z6, Qgc6z6, Ygc6z6, Ghc6z6;
wire Ohc6z6, Whc6z6, Eic6z6, Mic6z6, Uic6z6, Cjc6z6, Kjc6z6, Sjc6z6, Akc6z6, Ikc6z6;
wire Qkc6z6, Ykc6z6, Glc6z6, Olc6z6, Wlc6z6, Emc6z6, Mmc6z6, Umc6z6, Cnc6z6, Knc6z6;
wire Snc6z6, Aoc6z6, Ioc6z6, Qoc6z6, Yoc6z6, Gpc6z6, Opc6z6, Wpc6z6, Eqc6z6, Mqc6z6;
wire Uqc6z6, Crc6z6, Krc6z6, Src6z6, Asc6z6, Isc6z6, Qsc6z6, Ysc6z6, Gtc6z6, Otc6z6;
wire Wtc6z6, Euc6z6, Muc6z6, Uuc6z6, Cvc6z6, Kvc6z6, Svc6z6, Awc6z6, Iwc6z6, Qwc6z6;
wire Ywc6z6, Gxc6z6, Oxc6z6, Wxc6z6, Eyc6z6, Myc6z6, Uyc6z6, Czc6z6, Kzc6z6, Szc6z6;
wire A0d6z6, I0d6z6, Q0d6z6, Y0d6z6, G1d6z6, O1d6z6, W1d6z6, E2d6z6, M2d6z6, U2d6z6;
wire C3d6z6, K3d6z6, S3d6z6, A4d6z6, I4d6z6, Q4d6z6, Y4d6z6, G5d6z6, O5d6z6, W5d6z6;
wire E6d6z6, M6d6z6, U6d6z6, C7d6z6, K7d6z6, S7d6z6, A8d6z6, I8d6z6, Q8d6z6, Y8d6z6;
wire G9d6z6, O9d6z6, W9d6z6, Ead6z6, Mad6z6, Uad6z6, Cbd6z6, Kbd6z6, Sbd6z6, Acd6z6;
wire Icd6z6, Qcd6z6, Ycd6z6, Gdd6z6, Odd6z6, Wdd6z6, Eed6z6, Med6z6, Ued6z6, Cfd6z6;
wire Kfd6z6, Sfd6z6, Agd6z6, Igd6z6, Qgd6z6, Ygd6z6, Ghd6z6, Ohd6z6, Whd6z6, Eid6z6;
wire Mid6z6, Uid6z6, Cjd6z6, Kjd6z6, Sjd6z6, Akd6z6, Ikd6z6, Qkd6z6, Ykd6z6, Gld6z6;
wire Old6z6, Wld6z6, Emd6z6, Mmd6z6, Umd6z6, Cnd6z6, Knd6z6, Snd6z6, Aod6z6, Iod6z6;
wire Qod6z6, Yod6z6, Gpd6z6, Opd6z6, Wpd6z6, Eqd6z6, Mqd6z6, Uqd6z6, Crd6z6, Krd6z6;
wire Srd6z6, Asd6z6, Isd6z6, Qsd6z6, Ysd6z6, Gtd6z6, Otd6z6, Wtd6z6, Eud6z6, Mud6z6;
wire Uud6z6, Cvd6z6, Kvd6z6, Svd6z6, Awd6z6, Iwd6z6, Qwd6z6, Ywd6z6, Gxd6z6, Oxd6z6;
wire Wxd6z6, Eyd6z6, Myd6z6, Uyd6z6, Czd6z6, Kzd6z6, Szd6z6, A0e6z6, I0e6z6, Q0e6z6;
wire Y0e6z6, G1e6z6, O1e6z6, W1e6z6, E2e6z6, M2e6z6, U2e6z6, C3e6z6, K3e6z6, S3e6z6;
wire A4e6z6, I4e6z6, Q4e6z6, Y4e6z6, G5e6z6, O5e6z6, W5e6z6, E6e6z6, M6e6z6, U6e6z6;
wire C7e6z6, K7e6z6, S7e6z6, A8e6z6, I8e6z6, Q8e6z6, Y8e6z6, G9e6z6, O9e6z6, W9e6z6;
wire Eae6z6, Mae6z6, Uae6z6, Cbe6z6, Kbe6z6, Sbe6z6, Ace6z6, Ice6z6, Qce6z6, Yce6z6;
wire Gde6z6, Ode6z6, Wde6z6, Eee6z6, Mee6z6, Uee6z6, Cfe6z6, Kfe6z6, Sfe6z6, Age6z6;
wire Ige6z6, Qge6z6, Yge6z6, Ghe6z6, Ohe6z6, Whe6z6, Eie6z6, Mie6z6, Uie6z6, Cje6z6;
wire Kje6z6, Sje6z6, Ake6z6, Ike6z6, Qke6z6, Yke6z6, Gle6z6, Ole6z6, Wle6z6, Eme6z6;
wire Mme6z6, Ume6z6, Cne6z6, Kne6z6, Sne6z6, Aoe6z6, Ioe6z6, Qoe6z6, Yoe6z6, Gpe6z6;
wire Ope6z6, Wpe6z6, Eqe6z6, Mqe6z6, Uqe6z6, Cre6z6, Kre6z6, Sre6z6, Ase6z6, Ise6z6;
wire Qse6z6, Yse6z6, Gte6z6, Ote6z6, Wte6z6, Eue6z6, Mue6z6, Uue6z6, Cve6z6, Kve6z6;
wire Sve6z6, Awe6z6, Iwe6z6, Qwe6z6, Ywe6z6, Gxe6z6, Oxe6z6, Wxe6z6, Eye6z6, Mye6z6;
wire Uye6z6, Cze6z6, Kze6z6, Sze6z6, A0f6z6, I0f6z6, Q0f6z6, Y0f6z6, G1f6z6, O1f6z6;
wire W1f6z6, E2f6z6, M2f6z6, U2f6z6, C3f6z6, K3f6z6, S3f6z6, A4f6z6, I4f6z6, Q4f6z6;
wire Y4f6z6, G5f6z6, O5f6z6, W5f6z6, E6f6z6, M6f6z6, U6f6z6, C7f6z6, K7f6z6, S7f6z6;
wire A8f6z6, I8f6z6, Q8f6z6, Y8f6z6, G9f6z6, O9f6z6, W9f6z6, Eaf6z6, Maf6z6, Uaf6z6;
wire Cbf6z6, Kbf6z6, Sbf6z6, Acf6z6, Icf6z6, Qcf6z6, Ycf6z6, Gdf6z6, Odf6z6, Wdf6z6;
wire Eef6z6, Mef6z6, Uef6z6, Cff6z6, Kff6z6, Sff6z6, Agf6z6, Igf6z6, Qgf6z6, Ygf6z6;
wire Ghf6z6, Ohf6z6, Whf6z6, Eif6z6, Mif6z6, Uif6z6, Cjf6z6, Kjf6z6, Sjf6z6, Akf6z6;
wire Ikf6z6, Qkf6z6, Ykf6z6, Glf6z6, Olf6z6, Wlf6z6, Emf6z6, Mmf6z6, Umf6z6, Cnf6z6;
wire Knf6z6, Snf6z6, Aof6z6, Iof6z6, Qof6z6, Yof6z6, Gpf6z6, Opf6z6, Wpf6z6, Eqf6z6;
wire Mqf6z6, Uqf6z6, Crf6z6, Krf6z6, Srf6z6, Asf6z6, Isf6z6, Qsf6z6, Ysf6z6, Gtf6z6;
wire Otf6z6, Wtf6z6, Euf6z6, Muf6z6, Uuf6z6, Cvf6z6, Kvf6z6, Svf6z6, Awf6z6, Iwf6z6;
wire Qwf6z6, Ywf6z6, Gxf6z6, Oxf6z6, Wxf6z6, Eyf6z6, Myf6z6, Uyf6z6, Czf6z6, Kzf6z6;
wire Szf6z6, A0g6z6, I0g6z6, Q0g6z6, Y0g6z6, G1g6z6, O1g6z6, W1g6z6, E2g6z6, M2g6z6;
wire U2g6z6, C3g6z6, K3g6z6, S3g6z6, A4g6z6, I4g6z6, Q4g6z6, Y4g6z6, G5g6z6, O5g6z6;
wire W5g6z6, E6g6z6, M6g6z6, U6g6z6, C7g6z6, K7g6z6, S7g6z6, A8g6z6, I8g6z6, Q8g6z6;
wire Y8g6z6, G9g6z6, O9g6z6, W9g6z6, Eag6z6, Mag6z6, Uag6z6, Cbg6z6, Kbg6z6, Sbg6z6;
wire Acg6z6, Icg6z6, Qcg6z6, Ycg6z6, Gdg6z6, Odg6z6, Wdg6z6, Eeg6z6, Meg6z6, Ueg6z6;
wire Cfg6z6, Kfg6z6, Sfg6z6, Agg6z6, Igg6z6, Qgg6z6, Ygg6z6, Ghg6z6, Ohg6z6, Whg6z6;
wire Eig6z6, Mig6z6, Uig6z6, Cjg6z6, Kjg6z6, Sjg6z6, Akg6z6, Ikg6z6, Qkg6z6, Ykg6z6;
wire Glg6z6, Olg6z6, Wlg6z6, Emg6z6, Mmg6z6, Umg6z6, Cng6z6, Kng6z6, Sng6z6, Aog6z6;
wire Iog6z6, Qog6z6, Yog6z6, Gpg6z6, Opg6z6, Wpg6z6, Eqg6z6, Mqg6z6, Uqg6z6, Crg6z6;
wire Krg6z6, Srg6z6, Asg6z6, Isg6z6, Qsg6z6, Ysg6z6, Gtg6z6, Otg6z6, Wtg6z6, Eug6z6;
wire Mug6z6, Uug6z6, Cvg6z6, Kvg6z6, Svg6z6, Awg6z6, Iwg6z6, Qwg6z6, Ywg6z6, Gxg6z6;
wire Oxg6z6, Wxg6z6, Eyg6z6, Myg6z6, Uyg6z6, Czg6z6, Kzg6z6, Szg6z6, A0h6z6, I0h6z6;
wire Q0h6z6, Y0h6z6, G1h6z6, O1h6z6, W1h6z6, E2h6z6, M2h6z6, U2h6z6, C3h6z6, K3h6z6;
wire S3h6z6, A4h6z6, I4h6z6, Q4h6z6, Y4h6z6, G5h6z6, O5h6z6, W5h6z6, E6h6z6, M6h6z6;
wire U6h6z6, C7h6z6, K7h6z6, S7h6z6, A8h6z6, I8h6z6, Q8h6z6, Y8h6z6, G9h6z6, O9h6z6;
wire W9h6z6, Eah6z6, Mah6z6, Uah6z6, Cbh6z6, Kbh6z6, Sbh6z6, Ach6z6, Ich6z6, Qch6z6;
wire Ych6z6, Gdh6z6, Odh6z6, Wdh6z6, Eeh6z6, Meh6z6, Ueh6z6, Cfh6z6, Kfh6z6, Sfh6z6;
wire Agh6z6, Igh6z6, Qgh6z6, Ygh6z6, Ghh6z6, Ohh6z6, Whh6z6, Eih6z6, Mih6z6, Uih6z6;
wire Cjh6z6, Kjh6z6, Sjh6z6, Akh6z6, Ikh6z6, Qkh6z6, Ykh6z6, Glh6z6, Olh6z6, Wlh6z6;
wire Emh6z6, Mmh6z6, Umh6z6, Cnh6z6, Knh6z6, Snh6z6, Aoh6z6, Ioh6z6, Qoh6z6, Yoh6z6;
wire Gph6z6, Oph6z6, Wph6z6, Eqh6z6, Mqh6z6, Uqh6z6, Crh6z6, Krh6z6, Srh6z6, Ash6z6;
wire Ish6z6, Qsh6z6, Ysh6z6, Gth6z6, Oth6z6, Wth6z6, Euh6z6, Muh6z6, Uuh6z6, Cvh6z6;
wire Kvh6z6, Svh6z6, Awh6z6, Iwh6z6, Qwh6z6, Ywh6z6, Gxh6z6, Oxh6z6, Wxh6z6, Eyh6z6;
wire Myh6z6, Uyh6z6, Czh6z6, Kzh6z6, Szh6z6, A0i6z6, I0i6z6, Q0i6z6, Y0i6z6, G1i6z6;
wire O1i6z6, W1i6z6, E2i6z6, M2i6z6, U2i6z6, C3i6z6, K3i6z6, S3i6z6, A4i6z6, I4i6z6;
wire Q4i6z6, Y4i6z6, G5i6z6, O5i6z6, W5i6z6, E6i6z6, M6i6z6, U6i6z6, C7i6z6, K7i6z6;
wire S7i6z6, A8i6z6, I8i6z6, Q8i6z6, Y8i6z6, G9i6z6, O9i6z6, W9i6z6, Eai6z6, Mai6z6;
wire Uai6z6, Cbi6z6, Kbi6z6, Sbi6z6, Aci6z6, Ici6z6, Qci6z6, Yci6z6, Gdi6z6, Odi6z6;
wire Wdi6z6, Eei6z6, Mei6z6, Uei6z6, Cfi6z6, Kfi6z6, Sfi6z6, Agi6z6, Igi6z6, Qgi6z6;
wire Ygi6z6, Ghi6z6, Ohi6z6, Whi6z6, Eii6z6, Mii6z6, Uii6z6, Cji6z6, Kji6z6, Sji6z6;
wire Aki6z6, Iki6z6, Qki6z6, Yki6z6, Gli6z6, Oli6z6, Wli6z6, Emi6z6, Mmi6z6, Umi6z6;
wire Cni6z6, Kni6z6, Sni6z6, Aoi6z6, Ioi6z6, Qoi6z6, Yoi6z6, Gpi6z6, Opi6z6, Wpi6z6;
wire Eqi6z6, Mqi6z6, Uqi6z6, Cri6z6, Kri6z6, Sri6z6, Asi6z6, Isi6z6, Qsi6z6, Ysi6z6;
wire Gti6z6, Oti6z6, Wti6z6, Eui6z6, Mui6z6, Uui6z6, Cvi6z6, Kvi6z6, Svi6z6, Awi6z6;
wire Iwi6z6, Qwi6z6, Ywi6z6, Gxi6z6, Oxi6z6, Wxi6z6, Eyi6z6, Myi6z6, Uyi6z6, Czi6z6;
wire Kzi6z6, Szi6z6, A0j6z6, I0j6z6, Q0j6z6, Y0j6z6, G1j6z6, O1j6z6, W1j6z6, E2j6z6;
wire M2j6z6, U2j6z6, C3j6z6, K3j6z6, S3j6z6, A4j6z6, I4j6z6, Q4j6z6, Y4j6z6, G5j6z6;
wire O5j6z6, W5j6z6, E6j6z6, M6j6z6, U6j6z6, C7j6z6, K7j6z6, S7j6z6, A8j6z6, I8j6z6;
wire Q8j6z6, Y8j6z6, G9j6z6, O9j6z6, W9j6z6, Eaj6z6, Maj6z6, Uaj6z6, Cbj6z6, Kbj6z6;
wire Sbj6z6, Acj6z6, Icj6z6, Qcj6z6, Ycj6z6, Gdj6z6, Odj6z6, Wdj6z6, Eej6z6, Mej6z6;
wire Uej6z6, Cfj6z6, Kfj6z6, Sfj6z6, Agj6z6, Igj6z6, Qgj6z6, Ygj6z6, Ghj6z6, Ohj6z6;
wire Whj6z6, Eij6z6, Mij6z6, Uij6z6, Cjj6z6, Kjj6z6, Sjj6z6, Akj6z6, Ikj6z6, Qkj6z6;
wire Ykj6z6, Glj6z6, Olj6z6, Wlj6z6, Emj6z6, Mmj6z6, Umj6z6, Cnj6z6, Knj6z6, Snj6z6;
wire Aoj6z6, Ioj6z6, Qoj6z6, Yoj6z6, Gpj6z6, Opj6z6, Wpj6z6, Eqj6z6, Mqj6z6, Uqj6z6;
wire Crj6z6, Krj6z6, Srj6z6, Asj6z6, Isj6z6, Qsj6z6, Ysj6z6, Gtj6z6, Otj6z6, Wtj6z6;
wire Euj6z6, Muj6z6, Uuj6z6, Cvj6z6, Kvj6z6, Svj6z6, Awj6z6, Iwj6z6, Qwj6z6, Ywj6z6;
wire Gxj6z6, Oxj6z6, Wxj6z6, Eyj6z6, Myj6z6, Uyj6z6, Czj6z6, Kzj6z6, Szj6z6, A0k6z6;
wire I0k6z6, Q0k6z6, Y0k6z6, G1k6z6, O1k6z6, W1k6z6, E2k6z6, M2k6z6, U2k6z6, C3k6z6;
wire K3k6z6, S3k6z6, A4k6z6, I4k6z6, Q4k6z6, Y4k6z6, G5k6z6, O5k6z6, W5k6z6, E6k6z6;
wire M6k6z6, U6k6z6, C7k6z6, K7k6z6, S7k6z6, A8k6z6, I8k6z6, Q8k6z6, Y8k6z6, G9k6z6;
wire O9k6z6, W9k6z6, Eak6z6, Mak6z6, Uak6z6, Cbk6z6, Kbk6z6, Sbk6z6, Ack6z6, Ick6z6;
wire Qck6z6, Yck6z6, Gdk6z6, Odk6z6, Wdk6z6, Eek6z6, Mek6z6, Uek6z6, Cfk6z6, Kfk6z6;
wire Sfk6z6, Agk6z6, Igk6z6, Qgk6z6, Ygk6z6, Ghk6z6, Ohk6z6, Whk6z6, Eik6z6, Mik6z6;
wire Uik6z6, Cjk6z6, Kjk6z6, Sjk6z6, Akk6z6, Ikk6z6, Qkk6z6, Ykk6z6, Glk6z6, Olk6z6;
wire Wlk6z6, Emk6z6, Mmk6z6, Umk6z6, Cnk6z6, Knk6z6, Snk6z6, Aok6z6, Iok6z6, Qok6z6;
wire Yok6z6, Gpk6z6, Opk6z6, Wpk6z6, Eqk6z6, Mqk6z6, Uqk6z6, Crk6z6, Krk6z6, Srk6z6;
wire Ask6z6, Isk6z6, Qsk6z6, Ysk6z6, Gtk6z6, Otk6z6, Wtk6z6, Euk6z6, Muk6z6, Uuk6z6;
wire Cvk6z6, Kvk6z6, Svk6z6, Awk6z6, Iwk6z6, Qwk6z6, Ywk6z6, Gxk6z6, Oxk6z6, Wxk6z6;
wire Eyk6z6, Myk6z6, Uyk6z6, Czk6z6, Kzk6z6, Szk6z6, A0l6z6, I0l6z6, Q0l6z6, Y0l6z6;
wire G1l6z6, O1l6z6, W1l6z6, E2l6z6, M2l6z6, U2l6z6, C3l6z6, K3l6z6, S3l6z6, A4l6z6;
wire I4l6z6, Q4l6z6, Y4l6z6, G5l6z6, O5l6z6, W5l6z6, E6l6z6, M6l6z6, U6l6z6, C7l6z6;
wire K7l6z6, S7l6z6, A8l6z6, I8l6z6, Q8l6z6, Y8l6z6, G9l6z6, O9l6z6, W9l6z6, Eal6z6;
wire Mal6z6, Ual6z6, Cbl6z6, Kbl6z6, Sbl6z6, Acl6z6, Icl6z6, Qcl6z6, Ycl6z6, Gdl6z6;
wire Odl6z6, Wdl6z6, Eel6z6, Mel6z6, Uel6z6, Cfl6z6, Kfl6z6, Sfl6z6, Agl6z6, Igl6z6;
wire Qgl6z6, Ygl6z6, Ghl6z6, Ohl6z6, Whl6z6, Eil6z6, Mil6z6, Uil6z6, Cjl6z6, Kjl6z6;
wire Sjl6z6, Akl6z6, Ikl6z6, Qkl6z6, Ykl6z6, Gll6z6, Oll6z6, Wll6z6, Eml6z6, Mml6z6;
wire Uml6z6, Cnl6z6, Knl6z6, Snl6z6, Aol6z6, Iol6z6, Qol6z6, Yol6z6, Gpl6z6, Opl6z6;
wire Wpl6z6, Eql6z6, Mql6z6, Uql6z6, Crl6z6, Krl6z6, Srl6z6, Asl6z6, Isl6z6, Qsl6z6;
wire Ysl6z6, Gtl6z6, Otl6z6, Wtl6z6, Eul6z6, Mul6z6, Uul6z6, Cvl6z6, Kvl6z6, Svl6z6;
wire Awl6z6, Iwl6z6, Qwl6z6, Ywl6z6, Gxl6z6, Oxl6z6, Wxl6z6, Eyl6z6, Myl6z6, Uyl6z6;
wire Czl6z6, Kzl6z6, Szl6z6, A0m6z6, I0m6z6, Q0m6z6, Y0m6z6, G1m6z6, O1m6z6, W1m6z6;
wire E2m6z6, M2m6z6, U2m6z6, C3m6z6, K3m6z6, S3m6z6, A4m6z6, I4m6z6, Q4m6z6, Y4m6z6;
wire G5m6z6, O5m6z6, W5m6z6, E6m6z6, M6m6z6, U6m6z6, C7m6z6, K7m6z6, S7m6z6, A8m6z6;
wire I8m6z6, Q8m6z6, Y8m6z6, G9m6z6, O9m6z6, W9m6z6, Eam6z6, Mam6z6, Uam6z6, Cbm6z6;
wire Kbm6z6, Sbm6z6, Acm6z6, Icm6z6, Qcm6z6, Ycm6z6, Gdm6z6, Odm6z6, Wdm6z6, Eem6z6;
wire Mem6z6, Uem6z6, Cfm6z6, Kfm6z6, Sfm6z6, Agm6z6, Igm6z6, Qgm6z6, Ygm6z6, Ghm6z6;
wire Ohm6z6, Whm6z6, Eim6z6, Mim6z6, Uim6z6, Cjm6z6, Kjm6z6, Sjm6z6, Akm6z6, Ikm6z6;
wire Qkm6z6, Ykm6z6, Glm6z6, Olm6z6, Wlm6z6, Emm6z6, Mmm6z6, Umm6z6, Cnm6z6, Knm6z6;
wire Snm6z6, Aom6z6, Iom6z6, Qom6z6, Yom6z6, Gpm6z6, Opm6z6, Wpm6z6, Eqm6z6, Mqm6z6;
wire Uqm6z6, Crm6z6, Krm6z6, Srm6z6, Asm6z6, Ism6z6, Qsm6z6, Ysm6z6, Gtm6z6, Otm6z6;
wire Wtm6z6, Eum6z6, Mum6z6, Uum6z6, Cvm6z6, Kvm6z6, Svm6z6, Awm6z6, Iwm6z6, Qwm6z6;
wire Ywm6z6, Gxm6z6, Oxm6z6, Wxm6z6, Eym6z6, Mym6z6, Uym6z6, Czm6z6, Kzm6z6, Szm6z6;
wire A0n6z6, I0n6z6, Q0n6z6, Y0n6z6, G1n6z6, O1n6z6, W1n6z6, E2n6z6, M2n6z6, U2n6z6;
wire C3n6z6, K3n6z6, S3n6z6, A4n6z6, I4n6z6, Q4n6z6, Y4n6z6, G5n6z6, O5n6z6, W5n6z6;
wire E6n6z6, M6n6z6, U6n6z6, C7n6z6, K7n6z6, S7n6z6, A8n6z6, I8n6z6, Q8n6z6, Y8n6z6;
wire G9n6z6, O9n6z6, W9n6z6, Ean6z6, Man6z6, Uan6z6, Cbn6z6, Kbn6z6, Sbn6z6, Acn6z6;
wire Icn6z6, Qcn6z6, Ycn6z6, Gdn6z6, Odn6z6, Wdn6z6, Een6z6, Men6z6, Uen6z6, Cfn6z6;
wire Kfn6z6, Sfn6z6, Agn6z6, Ign6z6, Qgn6z6, Ygn6z6, Ghn6z6, Ohn6z6, Whn6z6, Ein6z6;
wire Min6z6, Uin6z6, Cjn6z6, Kjn6z6, Sjn6z6, Akn6z6, Ikn6z6, Qkn6z6, Ykn6z6, Gln6z6;
wire Oln6z6, Wln6z6, Emn6z6, Mmn6z6, Umn6z6, Cnn6z6, Knn6z6, Snn6z6, Aon6z6, Ion6z6;
wire Qon6z6, Yon6z6, Gpn6z6, Opn6z6, Wpn6z6, Eqn6z6, Mqn6z6, Uqn6z6, Crn6z6, Krn6z6;
wire Srn6z6, Asn6z6, Isn6z6, Qsn6z6, Ysn6z6, Gtn6z6, Otn6z6, Wtn6z6, Eun6z6, Mun6z6;
wire Uun6z6, Cvn6z6, Kvn6z6, Svn6z6, Awn6z6, Iwn6z6, Qwn6z6, Ywn6z6, Gxn6z6, Oxn6z6;
wire Wxn6z6, Eyn6z6, Myn6z6, Uyn6z6, Czn6z6, Kzn6z6, Szn6z6, A0o6z6, I0o6z6, Q0o6z6;
wire Y0o6z6, G1o6z6, O1o6z6, W1o6z6, E2o6z6, M2o6z6, U2o6z6, C3o6z6, K3o6z6, S3o6z6;
wire A4o6z6, I4o6z6, Q4o6z6, Y4o6z6, G5o6z6, O5o6z6, W5o6z6, E6o6z6, M6o6z6, U6o6z6;
wire C7o6z6, K7o6z6, S7o6z6, A8o6z6, I8o6z6, Q8o6z6, Y8o6z6, G9o6z6, O9o6z6, W9o6z6;
wire Eao6z6, Mao6z6, Uao6z6, Cbo6z6, Kbo6z6, Sbo6z6, Aco6z6, Ico6z6, Qco6z6, Yco6z6;
wire Gdo6z6, Odo6z6, Wdo6z6, Eeo6z6, Meo6z6, Ueo6z6, Cfo6z6, Kfo6z6, Sfo6z6, Ago6z6;
wire Igo6z6, Qgo6z6, Ygo6z6, Gho6z6, Oho6z6, Who6z6, Eio6z6, Mio6z6, Uio6z6, Cjo6z6;
wire Kjo6z6, Sjo6z6, Ako6z6, Iko6z6, Qko6z6, Yko6z6, Glo6z6, Olo6z6, Wlo6z6, Emo6z6;
wire Mmo6z6, Umo6z6, Cno6z6, Kno6z6, Sno6z6, Aoo6z6, Ioo6z6, Qoo6z6, Yoo6z6, Gpo6z6;
wire Opo6z6, Wpo6z6, Eqo6z6, Mqo6z6, Uqo6z6, Cro6z6, Kro6z6, Sro6z6, Aso6z6, Iso6z6;
wire Qso6z6, Yso6z6, Gto6z6, Oto6z6, Wto6z6, Euo6z6, Muo6z6, Uuo6z6, Cvo6z6, Kvo6z6;
wire Svo6z6, Awo6z6, Iwo6z6, Qwo6z6, Ywo6z6, Gxo6z6, Oxo6z6, Wxo6z6, Eyo6z6, Myo6z6;
wire Uyo6z6, Czo6z6, Kzo6z6, Szo6z6, A0p6z6, I0p6z6, Q0p6z6, Y0p6z6, G1p6z6, O1p6z6;
wire W1p6z6, E2p6z6, M2p6z6, U2p6z6, C3p6z6, K3p6z6, S3p6z6, A4p6z6, I4p6z6, Q4p6z6;
wire Y4p6z6, G5p6z6, O5p6z6, W5p6z6, E6p6z6, M6p6z6, U6p6z6, C7p6z6, K7p6z6, S7p6z6;
wire A8p6z6, I8p6z6, Q8p6z6, Y8p6z6, G9p6z6, O9p6z6, W9p6z6, Eap6z6, Map6z6, Uap6z6;
wire Cbp6z6, Kbp6z6, Sbp6z6, Acp6z6, Icp6z6, Qcp6z6, Ycp6z6, Gdp6z6, Odp6z6, Wdp6z6;
wire Eep6z6, Mep6z6, Uep6z6, Cfp6z6, Kfp6z6, Sfp6z6, Agp6z6, Igp6z6, Qgp6z6, Ygp6z6;
wire Ghp6z6, Ohp6z6, Whp6z6, Eip6z6, Mip6z6, Uip6z6, Cjp6z6, Kjp6z6, Sjp6z6, Akp6z6;
wire Ikp6z6, Qkp6z6, Ykp6z6, Glp6z6, Olp6z6, Wlp6z6, Emp6z6, Mmp6z6, Ump6z6, Cnp6z6;
wire Knp6z6, Snp6z6, Aop6z6, Iop6z6, Qop6z6, Yop6z6, Gpp6z6, Opp6z6, Wpp6z6, Eqp6z6;
wire Mqp6z6, Uqp6z6, Crp6z6, Krp6z6, Srp6z6, Asp6z6, Isp6z6, Qsp6z6, Ysp6z6, Gtp6z6;
wire Otp6z6, Wtp6z6, Eup6z6, Mup6z6, Uup6z6, Cvp6z6, Kvp6z6, Svp6z6, Awp6z6, Iwp6z6;
wire Qwp6z6, Ywp6z6, Gxp6z6, Oxp6z6, Wxp6z6, Eyp6z6, Myp6z6, Uyp6z6, Czp6z6, Kzp6z6;
wire Szp6z6, A0q6z6, I0q6z6, Q0q6z6, Y0q6z6, G1q6z6, O1q6z6, W1q6z6, E2q6z6, M2q6z6;
wire U2q6z6, C3q6z6, K3q6z6, S3q6z6, A4q6z6, I4q6z6, Q4q6z6, Y4q6z6, G5q6z6, O5q6z6;
wire W5q6z6, E6q6z6, M6q6z6, U6q6z6, C7q6z6, K7q6z6, S7q6z6, A8q6z6, I8q6z6, Q8q6z6;
wire Y8q6z6, G9q6z6, O9q6z6, W9q6z6, Eaq6z6, Maq6z6, Uaq6z6, Cbq6z6, Kbq6z6, Sbq6z6;
wire Acq6z6, Icq6z6, Qcq6z6, Ycq6z6, Gdq6z6, Odq6z6, Wdq6z6, Eeq6z6, Meq6z6, Ueq6z6;
wire Cfq6z6, Kfq6z6, Sfq6z6, Agq6z6, Igq6z6, Qgq6z6, Ygq6z6, Ghq6z6, Ohq6z6, Whq6z6;
wire Eiq6z6, Miq6z6, Uiq6z6, Cjq6z6, Kjq6z6, Sjq6z6, Akq6z6, Ikq6z6, Qkq6z6, Ykq6z6;
wire Glq6z6, Olq6z6, Wlq6z6, Emq6z6, Mmq6z6, Umq6z6, Cnq6z6, Knq6z6, Snq6z6, Aoq6z6;
wire Ioq6z6, Qoq6z6, Yoq6z6, Gpq6z6, Opq6z6, Wpq6z6, Eqq6z6, Mqq6z6, Uqq6z6, Crq6z6;
wire Krq6z6, Srq6z6, Asq6z6, Isq6z6, Qsq6z6, Ysq6z6, Gtq6z6, Otq6z6, Wtq6z6, Euq6z6;
wire Muq6z6, Uuq6z6, Cvq6z6, Kvq6z6, Svq6z6, Awq6z6, Iwq6z6, Qwq6z6, Ywq6z6, Gxq6z6;
wire Oxq6z6, Wxq6z6, Eyq6z6, Myq6z6, Uyq6z6, Czq6z6, Kzq6z6, Szq6z6, A0r6z6, I0r6z6;
wire Q0r6z6, Y0r6z6, G1r6z6, O1r6z6, W1r6z6, E2r6z6, M2r6z6, U2r6z6, C3r6z6, K3r6z6;
wire S3r6z6, A4r6z6, I4r6z6, Q4r6z6, Y4r6z6, G5r6z6, O5r6z6, W5r6z6, E6r6z6, M6r6z6;
wire U6r6z6, C7r6z6, K7r6z6, S7r6z6, A8r6z6, I8r6z6, Q8r6z6, Y8r6z6, G9r6z6, O9r6z6;
wire W9r6z6, Ear6z6, Mar6z6, Uar6z6, Cbr6z6, Kbr6z6, Sbr6z6, Acr6z6, Icr6z6, Qcr6z6;
wire Ycr6z6, Gdr6z6, Odr6z6, Wdr6z6, Eer6z6, Mer6z6, Uer6z6, Cfr6z6, Kfr6z6, Sfr6z6;
wire Agr6z6, Igr6z6, Qgr6z6, Ygr6z6, Ghr6z6, Ohr6z6, Whr6z6, Eir6z6, Mir6z6, Uir6z6;
wire Cjr6z6, Kjr6z6, Sjr6z6, Akr6z6, Ikr6z6, Qkr6z6, Ykr6z6, Glr6z6, Olr6z6, Wlr6z6;
wire Emr6z6, Mmr6z6, Umr6z6, Cnr6z6, Knr6z6, Snr6z6, Aor6z6, Ior6z6, Qor6z6, Yor6z6;
wire Gpr6z6, Opr6z6, Wpr6z6, Eqr6z6, Mqr6z6, Uqr6z6, Crr6z6, Krr6z6, Srr6z6, Asr6z6;
wire Isr6z6, Qsr6z6, Ysr6z6, Gtr6z6, Otr6z6, Wtr6z6, Eur6z6, Mur6z6, Uur6z6, Cvr6z6;
wire Kvr6z6, Svr6z6, Awr6z6, Iwr6z6, Qwr6z6, Ywr6z6, Gxr6z6, Oxr6z6, Wxr6z6, Eyr6z6;
wire Myr6z6, Uyr6z6, Czr6z6, Kzr6z6, Szr6z6, A0s6z6, I0s6z6, Q0s6z6, Y0s6z6, G1s6z6;
wire O1s6z6, W1s6z6, E2s6z6, M2s6z6, U2s6z6, C3s6z6, K3s6z6, S3s6z6, A4s6z6, I4s6z6;
wire Q4s6z6, Y4s6z6, G5s6z6, O5s6z6, W5s6z6, E6s6z6, M6s6z6, U6s6z6, C7s6z6, K7s6z6;
wire S7s6z6, A8s6z6, I8s6z6, Q8s6z6, Y8s6z6, G9s6z6, O9s6z6, W9s6z6, Eas6z6, Mas6z6;
wire Uas6z6, Cbs6z6, Kbs6z6, Sbs6z6, Acs6z6, Ics6z6, Qcs6z6, Ycs6z6, Gds6z6, Ods6z6;
wire Wds6z6, Ees6z6, Mes6z6, Ues6z6, Cfs6z6, Kfs6z6, Sfs6z6, Ags6z6, Igs6z6, Qgs6z6;
wire Ygs6z6, Ghs6z6, Ohs6z6, Whs6z6, Eis6z6, Mis6z6, Uis6z6, Cjs6z6, Kjs6z6, Sjs6z6;
wire Aks6z6, Iks6z6, Qks6z6, Yks6z6, Gls6z6, Ols6z6, Wls6z6, Ems6z6, Mms6z6, Ums6z6;
wire Cns6z6, Kns6z6, Sns6z6, Aos6z6, Ios6z6, Qos6z6, Yos6z6, Gps6z6, Ops6z6, Wps6z6;
wire Eqs6z6, Mqs6z6, Uqs6z6, Crs6z6, Krs6z6, Srs6z6, Ass6z6, Iss6z6, Qss6z6, Yss6z6;
wire Gts6z6, Ots6z6, Wts6z6, Eus6z6, Mus6z6, Uus6z6, Cvs6z6, Kvs6z6, Svs6z6, Aws6z6;
wire Iws6z6, Qws6z6, Yws6z6, Gxs6z6, Oxs6z6, Wxs6z6, Eys6z6, Mys6z6, Uys6z6, Czs6z6;
wire Kzs6z6, Szs6z6, A0t6z6, I0t6z6, Q0t6z6, Y0t6z6, G1t6z6, O1t6z6, W1t6z6, E2t6z6;
wire M2t6z6, U2t6z6, C3t6z6, K3t6z6, S3t6z6, A4t6z6, I4t6z6, Q4t6z6, Y4t6z6, G5t6z6;
wire O5t6z6, W5t6z6, E6t6z6, M6t6z6, U6t6z6, C7t6z6, K7t6z6, S7t6z6, A8t6z6, I8t6z6;
wire Q8t6z6, Y8t6z6, G9t6z6, O9t6z6, W9t6z6, Eat6z6, Mat6z6, Uat6z6, Cbt6z6, Kbt6z6;
wire Sbt6z6, Act6z6, Ict6z6, Qct6z6, Yct6z6, Gdt6z6, Odt6z6, Wdt6z6, Eet6z6, Met6z6;
wire Uet6z6, Cft6z6, Kft6z6, Sft6z6, Agt6z6, Igt6z6, Qgt6z6, Ygt6z6, Ght6z6, Oht6z6;
wire Wht6z6, Eit6z6, Mit6z6, Uit6z6, Cjt6z6, Kjt6z6, Sjt6z6, Akt6z6, Ikt6z6, Qkt6z6;
wire Ykt6z6, Glt6z6, Olt6z6, Wlt6z6, Emt6z6, Mmt6z6, Umt6z6, Cnt6z6, Knt6z6, Snt6z6;
wire Aot6z6, Iot6z6, Qot6z6, Yot6z6, Gpt6z6, Opt6z6, Wpt6z6, Eqt6z6, Mqt6z6, Uqt6z6;
wire Crt6z6, Krt6z6, Srt6z6, Ast6z6, Ist6z6, Qst6z6, Yst6z6, Gtt6z6, Ott6z6, Wtt6z6;
wire Eut6z6, Mut6z6, Uut6z6, Cvt6z6, Kvt6z6, Svt6z6, Awt6z6, Iwt6z6, Qwt6z6, Ywt6z6;
wire Gxt6z6, Oxt6z6, Wxt6z6, Eyt6z6, Myt6z6, Uyt6z6, Czt6z6, Kzt6z6, Szt6z6, A0u6z6;
wire I0u6z6, Q0u6z6, Y0u6z6, G1u6z6, O1u6z6, W1u6z6, E2u6z6, M2u6z6, U2u6z6, C3u6z6;
wire K3u6z6, S3u6z6, A4u6z6, I4u6z6, Q4u6z6, Y4u6z6, G5u6z6, O5u6z6, W5u6z6, E6u6z6;
wire M6u6z6, U6u6z6, C7u6z6, K7u6z6, S7u6z6, A8u6z6, I8u6z6, Q8u6z6, Y8u6z6, G9u6z6;
wire O9u6z6, W9u6z6, Eau6z6, Mau6z6, Uau6z6, Cbu6z6, Kbu6z6, Sbu6z6, Acu6z6, Icu6z6;
wire Qcu6z6, Ycu6z6, Gdu6z6, Odu6z6, Wdu6z6, Eeu6z6, Meu6z6, Ueu6z6, Cfu6z6, Kfu6z6;
wire Sfu6z6, Agu6z6, Igu6z6, Qgu6z6, Ygu6z6, Ghu6z6, Ohu6z6, Whu6z6, Eiu6z6, Miu6z6;
wire Uiu6z6, Cju6z6, Kju6z6, Sju6z6, Aku6z6, Iku6z6, Qku6z6, Yku6z6, Glu6z6, Olu6z6;
wire Wlu6z6, Emu6z6, Mmu6z6, Umu6z6, Cnu6z6, Knu6z6, Snu6z6, Aou6z6, Iou6z6, Qou6z6;
wire You6z6, Gpu6z6, Opu6z6, Wpu6z6, Equ6z6, Mqu6z6, Uqu6z6, Cru6z6, Kru6z6, Sru6z6;
wire Asu6z6, Isu6z6, Qsu6z6, Ysu6z6, Gtu6z6, Otu6z6, Wtu6z6, Euu6z6, Muu6z6, Uuu6z6;
wire Cvu6z6, Kvu6z6, Svu6z6, Awu6z6, Iwu6z6, Qwu6z6, Ywu6z6, Gxu6z6, Oxu6z6, Wxu6z6;
wire Eyu6z6, Myu6z6, Uyu6z6, Czu6z6, Kzu6z6, Szu6z6, A0v6z6, I0v6z6, Q0v6z6, Y0v6z6;
wire G1v6z6, O1v6z6, W1v6z6, E2v6z6, M2v6z6, U2v6z6, C3v6z6, K3v6z6, S3v6z6, A4v6z6;
wire I4v6z6, Q4v6z6, Y4v6z6, G5v6z6, O5v6z6, W5v6z6, E6v6z6, M6v6z6, U6v6z6, C7v6z6;
wire K7v6z6, S7v6z6, A8v6z6, I8v6z6, Q8v6z6, Y8v6z6, G9v6z6, O9v6z6, W9v6z6, Eav6z6;
wire Mav6z6, Uav6z6, Cbv6z6, Kbv6z6, Sbv6z6, Acv6z6, Icv6z6, Qcv6z6, Ycv6z6, Gdv6z6;
wire Odv6z6, Wdv6z6, Eev6z6, Mev6z6, Uev6z6, Cfv6z6, Kfv6z6, Sfv6z6, Agv6z6, Igv6z6;
wire Qgv6z6, Ygv6z6, Ghv6z6, Ohv6z6, Whv6z6, Eiv6z6, Miv6z6, Uiv6z6, Cjv6z6, Kjv6z6;
wire Sjv6z6, Akv6z6, Ikv6z6, Qkv6z6, Ykv6z6, Glv6z6, Olv6z6, Wlv6z6, Emv6z6, Mmv6z6;
wire Umv6z6, Cnv6z6, Knv6z6, Snv6z6, Aov6z6, Iov6z6, Qov6z6, Yov6z6, Gpv6z6, Opv6z6;
wire Wpv6z6, Eqv6z6, Mqv6z6, Uqv6z6, Crv6z6, Krv6z6, Srv6z6, Asv6z6, Isv6z6, Qsv6z6;
wire Ysv6z6, Gtv6z6, Otv6z6, Wtv6z6, Euv6z6, Muv6z6, Uuv6z6, Cvv6z6, Kvv6z6, Svv6z6;
wire Awv6z6, Iwv6z6, Qwv6z6, Ywv6z6, Gxv6z6, Oxv6z6, Wxv6z6, Eyv6z6, Myv6z6, Uyv6z6;
wire Czv6z6, Kzv6z6, Szv6z6, A0w6z6, I0w6z6, Q0w6z6, Y0w6z6, G1w6z6, O1w6z6, W1w6z6;
wire E2w6z6, M2w6z6, U2w6z6, C3w6z6, K3w6z6, S3w6z6, A4w6z6, I4w6z6, Q4w6z6, Y4w6z6;
wire G5w6z6, O5w6z6, W5w6z6, E6w6z6, M6w6z6, U6w6z6, C7w6z6, K7w6z6, S7w6z6, A8w6z6;
wire I8w6z6, Q8w6z6, Y8w6z6, G9w6z6, O9w6z6, W9w6z6, Eaw6z6, Maw6z6, Uaw6z6, Cbw6z6;
wire Kbw6z6, Sbw6z6, Acw6z6, Icw6z6, Qcw6z6, Ycw6z6, Gdw6z6, Odw6z6, Wdw6z6, Eew6z6;
wire Mew6z6, Uew6z6, Cfw6z6, Kfw6z6, Sfw6z6, Agw6z6, Igw6z6, Qgw6z6, Ygw6z6, Ghw6z6;
wire Ohw6z6, Whw6z6, Eiw6z6, Miw6z6, Uiw6z6, Cjw6z6, Kjw6z6, Sjw6z6, Akw6z6, Ikw6z6;
wire Qkw6z6, Ykw6z6, Glw6z6, Olw6z6, Wlw6z6, Emw6z6, Mmw6z6, Umw6z6, Cnw6z6, Knw6z6;
wire Snw6z6, Aow6z6, Iow6z6, Qow6z6, Yow6z6, Gpw6z6, Opw6z6, Wpw6z6, Eqw6z6, Mqw6z6;
wire Uqw6z6, Crw6z6, Krw6z6, Srw6z6, Asw6z6, Isw6z6, Qsw6z6, Ysw6z6, Gtw6z6, Otw6z6;
wire Wtw6z6, Euw6z6, Muw6z6, Uuw6z6, Cvw6z6, Kvw6z6, Svw6z6, Aww6z6, Iww6z6, Qww6z6;
wire Yww6z6, Gxw6z6, Oxw6z6, Wxw6z6, Eyw6z6, Myw6z6, Uyw6z6, Czw6z6, Kzw6z6, Szw6z6;
wire A0x6z6, I0x6z6, Q0x6z6, Y0x6z6, G1x6z6, O1x6z6, W1x6z6, E2x6z6, M2x6z6, U2x6z6;
wire C3x6z6, K3x6z6, S3x6z6, A4x6z6, I4x6z6, Q4x6z6, Y4x6z6, G5x6z6, O5x6z6, W5x6z6;
wire E6x6z6, M6x6z6, U6x6z6, C7x6z6, K7x6z6, S7x6z6, A8x6z6, I8x6z6, Q8x6z6, Y8x6z6;
wire G9x6z6, O9x6z6, W9x6z6, Eax6z6, Max6z6, Uax6z6, Cbx6z6, Kbx6z6, Sbx6z6, Acx6z6;
wire Icx6z6, Qcx6z6, Ycx6z6, Gdx6z6, Odx6z6, Wdx6z6, Eex6z6, Mex6z6, Uex6z6, Cfx6z6;
wire Kfx6z6, Sfx6z6, Agx6z6, Igx6z6, Qgx6z6, Ygx6z6, Ghx6z6, Ohx6z6, Whx6z6, Eix6z6;
wire Mix6z6, Uix6z6, Cjx6z6, Kjx6z6, Sjx6z6, Akx6z6, Ikx6z6, Qkx6z6, Ykx6z6, Glx6z6;
wire Olx6z6, Wlx6z6, Emx6z6, Mmx6z6, Umx6z6, Cnx6z6, Knx6z6, Snx6z6, Aox6z6, Iox6z6;
wire Qox6z6, Yox6z6, Gpx6z6, Opx6z6, Wpx6z6, Eqx6z6, Mqx6z6, Uqx6z6, Crx6z6, Krx6z6;
wire Srx6z6, Asx6z6, Isx6z6, Qsx6z6, Ysx6z6, Gtx6z6, Otx6z6, Wtx6z6, Eux6z6, Mux6z6;
wire Uux6z6, Cvx6z6, Kvx6z6, Svx6z6, Awx6z6, Iwx6z6, Qwx6z6, Ywx6z6, Gxx6z6, Oxx6z6;
wire Wxx6z6, Eyx6z6, Myx6z6, Uyx6z6, Czx6z6, Kzx6z6, Szx6z6, A0y6z6, I0y6z6, Q0y6z6;
wire Y0y6z6, G1y6z6, O1y6z6, W1y6z6, E2y6z6, M2y6z6, U2y6z6, C3y6z6, K3y6z6, S3y6z6;
wire A4y6z6, I4y6z6, Q4y6z6, Y4y6z6, G5y6z6, O5y6z6, W5y6z6, E6y6z6, M6y6z6, U6y6z6;
wire C7y6z6, K7y6z6, S7y6z6, A8y6z6, I8y6z6, Q8y6z6, Y8y6z6, G9y6z6, O9y6z6, W9y6z6;
wire Eay6z6, May6z6, Uay6z6, Cby6z6, Kby6z6, Sby6z6, Acy6z6, Icy6z6, Qcy6z6, Ycy6z6;
wire Gdy6z6, Ody6z6, Wdy6z6, Eey6z6, Mey6z6, Uey6z6, Cfy6z6, Kfy6z6, Sfy6z6, Agy6z6;
wire Igy6z6, Qgy6z6, Ygy6z6, Ghy6z6, Ohy6z6, Why6z6, Eiy6z6, Miy6z6, Uiy6z6, Cjy6z6;
wire Kjy6z6, Sjy6z6, Aky6z6, Iky6z6, Qky6z6, Yky6z6, Gly6z6, Oly6z6, Wly6z6, Emy6z6;
wire Mmy6z6, Umy6z6, Cny6z6, Kny6z6, Sny6z6, Aoy6z6, Ioy6z6, Qoy6z6, Yoy6z6, Gpy6z6;
wire Opy6z6, Wpy6z6, Eqy6z6, Mqy6z6, Uqy6z6, Cry6z6, Kry6z6, Sry6z6, Asy6z6, Isy6z6;
wire Qsy6z6, Ysy6z6, Gty6z6, Oty6z6, Wty6z6, Euy6z6, Muy6z6, Uuy6z6, Cvy6z6, Kvy6z6;
wire Svy6z6, Awy6z6, Iwy6z6, Qwy6z6, Ywy6z6, Gxy6z6, Oxy6z6, Wxy6z6, Eyy6z6, Myy6z6;
wire Uyy6z6, Czy6z6, Kzy6z6, Szy6z6, A0z6z6, I0z6z6, Q0z6z6, Y0z6z6, G1z6z6, O1z6z6;
wire W1z6z6, E2z6z6, M2z6z6, U2z6z6, C3z6z6, K3z6z6, S3z6z6, A4z6z6, I4z6z6, Q4z6z6;
wire Y4z6z6, G5z6z6, O5z6z6, W5z6z6, E6z6z6, M6z6z6, U6z6z6, C7z6z6, K7z6z6, S7z6z6;
wire A8z6z6, I8z6z6, Q8z6z6, Y8z6z6, G9z6z6, O9z6z6, W9z6z6, Eaz6z6, Maz6z6, Uaz6z6;
wire Cbz6z6, Kbz6z6, Sbz6z6, Acz6z6, Icz6z6, Qcz6z6, Ycz6z6, Gdz6z6, Odz6z6, Wdz6z6;
wire Eez6z6, Mez6z6, Uez6z6, Cfz6z6, Kfz6z6, Sfz6z6, Agz6z6, Igz6z6, Qgz6z6, Ygz6z6;
wire Ghz6z6, Ohz6z6, Whz6z6, Eiz6z6, Miz6z6, Uiz6z6, Cjz6z6, Kjz6z6, Sjz6z6, Akz6z6;
wire Ikz6z6, Qkz6z6, Ykz6z6, Glz6z6, Olz6z6, Wlz6z6, Emz6z6, Mmz6z6, Umz6z6, Cnz6z6;
wire Knz6z6, Snz6z6, Aoz6z6, Ioz6z6, Qoz6z6, Yoz6z6, Gpz6z6, Opz6z6, Wpz6z6, Eqz6z6;
wire Mqz6z6, Uqz6z6, Crz6z6, Krz6z6, Srz6z6, Asz6z6, Isz6z6, Qsz6z6, Ysz6z6, Gtz6z6;
wire Otz6z6, Wtz6z6, Euz6z6, Muz6z6, Uuz6z6, Cvz6z6, Kvz6z6, Svz6z6, Awz6z6, Iwz6z6;
wire Qwz6z6, Ywz6z6, Gxz6z6, Oxz6z6, Wxz6z6, Eyz6z6, Myz6z6, Uyz6z6, Czz6z6, Kzz6z6;
wire Szz6z6, A007z6, I007z6, Q007z6, Y007z6, G107z6, O107z6, W107z6, E207z6, M207z6;
wire U207z6, C307z6, K307z6, S307z6, A407z6, I407z6, Q407z6, Y407z6, G507z6, O507z6;
wire W507z6, E607z6, M607z6, U607z6, C707z6, K707z6, S707z6, A807z6, I807z6, Q807z6;
wire Y807z6, G907z6, O907z6, W907z6, Ea07z6, Ma07z6, Ua07z6, Cb07z6, Kb07z6, Sb07z6;
wire Ac07z6, Ic07z6, Qc07z6, Yc07z6, Gd07z6, Od07z6, Wd07z6, Ee07z6, Me07z6, Ue07z6;
wire Cf07z6, Kf07z6, Sf07z6, Ag07z6, Ig07z6, Qg07z6, Yg07z6, Gh07z6, Oh07z6, Wh07z6;
wire Ei07z6, Mi07z6, Ui07z6, Cj07z6, Kj07z6, Sj07z6, Ak07z6, Ik07z6, Qk07z6, Yk07z6;
wire Gl07z6, Ol07z6, Wl07z6, Em07z6, Mm07z6, Um07z6, Cn07z6, Kn07z6, Sn07z6, Ao07z6;
wire Io07z6, Qo07z6, Yo07z6, Gp07z6, Op07z6, Wp07z6, Eq07z6, Mq07z6, Uq07z6, Cr07z6;
wire Kr07z6, Sr07z6, As07z6, Is07z6, Qs07z6, Ys07z6, Gt07z6, Ot07z6, Wt07z6, Eu07z6;
wire Mu07z6, Uu07z6, Cv07z6, Kv07z6, Sv07z6, Aw07z6, Iw07z6, Qw07z6, Yw07z6, Gx07z6;
wire Ox07z6, Wx07z6, Ey07z6, My07z6, Uy07z6, Cz07z6, Kz07z6, Sz07z6, A017z6, I017z6;
wire Q017z6, Y017z6, G117z6, O117z6, W117z6, E217z6, M217z6, U217z6, C317z6, K317z6;
wire S317z6, A417z6, I417z6, Q417z6, Y417z6, G517z6, O517z6, W517z6, E617z6, M617z6;
wire U617z6, C717z6, K717z6, S717z6, A817z6, I817z6, Q817z6, Y817z6, G917z6, O917z6;
wire W917z6, Ea17z6, Ma17z6, Ua17z6, Cb17z6, Kb17z6, Sb17z6, Ac17z6, Ic17z6, Qc17z6;
wire Yc17z6, Gd17z6, Od17z6, Wd17z6, Ee17z6, Me17z6, Ue17z6, Cf17z6, Kf17z6, Sf17z6;
wire Ag17z6, Ig17z6, Qg17z6, Yg17z6, Gh17z6, Oh17z6, Wh17z6, Ei17z6, Mi17z6, Ui17z6;
wire Cj17z6, Kj17z6, Sj17z6, Ak17z6, Ik17z6, Qk17z6, Yk17z6, Gl17z6, Ol17z6, Wl17z6;
wire Em17z6, Mm17z6, Um17z6, Cn17z6, Kn17z6, Sn17z6, Ao17z6, Io17z6, Qo17z6, Yo17z6;
wire Gp17z6, Op17z6, Wp17z6, Eq17z6, Mq17z6, Uq17z6, Cr17z6, Kr17z6, Sr17z6, As17z6;
wire Is17z6, Qs17z6, Ys17z6, Gt17z6, Ot17z6, Wt17z6, Eu17z6, Mu17z6, Uu17z6, Cv17z6;
wire Kv17z6, Sv17z6, Aw17z6, Iw17z6, Qw17z6, Yw17z6, Gx17z6, Ox17z6, Wx17z6, Ey17z6;
wire My17z6, Uy17z6, Cz17z6, Kz17z6, Sz17z6, A027z6, I027z6, Q027z6, Y027z6, G127z6;
wire O127z6, W127z6, E227z6, M227z6, U227z6, C327z6, K327z6, S327z6, A427z6, I427z6;
wire Q427z6, Y427z6, G527z6, O527z6, W527z6, E627z6, M627z6, U627z6, C727z6, K727z6;
wire S727z6, A827z6, I827z6, Q827z6, Y827z6, G927z6, O927z6, W927z6, Ea27z6, Ma27z6;
wire Ua27z6, Cb27z6, Kb27z6, Sb27z6, Ac27z6, Ic27z6, Qc27z6, Yc27z6, Gd27z6, Od27z6;
wire Wd27z6, Ee27z6, Me27z6, Ue27z6, Cf27z6, Kf27z6, Sf27z6, Ag27z6, Ig27z6, Qg27z6;
wire Yg27z6, Gh27z6, Oh27z6, Wh27z6, Ei27z6, Mi27z6, Ui27z6, Cj27z6, Kj27z6, Sj27z6;
wire Ak27z6, Ik27z6, Qk27z6, Yk27z6, Gl27z6, Ol27z6, Wl27z6, Em27z6, Mm27z6, Um27z6;
wire Cn27z6, Kn27z6, Sn27z6, Ao27z6, Io27z6, Qo27z6, Yo27z6, Gp27z6, Op27z6, Wp27z6;
wire Eq27z6, Mq27z6, Uq27z6, Cr27z6, Kr27z6, Sr27z6, As27z6, Is27z6, Qs27z6, Ys27z6;
wire Gt27z6, Ot27z6, Wt27z6, Eu27z6, Mu27z6, Uu27z6, Cv27z6, Kv27z6, Sv27z6, Aw27z6;
wire Iw27z6, Qw27z6, Yw27z6, Gx27z6, Ox27z6, Wx27z6, Ey27z6, My27z6, Uy27z6, Cz27z6;
wire Kz27z6, Sz27z6, A037z6, I037z6, Q037z6, Y037z6, G137z6, O137z6, W137z6, E237z6;
wire M237z6, U237z6, C337z6, K337z6, S337z6, A437z6, I437z6, Q437z6, Y437z6, G537z6;
wire O537z6, W537z6, E637z6, M637z6, U637z6, C737z6, K737z6, S737z6, A837z6, I837z6;
wire Q837z6, Y837z6, G937z6, O937z6, W937z6, Ea37z6, Ma37z6, Ua37z6, Cb37z6, Kb37z6;
wire Sb37z6, Ac37z6, Ic37z6, Qc37z6, Yc37z6, Gd37z6, Od37z6, Wd37z6, Ee37z6, Me37z6;
wire Ue37z6, Cf37z6, Kf37z6, Sf37z6, Ag37z6, Ig37z6, Qg37z6, Yg37z6, Gh37z6, Oh37z6;
wire Wh37z6, Ei37z6, Mi37z6, Ui37z6, Cj37z6, Kj37z6, Sj37z6, Ak37z6, Ik37z6, Qk37z6;
wire Yk37z6, Gl37z6, Ol37z6, Wl37z6, Em37z6, Mm37z6, Um37z6, Cn37z6, Kn37z6, Sn37z6;
wire Ao37z6, Io37z6, Qo37z6, Yo37z6, Gp37z6, Op37z6, Wp37z6, Eq37z6, Mq37z6, Uq37z6;
wire Cr37z6, Kr37z6, Sr37z6, As37z6, Is37z6, Qs37z6, Ys37z6, Gt37z6, Ot37z6, Wt37z6;
wire Eu37z6, Mu37z6, Uu37z6, Cv37z6, Kv37z6, Sv37z6, Aw37z6, Iw37z6, Qw37z6, Yw37z6;
wire Gx37z6, Ox37z6, Wx37z6, Ey37z6, My37z6, Uy37z6, Cz37z6, Kz37z6, Sz37z6, A047z6;
wire I047z6, Q047z6, Y047z6, G147z6, O147z6, W147z6, E247z6, M247z6, U247z6, C347z6;
wire K347z6, S347z6, A447z6, I447z6, Q447z6, Y447z6, G547z6, O547z6, W547z6, E647z6;
wire M647z6, U647z6, C747z6, K747z6, S747z6, A847z6, I847z6, Q847z6, Y847z6, G947z6;
wire O947z6, W947z6, Ea47z6, Ma47z6, Ua47z6, Cb47z6, Kb47z6, Sb47z6, Ac47z6, Ic47z6;
wire Qc47z6, Yc47z6, Gd47z6, Od47z6, Wd47z6, Ee47z6, Me47z6, Ue47z6, Cf47z6, Kf47z6;
wire Sf47z6, Ag47z6, Ig47z6, Qg47z6, Yg47z6, Gh47z6, Oh47z6, Wh47z6, Ei47z6, Mi47z6;
wire Ui47z6, Cj47z6, Kj47z6, Sj47z6, Ak47z6, Ik47z6, Qk47z6, Yk47z6, Gl47z6, Ol47z6;
wire Wl47z6, Em47z6, Mm47z6, Um47z6, Cn47z6, Kn47z6, Sn47z6, Ao47z6, Io47z6, Qo47z6;
wire Yo47z6, Gp47z6, Op47z6, Wp47z6, Eq47z6, Mq47z6, Uq47z6, Cr47z6, Kr47z6, Sr47z6;
wire As47z6, Is47z6, Qs47z6, Ys47z6, Gt47z6, Ot47z6, Wt47z6, Eu47z6, Mu47z6, Uu47z6;
wire Cv47z6, Kv47z6, Sv47z6, Aw47z6, Iw47z6, Qw47z6, Yw47z6, Gx47z6, Ox47z6, Wx47z6;
wire Ey47z6, My47z6, Uy47z6, Cz47z6, Kz47z6, Sz47z6, A057z6, I057z6, Q057z6, Y057z6;
wire G157z6, O157z6, W157z6, E257z6, M257z6, U257z6, C357z6, K357z6, S357z6, A457z6;
wire I457z6, Q457z6, Y457z6, G557z6, O557z6, W557z6, E657z6, M657z6, U657z6, C757z6;
wire K757z6, S757z6, A857z6, I857z6, Q857z6, Y857z6, G957z6, O957z6, W957z6, Ea57z6;
wire Ma57z6, Ua57z6, Cb57z6, Kb57z6, Sb57z6, Ac57z6, Ic57z6, Qc57z6, Yc57z6, Gd57z6;
wire Od57z6, Wd57z6, Ee57z6, Me57z6, Ue57z6, Cf57z6, Kf57z6, Sf57z6, Ag57z6, Ig57z6;
wire Qg57z6, Yg57z6, Gh57z6, Oh57z6, Wh57z6, Ei57z6, Mi57z6, Ui57z6, Cj57z6, Kj57z6;
wire Sj57z6, Ak57z6, Ik57z6, Qk57z6, Yk57z6, Gl57z6, Ol57z6, Wl57z6, Em57z6, Mm57z6;
wire Um57z6, Cn57z6, Kn57z6, Sn57z6, Ao57z6, Io57z6, Qo57z6, Yo57z6, Gp57z6, Op57z6;
wire Wp57z6, Eq57z6, Mq57z6, Uq57z6, Cr57z6, Kr57z6, Sr57z6, As57z6, Is57z6, Qs57z6;
wire Ys57z6, Gt57z6, Ot57z6, Wt57z6, Eu57z6, Mu57z6, Uu57z6, Cv57z6, Kv57z6, Sv57z6;
wire Aw57z6, Iw57z6, Qw57z6, Yw57z6, Gx57z6, Ox57z6, Wx57z6, Ey57z6, My57z6, Uy57z6;
wire Cz57z6, Kz57z6, Sz57z6, A067z6, I067z6, Q067z6, Y067z6, G167z6, O167z6, W167z6;
wire E267z6, M267z6, U267z6, C367z6, K367z6, S367z6, A467z6, I467z6, Q467z6, Y467z6;
wire G567z6, O567z6, W567z6, E667z6, M667z6, U667z6, C767z6, K767z6, S767z6, A867z6;
wire I867z6, Q867z6, Y867z6, G967z6, O967z6, W967z6, Ea67z6, Ma67z6, Ua67z6, Cb67z6;
wire Kb67z6, Sb67z6, Ac67z6, Ic67z6, Qc67z6, Yc67z6, Gd67z6, Od67z6, Wd67z6, Ee67z6;
wire Me67z6, Ue67z6, Cf67z6, Kf67z6, Sf67z6, Ag67z6, Ig67z6, Qg67z6, Yg67z6, Gh67z6;
wire Oh67z6, Wh67z6, Ei67z6, Mi67z6, Ui67z6, Cj67z6, Kj67z6, Sj67z6, Ak67z6, Ik67z6;
wire Qk67z6, Yk67z6, Gl67z6, Ol67z6, Wl67z6, Em67z6, Mm67z6, Um67z6, Cn67z6, Kn67z6;
wire Sn67z6, Ao67z6, Io67z6, Qo67z6, Yo67z6, Gp67z6, Op67z6, Wp67z6, Eq67z6, Mq67z6;
wire Uq67z6, Cr67z6, Kr67z6, Sr67z6, As67z6, Is67z6, Qs67z6, Ys67z6, Gt67z6, Ot67z6;
wire Wt67z6, Eu67z6, Mu67z6, Uu67z6, Cv67z6, Kv67z6, Sv67z6, Aw67z6, Iw67z6, Qw67z6;
wire Yw67z6, Gx67z6, Ox67z6, Wx67z6, Ey67z6, My67z6, Uy67z6, Cz67z6, Kz67z6, Sz67z6;
wire A077z6, I077z6, Q077z6, Y077z6, G177z6, O177z6, W177z6, E277z6, M277z6, U277z6;
wire C377z6, K377z6, S377z6, A477z6, I477z6, Q477z6, Y477z6, G577z6, O577z6, W577z6;
wire E677z6, M677z6, U677z6, C777z6, K777z6, S777z6, A877z6, I877z6, Q877z6, Y877z6;
wire G977z6, O977z6, W977z6, Ea77z6, Ma77z6, Ua77z6, Cb77z6, Kb77z6, Sb77z6, Ac77z6;
wire Ic77z6, Qc77z6, Yc77z6, Gd77z6, Od77z6, Wd77z6, Ee77z6, Me77z6, Ue77z6, Cf77z6;
wire Kf77z6, Sf77z6, Ag77z6, Ig77z6, Qg77z6, Yg77z6, Gh77z6, Oh77z6, Wh77z6, Ei77z6;
wire Mi77z6, Ui77z6, Cj77z6, Kj77z6, Sj77z6, Ak77z6, Ik77z6, Qk77z6, Yk77z6, Gl77z6;
wire Ol77z6, Wl77z6, Em77z6, Mm77z6, Um77z6, Cn77z6, Kn77z6, Sn77z6, Ao77z6, Io77z6;
wire Qo77z6, Yo77z6, Gp77z6, Op77z6, Wp77z6, Eq77z6, Mq77z6, Uq77z6, Cr77z6, Kr77z6;
wire Sr77z6, As77z6, Is77z6, Qs77z6, Ys77z6, Gt77z6, Ot77z6, Wt77z6, Eu77z6, Mu77z6;
wire Uu77z6, Cv77z6, Kv77z6, Sv77z6, Aw77z6, Iw77z6, Qw77z6, Yw77z6, Gx77z6, Ox77z6;
wire Wx77z6, Ey77z6, My77z6, Uy77z6, Cz77z6, Kz77z6, Sz77z6, A087z6, I087z6, Q087z6;
wire Y087z6, G187z6, O187z6, W187z6, E287z6, M287z6, U287z6, C387z6, K387z6, S387z6;
wire A487z6, I487z6, Q487z6, Y487z6, G587z6, O587z6, W587z6, E687z6, M687z6, U687z6;
wire C787z6, K787z6, S787z6, A887z6, I887z6, Q887z6, Y887z6, G987z6, O987z6, W987z6;
wire Ea87z6, Ma87z6, Ua87z6, Cb87z6, Kb87z6, Sb87z6, Ac87z6, Ic87z6, Qc87z6, Yc87z6;
wire Gd87z6, Od87z6, Wd87z6, Ee87z6, Me87z6, Ue87z6, Cf87z6, Kf87z6, Sf87z6, Ag87z6;
wire Ig87z6, Qg87z6, Yg87z6, Gh87z6, Oh87z6, Wh87z6, Ei87z6, Mi87z6, Ui87z6, Cj87z6;
wire Kj87z6, Sj87z6, Ak87z6, Ik87z6, Qk87z6, Yk87z6, Gl87z6, Ol87z6, Wl87z6, Em87z6;
wire Mm87z6, Um87z6, Cn87z6, Kn87z6, Sn87z6, Ao87z6, Io87z6, Qo87z6, Yo87z6, Gp87z6;
wire Op87z6, Wp87z6, Eq87z6, Mq87z6, Uq87z6, Cr87z6, Kr87z6, Sr87z6, As87z6, Is87z6;
wire Qs87z6, Ys87z6, Gt87z6, Ot87z6, Wt87z6, Eu87z6, Mu87z6, Uu87z6, Cv87z6, Kv87z6;
wire Sv87z6, Aw87z6, Iw87z6, Qw87z6, Yw87z6, Gx87z6, Ox87z6, Wx87z6, Ey87z6, My87z6;
wire Uy87z6, Cz87z6, Kz87z6, Sz87z6, A097z6, I097z6, Q097z6, Y097z6, G197z6, O197z6;
wire W197z6, E297z6, M297z6, U297z6, C397z6, K397z6, S397z6, A497z6, I497z6, Q497z6;
wire Y497z6, G597z6, O597z6, W597z6, E697z6, M697z6, U697z6, C797z6, K797z6, S797z6;
wire A897z6, I897z6, Q897z6, Y897z6, G997z6, O997z6, W997z6, Ea97z6, Ma97z6, Ua97z6;
wire Cb97z6, Kb97z6, Sb97z6, Ac97z6, Ic97z6, Qc97z6, Yc97z6, Gd97z6, Od97z6, Wd97z6;
wire Ee97z6, Me97z6, Ue97z6, Cf97z6, Kf97z6, Sf97z6, Ag97z6, Ig97z6, Qg97z6, Yg97z6;
wire Gh97z6, Oh97z6, Wh97z6, Ei97z6, Mi97z6, Ui97z6, Cj97z6, Kj97z6, Sj97z6, Ak97z6;
wire Ik97z6, Qk97z6, Yk97z6, Gl97z6, Ol97z6, Wl97z6, Em97z6, Mm97z6, Um97z6, Cn97z6;
wire Kn97z6, Sn97z6, Ao97z6, Io97z6, Qo97z6, Yo97z6, Gp97z6, Op97z6, Wp97z6, Eq97z6;
wire Mq97z6, Uq97z6, Cr97z6, Kr97z6, Sr97z6, As97z6, Is97z6, Qs97z6, Ys97z6, Gt97z6;
wire Ot97z6, Wt97z6, Eu97z6, Mu97z6, Uu97z6, Cv97z6, Kv97z6, Sv97z6, Aw97z6, Iw97z6;
wire Qw97z6, Yw97z6, Gx97z6, Ox97z6, Wx97z6, Ey97z6, My97z6, Uy97z6, Cz97z6, Kz97z6;
wire Sz97z6, A0a7z6, I0a7z6, Q0a7z6, Y0a7z6, G1a7z6, O1a7z6, W1a7z6, E2a7z6, M2a7z6;
wire U2a7z6, C3a7z6, K3a7z6, S3a7z6, A4a7z6, I4a7z6, Q4a7z6, Y4a7z6, G5a7z6, O5a7z6;
wire W5a7z6, E6a7z6, M6a7z6, U6a7z6, C7a7z6, K7a7z6, S7a7z6, A8a7z6, I8a7z6, Q8a7z6;
wire Y8a7z6, G9a7z6, O9a7z6, W9a7z6, Eaa7z6, Maa7z6, Uaa7z6, Cba7z6, Kba7z6, Sba7z6;
wire Aca7z6, Ica7z6, Qca7z6, Yca7z6, Gda7z6, Oda7z6, Wda7z6, Eea7z6, Mea7z6, Uea7z6;
wire Cfa7z6, Kfa7z6, Sfa7z6, Aga7z6, Iga7z6, Qga7z6, Yga7z6, Gha7z6, Oha7z6, Wha7z6;
wire Eia7z6, Mia7z6, Uia7z6, Cja7z6, Kja7z6, Sja7z6, Aka7z6, Xka7z6, Ula7z6, Rma7z6;
wire Ona7z6, Loa7z6, Ipa7z6, Fqa7z6, Cra7z6, Zra7z6, Xsa7z6, Vta7z6, Tua7z6, Rva7z6;
wire Pwa7z6, Nxa7z6, Lya7z6, Jza7z6, H0b7z6, F1b7z6, D2b7z6, B3b7z6, Z3b7z6, X4b7z6;
wire V5b7z6, T6b7z6, R7b7z6, P8b7z6, N9b7z6, Lab7z6, Jbb7z6, Hcb7z6, Fdb7z6, Deb7z6;
wire Bfb7z6, Zfb7z6, Xgb7z6, Vhb7z6;
wire [63:0] Tib7z6;
wire [66:0] Fjb7z6;
wire [19:2] Pjb7z6;
wire [9:8] Zjb7z6;
wire [2:0] Wkb7z6;
wire [4:0] Tlb7z6;
wire [8:0] Qmb7z6;
wire [31:10] Pnb7z6;
wire [8:0] Nob7z6;
wire [7:5] Ppb7z6;
wire [6:0] Mqb7z6;
wire [1:0] Hrb7z6;
wire [1:0] Gsb7z6;
wire [31:0] Itb7z6;
wire [1:0] Hub7z6;
wire [31:2] Fvb7z6;
wire [5:0] Dwb7z6;
wire [31:0] Kxb7z6;
wire [4:0] Uyb7z6;
wire [1:0] I0c7z6;
wire [31:0] V1c7z6;
wire [4:0] E3c7z6;
wire [3:0] P4c7z6;
wire [4:0] D6c7z6;
wire [8:7] O7c7z6;
wire [3:0] Z8c7z6;
wire [3:0] Oac7z6;
wire [14:3] Ecc7z6;
wire [31:0] Pdc7z6;
wire [31:0] Zec7z6;
wire [3:0] Cgc7z6;
wire [31:5] Fhc7z6;
wire [31:0] Pic7z6;
wire [31:1] Vjc7z6;
wire [31:1] Flc7z6;
wire [2:0] Pmc7z6;
wire [1:0] Lpc7z6;
wire [1:0] Fsc7z6;
wire [31:0] Dvc7z6;
wire [31:0] Byc7z6;
wire [31:2] X0d7z6;
wire [5:0] U3d7z6;
wire [2:0] P6d7z6;
wire [5:0] L9d7z6;
wire [5:0] Gcd7z6;
wire [5:0] Bfd7z6;
wire [31:2] Xhd7z6;
wire [31:1] Wkd7z6;
wire [31:1] Vnd7z6;
wire [22:17] Uqd7z6;
wire [2:1] Osd7z6;
wire [6:0] Gvd7z6;
wire [1:0] Yxd7z6;
wire [5:0] S0e7z6;
wire [1:0] M3e7z6;
wire [1:0] M5e7z6;
wire [1:0] K7e7z6;
wire [2:0] I9e7z6;
wire [4:0] Ibe7z6;
wire [3:0] Ide7z6;
wire [7:3] Mfe7z6;
wire [7:1] Ohe7z6;
wire [31:0] Rje7z6;
wire [7:0] Ple7z6;
wire [1:0] Pne7z6;
wire [5:2] Mpe7z6;
wire [1:0] Fre7z6;
wire [20:0] Dte7z6;
wire [30:0] Cve7z6;
wire [3:0] Xwe7z6;
wire [5:0] Rze7z6;
wire [5:0] K2f7z6;
wire [5:0] D5f7z6;
wire [5:0] S7f7z6;
wire [5:0] Jaf7z6;
wire [3:0] Bdf7z6;
wire [30:0] Uff7z6;
wire [31:0] Kif7z6;
wire [31:0] Alf7z6;
wire [31:0] Onf7z6;
wire [15:0] Cqf7z6;
wire [15:0] Ssf7z6;
wire [15:0] Ivf7z6;
wire [34:0] Yxf7z6;
wire [32:0] L0g7z6;
wire [31:0] X2g7z6;
wire [31:0] J5g7z6;
wire [31:0] V7g7z6;
wire [31:0] Fag7z6;
wire [31:0] Pcg7z6;
wire [32:1] Zfg7z6;
wire [32:1] Jjg7z6;
wire [32:1] Tmg7z6;
wire [32:1] Dqg7z6;
wire [3:0] Ntg7z6;
wire [3:0] Lvg7z6;
wire [3:0] Pxg7z6;
wire [3:0] Nzg7z6;
wire [5:0] Q1h7z6;
wire [1:0] R3h7z6;
wire [3:0] O5h7z6;
wire [3:0] E8h7z6;
wire [5:0] Uah7z6;
wire [1:0] Edh7z6;
wire [1:0] Tfh7z6;
wire [1:0] Kih7z6;
wire [31:0] Zkh7z6;
wire [2:0] Xnh7z6;
wire [31:0] Nqh7z6;
wire [31:0] Fth7z6;
wire [31:0] Vvh7z6;
wire [31:0] Oyh7z6;
wire [31:0] K1i7z6;
wire [9:0] G4i7z6;
wire [1:0] U6i7z6;
wire [9:0] P9i7z6;
wire [1:0] Fci7z6;
wire [3:1] Zei7z6;
wire [31:1] Bhi7z6;
wire [31:1] Eji7z6;
wire [31:1] Gli7z6;
wire [31:1] Bni7z6;
wire [11:2] Toi7z6;
wire [3:0] Bqi7z6;
wire [31:0] Dri7z6;
wire [2:0] Hsi7z6;
wire [9:7] Qti7z6;
wire [31:0] Wui7z6;
wire [31:0] Bwi7z6;
wire [4:0] Bxi7z6;
wire [31:1] Byi7z6;
wire [25:0] Bzi7z6;
wire [23:0] A0j7z6;
wire [23:0] H1j7z6;
wire [6:0] P2j7z6;
wire [15:0] Z3j7z6;
wire [63:0] G5j7z6;
wire [63:0] M6j7z6;
wire [2:0] T7j7z6;
wire [2:0] Z8j7z6;
wire [2:0] Gaj7z6;
wire [2:0] Nbj7z6;
wire [2:0] Tcj7z6;
wire [2:0] Zdj7z6;
wire [2:0] Ffj7z6;
wire [191:0] Lgj7z6;
wire [63:0] Ohj7z6;
wire [6:0] Qij7z6;
wire [63:0] Qkj7z6;
wire [5:1] Qmj7z6;
wire [2:0] Moj7z6;
wire [72:0] Jqj7z6;
wire [5:2] Dtj7z6;
wire [3:0] Pvj7z6;
wire [7:0] Hyj7z6;
wire [31:5] X0k7z6;
wire [31:2] N3k7z6;
wire [31:5] V5k7z6;
wire [7:0] H8k7z6;
wire [23:0] Rbk7z6;
wire [31:5] Dfk7z6;
wire [7:0] Pik7z6;
wire [23:0] Zlk7z6;
wire [24:5] Lpk7z6;
wire [7:0] Xsk7z6;
wire [23:0] Hwk7z6;
wire [24:5] Tzk7z6;
wire [7:0] F3l7z6;
wire [23:0] P6l7z6;
wire [24:5] Bal7z6;
wire [7:0] Ndl7z6;
wire [23:0] Xgl7z6;
wire [31:5] Jkl7z6;
wire [7:0] Vnl7z6;
wire [23:0] Frl7z6;
wire [24:5] Rul7z6;
wire [7:0] Dyl7z6;
wire [23:0] N1m7z6;
wire [24:5] Z4m7z6;
wire [7:0] L8m7z6;
wire [23:0] Vbm7z6;
wire [25:5] Hfm7z6;
wire [31:0] Tim7z6;
wire [1:0] Dkm7z6;
wire [31:0] Cmm7z6;
wire [2:0] Rnm7z6;
wire [2:0] Kqm7z6;
wire [3:0] Dtm7z6;
wire [1:0] Qvm7z6;
wire [3:1] Aym7z6;
wire [1:0] J0n7z6;
wire [1:0] W2n7z6;
wire [3:0] J5n7z6;
wire [1:0] S7n7z6;
wire [4:3] Ean7z6;
wire [31:0] Icn7z6;
wire [2:0] Ven7z6;
wire [31:0] Chn7z6;
wire [31:5] Hjn7z6;
wire [1:0] Qln7z6;
wire [3:0] Znn7z6;
wire [2:0] Eqn7z6;
wire [2:0] Ysn7z6;
wire [2:0] Svn7z6;
wire [2:0] Kyn7z6;
wire [1:0] C1o7z6;
wire [31:4] U3o7z6;
wire [7:2] F5o7z6;
wire [2:0] O7o7z6;
wire [3:0] Y9o7z6;
wire [6:4] Gco7z6;
wire [2:0] Oeo7z6;
wire [1:0] Ugo7z6;
wire [1:0] Ejo7z6;
wire [6:0] Klo7z6;
wire [31:2] Zmo7z6;
wire [31:2] Coo7z6;
wire [26:0] Fpo7z6;
wire [26:0] Nqo7z6;
wire [26:0] Vro7z6;
wire [1:0] Dto7z6;
wire [26:0] Ouo7z6;
wire [1:0] Wvo7z6;
wire [26:0] Hxo7z6;
wire [1:0] Pyo7z6;
wire [26:0] A0p7z6;
wire [1:0] I1p7z6;
wire [28:2] T2p7z6;
wire [28:2] W3p7z6;
wire [5:0] Z4p7z6;
wire [31:0] E6p7z6;
wire [3:0] I7p7z6;
wire [3:0] Q8p7z6;
wire [31:0] U9p7z6;
wire [1:0] Bbp7z6;
wire [1:0] Ncp7z6;
wire [3:0] Zdp7z6;
wire [3:0] Lfp7z6;
wire [3:0] Sgp7z6;
wire [3:0] Rip7z6;
wire [31:0] Mkp7z6;
wire [3:0] Hmp7z6;
wire [3:0] Gop7z6;
wire [31:0] Bqp7z6;
wire [1:0] Wrp7z6;
wire [1:0] Bup7z6;
wire [1:0] Gwp7z6;
wire [3:0] Hyp7z6;
wire [3:0] G0q7z6;
wire [31:0] B2q7z6;
wire [3:0] W3q7z6;
wire [1:0] W5q7z6;
wire [3:0] Y7q7z6;
wire [3:0] X9q7z6;
wire [7:0] Tbq7z6;
wire [7:0] Pdq7z6;
wire [7:0] Kfq7z6;
wire [7:0] Hhq7z6;
wire [7:0] Cjq7z6;
wire [22:12] Xkq7z6;
wire [6:3] Nmq7z6;
wire [14:1] Hoq7z6;
wire [14:0] Gqq7z6;
wire [31:0] Gsq7z6;
wire [14:1] Luq7z6;
wire [14:0] Kwq7z6;
wire [14:0] Kyq7z6;
wire [14:1] P0r7z6;
wire [14:0] O2r7z6;
wire [14:0] O4r7z6;
wire [31:1] T6r7z6;
wire [14:0] S8r7z6;
wire [31:0] Sar7z6;
wire [1:0] Xcr7z6;
wire [1:0] Dfr7z6;
wire [1:0] Jhr7z6;
wire [10:0] Tjr7z6;
wire [31:0] Wlr7z6;
wire [31:0] Cor7z6;
wire [31:1] Gqr7z6;
wire [1:0] Hsr7z6;
wire [1:0] Uur7z6;
wire [1:0] Ixr7z6;
wire [31:1] Rzr7z6;
wire [5:0] V1s7z6;
wire [1:0] C4s7z6;
wire [1:0] M6s7z6;
wire [30:8] P7s7z6;
wire [1:0] R8s7z6;
wire [39:0] X9s7z6;
wire [2:0] Zas7z6;
wire [3:0] Scs7z6;
wire [31:0] Ies7z6;
wire [11:7] Zfs7z6;
wire [3:0] Ihs7z6;
wire [5:0] Vis7z6;
wire [4:0] Nks7z6;
wire [8:0] Kms7z6;
wire [8:0] Cnvmz6;
wire [8:0] Xovmz6;
wire [8:0] Sqvmz6;
wire [8:0] Nsvmz6;
wire [8:4] Iuvmz6;
wire [4:0] Kwvmz6;
wire [8:0] Gyvmz6;
wire [8:0] K0wmz6;
wire [1:0] O2wmz6;
wire [1:0] Y4wmz6;
wire [8:0] J7wmz6;
wire [8:0] N9wmz6;
wire [1:0] Rbwmz6;
wire [1:0] Bewmz6;
wire [8:0] Mgwmz6;
wire [8:0] Qiwmz6;
wire [1:0] Ukwmz6;
wire [1:0] Enwmz6;
wire [8:0] Ppwmz6;
wire [8:0] Trwmz6;
wire [1:0] Xtwmz6;
wire [1:0] Hwwmz6;
wire [8:0] Sywmz6;
wire [8:0] W0xmz6;
wire [1:0] A3xmz6;
wire [1:0] K5xmz6;
wire [7:0] V7xmz6;
wire [2:0] O9xmz6;
wire [3:0] Fbxmz6;
wire [47:0] Vcxmz6;
wire [31:0] Jexmz6;
wire [11:0] Tfxmz6;
wire [3:0] Ogxmz6;
wire [1:0] Hhxmz6;
wire [31:0] Aixmz6;
wire [31:2] Uixmz6;
wire [11:0] Njxmz6;
wire [3:0] Ikxmz6;
wire [1:0] Blxmz6;
wire [31:0] Ulxmz6;
wire [31:2] Omxmz6;
wire [11:0] Hnxmz6;
wire [31:0] Coxmz6;
wire [5:0] Woxmz6;
wire [5:0] Fqxmz6;
wire [31:0] Krxmz6;
wire [1:0] Usxmz6;
wire [1:0] Fuxmz6;
wire [1:0] Ovxmz6;
wire [31:0] Cxxmz6;
wire [4:0] Myxmz6;
wire [4:0] Uzxmz6;
wire [5:0] B1ymz6;
wire [1:0] Q2ymz6;
wire [3:0] Z3ymz6;
wire [34:0] L5ymz6;
wire [3:0] W6ymz6;
wire [3:0] G8ymz6;
wire [3:0] R9ymz6;
wire [1:0] Dbymz6;
wire [4:1] Hcymz6;
wire [3:0] Jdymz6;
wire [3:0] Feymz6;
wire [2:0] Bfymz6;
wire [11:2] Xfymz6;
wire [10:0] Sgymz6;
wire [15:0] Biymz6;
wire [10:0] Ojymz6;
wire [3:0] Blymz6;
wire [3:0] Kmymz6;
wire [10:0] Unymz6;
wire [1:0] Ipymz6;
wire [1:0] Drymz6;
wire [15:0] Ctymz6;
wire [15:0] Ruymz6;
wire [3:0] Iwymz6;
wire [8:0] Zxymz6;
wire [3:0] Vzymz6;
wire [35:7] T1zmz6;
wire [31:7] P3zmz6;
wire [31:1] L5zmz6;
wire [31:1] I7zmz6;
wire [1:0] W8zmz6;
wire [8:0] Pazmz6;
wire [3:0] Lczmz6;
wire [35:1] Jezmz6;
wire [1:0] Fgzmz6;
wire [4:0] Yhzmz6;
wire [31:1] Rjzmz6;
wire [31:1] Slzmz6;
wire [46:0] Gnzmz6;
wire [7:0] Xozmz6;
wire [7:0] Nqzmz6;
wire [7:0] Dszmz6;
wire [7:0] Ttzmz6;
wire [7:0] Jvzmz6;
wire [7:0] Zwzmz6;
wire [7:0] Pyzmz6;
wire [7:0] F00nz6;
wire [7:0] V10nz6;
wire [7:0] L30nz6;
wire [7:0] B50nz6;
wire [7:0] R60nz6;
wire [7:0] H80nz6;
wire [7:0] X90nz6;
wire [7:0] Nb0nz6;
wire [7:0] Dd0nz6;
wire [7:0] Te0nz6;
wire [7:0] Jg0nz6;
wire [7:0] Zh0nz6;
wire [7:0] Pj0nz6;
wire [7:0] Fl0nz6;
wire [7:0] Vm0nz6;
wire [7:0] Lo0nz6;
wire [7:0] Bq0nz6;
wire [1:0] Rr0nz6;
wire [4:0] Ft0nz6;
wire [4:0] Uu0nz6;
wire [2:1] Hw0nz6;
wire [2:0] Ux0nz6;
wire [4:3] Mz0nz6;
wire [4:0] E11nz6;
wire [2:0] R21nz6;
wire [1:0] B41nz6;
wire [2:0] T51nz6;
wire [8:0] H71nz6;
wire [2:0] U81nz6;
wire [2:0] Ja1nz6;
wire [2:0] Yb1nz6;
wire [2:0] Md1nz6;
wire [2:0] Af1nz6;
wire [2:0] Fg1nz6;
wire [7:2] Kh1nz6;
wire [2:0] Hi1nz6;
wire [2:0] Lj1nz6;
wire [12:0] Pk1nz6;
wire [1:0] Nl1nz6;
wire [7:0] Mm1nz6;
wire [7:0] Nn1nz6;
wire [7:0] Oo1nz6;
wire [1:0] Pp1nz6;
wire [7:2] Xq1nz6;
wire [7:0] Yr1nz6;
wire [7:0] Zs1nz6;
wire [7:0] Au1nz6;
wire [1:0] Bv1nz6;
wire [3:0] Jw1nz6;
wire [1:0] Iy1nz6;
wire [11:2] J02nz6;
wire [7:0] Z12nz6;
wire [3:0] T32nz6;
wire [6:0] N52nz6;
wire [7:0] J72nz6;
wire [1:0] D92nz6;
wire [1:0] Qa2nz6;
wire [3:0] Ec2nz6;
wire [12:0] Td2nz6;
wire [2:0] Kf2nz6;
wire [2:0] Ah2nz6;
wire [5:0] Ti2nz6;
reg Sj2nz6, Ik2nz6, Zk2nz6, Ql2nz6, Im2nz6, Ym2nz6, Pn2nz6, Go2nz6, Yo2nz6, Eq2nz6;
reg Er2nz6, Hs2nz6, Et2nz6, Su2nz6, Aw2nz6, Ny2nz6, A13nz6, N33nz6, A63nz6, N83nz6;
reg Ab3nz6, Cd3nz6, Bf3nz6, Yg3nz6, Xh3nz6, Vj3nz6, Ul3nz6, Un3nz6, Ip3nz6, Vq3nz6;
reg Ms3nz6, Su3nz6, Mw3nz6, Sx3nz6, T04nz6, D34nz6, B64nz6, P84nz6, Ab4nz6, Pd4nz6;
reg Jf4nz6, Jh4nz6, Jj4nz6, Hl4nz6, Un4nz6, Nq4nz6, Gt4nz6, Yv4nz6, My4nz6, L15nz6;
reg R45nz6, H65nz6, G95nz6, Kc5nz6, Jf5nz6, Mi5nz6, Kl5nz6, Ho5nz6, Qq5nz6, Rs5nz6;
reg Ou5nz6, Zw5nz6, Oz5nz6, O16nz6, M36nz6, N66nz6, X86nz6, Vb6nz6, Pe6nz6, Jh6nz6;
reg Dk6nz6, Ym6nz6, Tp6nz6, Os6nz6, Jv6nz6, Ey6nz6, Z07nz6, A37nz6, P57nz6, H87nz6;
reg Z97nz6, Oc7nz6, Af7nz6, Qh7nz6, Fk7nz6, Cn7nz6, Cq7nz6, Ls7nz6, Jv7nz6, Dy7nz6;
reg X08nz6, S38nz6, N68nz6, I98nz6, Dc8nz6, Ye8nz6, Th8nz6, Uj8nz6, Rl8nz6, Co8nz6;
reg Rq8nz6, Rs8nz6, Pu8nz6, Qx8nz6, A09nz6, X29nz6, R59nz6, P89nz6, Lb9nz6, Le9nz6;
reg Oh9nz6, Ik9nz6, Gn9nz6, Fq9nz6, Ct9nz6, Av9nz6, Zv9nz6, Zw9nz6, Zx9nz6, Zy9nz6;
reg Zz9nz6, Z0anz6, Z1anz6, Z2anz6, Z3anz6, Z4anz6, A6anz6, B7anz6, C8anz6, D9anz6;
reg Eaanz6, Fbanz6, Gcanz6, Hdanz6, Ieanz6, Jfanz6, Kganz6, Lhanz6, Mianz6, Njanz6;
reg Okanz6, Planz6, Qmanz6, Rnanz6, Soanz6, Tpanz6, Uqanz6, Vranz6, Wsanz6, Xtanz6;
reg Yuanz6, Zvanz6, Axanz6, Byanz6, Czanz6, D0bnz6, E1bnz6, F2bnz6, G3bnz6, H4bnz6;
reg I5bnz6, J6bnz6, K7bnz6, L8bnz6, M9bnz6, Nabnz6, Obbnz6, Pcbnz6, Qdbnz6, Rebnz6;
reg Sfbnz6, Tgbnz6, Uhbnz6, Vibnz6, Wjbnz6, Xkbnz6, Ylbnz6, Zmbnz6, Aobnz6, Bpbnz6;
reg Cqbnz6, Drbnz6, Dsbnz6, Etbnz6, Fwbnz6, Hzbnz6, J2cnz6, L5cnz6, N8cnz6, Pbcnz6;
reg Recnz6, Thcnz6, Vkcnz6, Xncnz6, Zqcnz6, Bucnz6, Dxcnz6, F0dnz6, H3dnz6, J6dnz6;
reg L9dnz6, Ncdnz6, Pfdnz6, Ridnz6, Tldnz6, Vodnz6, Xrdnz6, Zudnz6, Bydnz6, D1enz6;
reg F4enz6, H7enz6, Jaenz6, Ldenz6, Ngenz6, Pjenz6, Rmenz6, Tpenz6, Vsenz6, Xvenz6;
reg Zyenz6, B2fnz6, D5fnz6, F8fnz6, Hbfnz6, Jefnz6, Lhfnz6, Nkfnz6, Pnfnz6, Rqfnz6;
reg Ttfnz6, Vwfnz6, Xzfnz6, Z2gnz6, B6gnz6, D9gnz6, Fcgnz6, Hfgnz6, Jignz6, Llgnz6;
reg Nognz6, Prgnz6, Rugnz6, Txgnz6, V0hnz6, X3hnz6, Z6hnz6, Bahnz6, Cdhnz6, Dghnz6;
reg Bjhnz6, Elhnz6, Cnhnz6, Hphnz6, Yrhnz6, Tuhnz6, Zxhnz6, Pzhnz6, O2inz6, S5inz6;
reg Q8inz6, Vainz6, Xdinz6, Zginz6, Bkinz6, Dninz6, Tpinz6, Osinz6, Kvinz6, Myinz6;
reg O1jnz6, N3jnz6, S5jnz6, Q7jnz6, P9jnz6, Objnz6, Qdjnz6, Wfjnz6, Bijnz6, Fkjnz6;
reg Gmjnz6, Qojnz6, Qrjnz6, Ztjnz6, Fxjnz6, Lzjnz6, P2knz6, D5knz6, O7knz6, Daknz6;
reg Dcknz6, Beknz6, Chknz6, Mjknz6, Kmknz6, Qoknz6, Vqknz6, Mtknz6, Jwknz6, Pzknz6;
reg J2lnz6, L5lnz6, L8lnz6, Ualnz6, Rdlnz6, Pglnz6, Uilnz6, Dllnz6, Aolnz6, Arlnz6;
reg Fulnz6, Exlnz6, Azlnz6, A1mnz6, X3mnz6, X6mnz6, G9mnz6, Qbmnz6, Zdmnz6, Wgmnz6;
reg Wjmnz6, Cnmnz6, Zpmnz6, Wsmnz6, Xvmnz6, Yymnz6, Z1nnz6, X4nnz6, T7nnz6, N9nnz6;
reg Gbnnz6, Wcnnz6, Sennz6, Dhnnz6, Sjnnz6, Plnnz6, Mnnnz6, Kpnnz6, Lsnnz6, Vunnz6;
reg Txnnz6, Vznnz6, W2onz6, G5onz6, E8onz6, U9onz6, Nbonz6, Ceonz6, Sgonz6, Ijonz6;
reg Xlonz6, Voonz6, Yronz6, Xuonz6, Cxonz6, Mzonz6, M2pnz6, V4pnz6, S7pnz6, P9pnz6;
reg Acpnz6, Pepnz6, Pgpnz6, Nipnz6, Olpnz6, Ynpnz6, Wqpnz6, Etpnz6, Svpnz6, Dypnz6;
reg S0qnz6, S2qnz6, Q4qnz6, R7qnz6, Baqnz6, Zcqnz6, Xfqnz6, Viqnz6, Zkqnz6, Ynqnz6;
reg Cqqnz6, Atqnz6, Evqnz6, Dyqnz6, H0rnz6, G3rnz6, K5rnz6, O8rnz6, Pbrnz6, Zdrnz6;
reg Xgrnz6, Yirnz6, Zlrnz6, Jornz6, Hrrnz6, Ntrnz6, Tvrnz6, Uyrnz6, E1snz6, C4snz6;
reg F6snz6, F8snz6, Hasnz6, Fcsnz6, Jesnz6, Hhsnz6, Kksnz6, Xmsnz6, Ypsnz6, Etsnz6;
reg Ewsnz6, Dzsnz6, H2tnz6, G5tnz6, M7tnz6, W9tnz6, Uctnz6, Oetnz6, Mgtnz6, Kitnz6;
reg Jktnz6, Hmtnz6, Fotnz6, Dqtnz6, Bstnz6, Wttnz6, Uvtnz6, Hytnz6, A1unz6, T3unz6;
reg G6unz6, Z8unz6, Sbunz6, Qdunz6, Ofunz6, Mhunz6, Kjunz6, Kmunz6, Tounz6, Qrunz6;
reg Stunz6, Uwunz6, Vzunz6, W2vnz6, U5vnz6, Y7vnz6, Cavnz6, Ccvnz6, Tevnz6, Khvnz6;
reg Pkvnz6, Smvnz6, Rovnz6, Prvnz6, Stvnz6, Wvvnz6, Yyvnz6, D1wnz6, N3wnz6, O5wnz6;
reg Q7wnz6, Rawnz6, Bdwnz6, Zfwnz6, Fiwnz6, Lkwnz6, Mnwnz6, Eqwnz6, Oswnz6, Yuwnz6;
reg Wxwnz6, Mzwnz6, K2xnz6, L5xnz6, V7xnz6, Baxnz6, Hcxnz6, Ifxnz6, Shxnz6, Qkxnz6;
reg Wmxnz6, Cpxnz6, Drxnz6, Ftxnz6, Gwxnz6, Qyxnz6, O1ynz6, L3ynz6, J5ynz6, E7ynz6;
reg Y8ynz6, Ebynz6, Kdynz6, Gfynz6, Chynz6, Yiynz6, Xkynz6, Rmynz6, Hoynz6, Gqynz6;
reg Gsynz6, Guynz6, Gwynz6, Gyynz6, G0znz6, Y2znz6, J5znz6, B8znz6, Maznz6, Xcznz6;
reg Ifznz6, Aiznz6, Skznz6, Dnznz6, Kpznz6, Isznz6, Jvznz6, Txznz6, R00oz6, P30oz6;
reg T50oz6, T70oz6, Ba0oz6, Ec0oz6, Ge0oz6, Jg0oz6, Ki0oz6, Ek0oz6, Em0oz6, Io0oz6;
reg Sq0oz6, Qs0oz6, Wu0oz6, Xw0oz6, Yy0oz6, V01oz6, Q21oz6, O41oz6, M61oz6, O81oz6;
reg Ra1oz6, Md1oz6, Eg1oz6, Ji1oz6, Pk1oz6, Ln1oz6, Qp1oz6, Or1oz6, Zt1oz6, Wv1oz6;
reg Jx1oz6, Oz1oz6, H12oz6, H32oz6, H52oz6, E72oz6, Z82oz6, Xa2oz6, Vc2oz6, Df2oz6;
reg Eh2oz6, Gj2oz6, Lm2oz6, Ip2oz6, Fs2oz6, Cv2oz6, Sx2oz6, J03oz6, A33oz6, Q53oz6;
reg Z73oz6, Ja3oz6, Hd3oz6, Tg3oz6, Sj3oz6, Lm3oz6, Mp3oz6, Wr3oz6, Uu3oz6, Ww3oz6;
reg Wy3oz6, A14oz6, J34oz6, S54oz6, B84oz6, Ka4oz6, Hc4oz6, Ce4oz6, Ag4oz6, Yh4oz6;
reg Ak4oz6, Dm4oz6, Vo4oz6, Ds4oz6, Gv4oz6, Ky4oz6, O15oz6, R45oz6, V75oz6, Za5oz6;
reg Ce5oz6, Fh5oz6, Jk5oz6, Nn5oz6, Qq5oz6, Ut5oz6, Yw5oz6, B06oz6, E36oz6, D66oz6;
reg A96oz6, Db6oz6, Hd6oz6, Ig6oz6, Jj6oz6, Mm6oz6, Pp6oz6, Rr6oz6, Yt6oz6, Ow6oz6;
reg Fz6oz6, O17oz6, O47oz6, O77oz6, Ka7oz6, Gd7oz6, Hf7oz6, Li7oz6, Kl7oz6, No7oz6;
reg Pr7oz6, Tu7oz6, Rx7oz6, U08oz6, T38oz6, V58oz6, X78oz6, Aa8oz6, Sc8oz6, Sf8oz6;
reg Ui8oz6, Xk8oz6, Ko8oz6, Hr8oz6, Vt8oz6, Jw8oz6, Mz8oz6, P29oz6, O59oz6, S89oz6;
reg Qb9oz6, Vd9oz6, Ng9oz6, Qj9oz6, Ql9oz6, Nn9oz6, Up9oz6, Zr9oz6, Gu9oz6, Gw9oz6;
reg Gy9oz6, G0aoz6, G2aoz6, B4aoz6, Z5aoz6, X7aoz6, Z9aoz6, Bcaoz6, Xeaoz6, Chaoz6;
reg Bkaoz6, Anaoz6, Wpaoz6, Bsaoz6, Avaoz6, Zxaoz6, R0boz6, G3boz6, K6boz6, O9boz6;
reg Ncboz6, Rfboz6, Qiboz6, Plboz6, Foboz6, Zqboz6, Qtboz6, Jwboz6, Wyboz6, Y1coz6;
reg Y3coz6, Q6coz6, L8coz6, Eacoz6, Xbcoz6, Qdcoz6, Jfcoz6, Chcoz6, Vicoz6, Okcoz6;
reg Hmcoz6, Aocoz6, Cqcoz6, Xrcoz6, Aucoz6, Pvcoz6, Fxcoz6, Vycoz6, J0doz6, X1doz6;
reg T3doz6, P5doz6, L7doz6, H9doz6, Dbdoz6, Zcdoz6, Vedoz6, Rgdoz6, Nidoz6, Jkdoz6;
reg Fmdoz6, Bodoz6, Updoz6, Nrdoz6, Gtdoz6, Zudoz6, Nwdoz6, Fydoz6, Xzdoz6, P1eoz6;
reg H3eoz6, Y4eoz6, P6eoz6, G8eoz6, X9eoz6, Nbeoz6, Edeoz6, Veeoz6, Ngeoz6, Djeoz6;
reg Ykeoz6, Rmeoz6, Koeoz6, Dqeoz6, Wreoz6, Pteoz6, Hveoz6, Zweoz6, Ryeoz6, I0foz6;
reg M2foz6, Q4foz6, U6foz6, Y8foz6, Cbfoz6, Gdfoz6, Lffoz6, Qhfoz6, Vjfoz6, Amfoz6;
reg Fofoz6, Kqfoz6, Psfoz6, Uufoz6, Zwfoz6, Ezfoz6, J1goz6, V2goz6, K4goz6, A6goz6;
reg X7goz6, V9goz6, Nbgoz6, Jdgoz6, Gfgoz6, Sggoz6, Ligoz6, Ckgoz6, Rlgoz6, Jngoz6;
reg Ipgoz6, Irgoz6, Ctgoz6, Evgoz6, Wwgoz6, Oygoz6, P0hoz6, A2hoz6, L3hoz6, Z5hoz6;
reg P8hoz6, Abhoz6, Uchoz6, Jehoz6, Wfhoz6, Ohhoz6, Cjhoz6, Ukhoz6, Imhoz6, Dohoz6;
reg Sphoz6, Wqhoz6, Urhoz6, Sthoz6, Rvhoz6, Kxhoz6, Pzhoz6, F2ioz6, X4ioz6, W7ioz6;
reg Faioz6, Mcioz6, Veioz6, Xhioz6, Xkioz6, Xnioz6, Arioz6, Utioz6, Twioz6, Pzioz6;
reg L2joz6, N5joz6, F8joz6, Fbjoz6, Jdjoz6, Cgjoz6, Eijoz6, Wkjoz6, Nnjoz6, Wpjoz6;
reg Yrjoz6, Yujoz6, Fxjoz6, Lzjoz6, R1koz6, X3koz6, D6koz6, J8koz6, Pakoz6, Vckoz6;
reg Bfkoz6, Hhkoz6, Ojkoz6, Vlkoz6, Cokoz6, Jqkoz6, Qskoz6, Xukoz6, Exkoz6, Lzkoz6;
reg S1loz6, Z3loz6, G6loz6, N8loz6, Ualoz6, Bdloz6, Ifloz6, Phloz6, Wjloz6, Gmloz6;
reg Eploz6, Srloz6, Vuloz6, Yxloz6, X0moz6, B4moz6, Z6moz6, W9moz6, Tcmoz6, Ufmoz6;
reg Dimoz6, Kkmoz6, Mmmoz6, Gpmoz6, Krmoz6, Ptmoz6, Tvmoz6, Wxmoz6, J0noz6, W2noz6;
reg G5noz6, Y6noz6, N8noz6, Eanoz6, Wbnoz6, Menoz6, Dhnoz6, Vjnoz6, Kmnoz6, Opnoz6;
reg Ssnoz6, Qvnoz6, Tynoz6, S1ooz6, S3ooz6, R5ooz6, O8ooz6, Kbooz6, Deooz6, Sgooz6;
reg Kjooz6, Flooz6, Xmooz6, Poooz6, Dqooz6, Yrooz6, Ltooz6, Yuooz6, Twooz6, Nyooz6;
reg E0poz6, V1poz6, O3poz6, C5poz6, U6poz6, M8poz6, Eapoz6, Wbpoz6, Ndpoz6, Efpoz6;
reg Wgpoz6, Mjpoz6, Zlpoz6, Nopoz6, Drpoz6, Ntpoz6, Fwpoz6, Yypoz6, L1qoz6, A4qoz6;
reg S6qoz6, J9qoz6, Bcqoz6, Vdqoz6, Mfqoz6, Dhqoz6, Fjqoz6, Zlqoz6, Qoqoz6, Grqoz6;
reg Ytqoz6, Tvqoz6, Lxqoz6, Dzqoz6, U0roz6, K2roz6, Y3roz6, M5roz6, A7roz6, O8roz6;
reg Earoz6, Ubroz6, Pdroz6, Bfroz6, Ogroz6, Hiroz6, Ujroz6, Wlroz6, Ynroz6, Aqroz6;
reg Csroz6, Furoz6, Iwroz6, Lyroz6, O0soz6, E3soz6, W5soz6, Z7soz6, Pasoz6, Hdsoz6;
reg Kfsoz6, Aisoz6, Sksoz6, Vmsoz6, Xosoz6, Pqsoz6, Hssoz6, Ttsoz6, Ivsoz6, Zwsoz6;
reg Bzsoz6, E1toz6, Z2toz6, C5toz6, U6toz6, X8toz6, Nbtoz6, Fetoz6, Xftoz6, Aitoz6;
reg Qktoz6, Odazz6, Gfazz6, Jhazz6, Ljazz6, Flazz6, Gnazz6, Zoazz6, Erazz6, Utazz6;
reg Mwazz6, Fyazz6, K0bzz6, L2bzz6, F4bzz6, H6bzz6, Z7bzz6, Cabzz6, Scbzz6, Kfbzz6;
reg Chbzz6, Fjbzz6, Hlbzz6, Bnbzz6, Cpbzz6, Vqbzz6, Atbzz6, Qvbzz6, Iybzz6, B0czz6;
reg G2czz6, H4czz6, B6czz6, D8czz6, V9czz6, Ybczz6, Oeczz6, Ghczz6, Yiczz6, Blczz6;
reg Dnczz6, Xoczz6, Yqczz6, Rsczz6, Wuczz6, Mxczz6, E0dzz6, X1dzz6, C4dzz6, D6dzz6;
reg X7dzz6, Z9dzz6, Rbdzz6, Uddzz6, Kgdzz6, Cjdzz6, Ukdzz6, Xmdzz6, Zodzz6, Tqdzz6;
reg Usdzz6, Nudzz6, Swdzz6, Izdzz6, A2ezz6, T3ezz6, Y5ezz6, Z7ezz6, T9ezz6, Vbezz6;
reg Ndezz6, Qfezz6, Giezz6, Ykezz6, Qmezz6, Toezz6, Vqezz6, Psezz6, Quezz6, Jwezz6;
reg Oyezz6, E1fzz6, W3fzz6, P5fzz6, U7fzz6, Kafzz6, Cdfzz6, Yefzz6, Vhfzz6, Pkfzz6;
reg Cnfzz6, Ppfzz6, Dsfzz6, Wufzz6, Jxfzz6, Xzfzz6, P2gzz6, P5gzz6, D8gzz6, Dbgzz6;
reg Degzz6, Dhgzz6, Dkgzz6, Cngzz6, Wpgzz6, Msgzz6, Jvgzz6, Bygzz6, D1hzz6, D4hzz6;
reg D7hzz6, Gahzz6, Jdhzz6, Ighzz6, Mjhzz6, Kmhzz6, Tohzz6, Prhzz6, Duhzz6, Rwhzz6;
reg Jzhzz6, D1izz6, U2izz6, L4izz6, N6izz6, Q8izz6, Haizz6, Ybizz6, Ldizz6, Dfizz6;
reg Hhizz6, Ziizz6, Dlizz6, Vmizz6, Zoizz6, Rqizz6, Vsizz6, Nuizz6, Ewizz6, Uyizz6;
reg M0jzz6, D2jzz6, X4jzz6, N7jzz6, Fajzz6, Zcjzz6, Mfjzz6, Bijzz6, Rkjzz6, Bnjzz6;
reg Xpjzz6, Osjzz6, Fvjzz6, Rxjzz6, H0kzz6, Y2kzz6, O5kzz6, G7kzz6, I9kzz6, Kbkzz6;
reg Ndkzz6, Qfkzz6, Thkzz6, Wjkzz6, Plkzz6, Knkzz6, Fpkzz6, Xqkzz6, Zskzz6, Qukzz6;
reg Gwkzz6, Wxkzz6, Mzkzz6, C1lzz6, S2lzz6, I4lzz6, Y5lzz6, S7lzz6, M9lzz6, Cclzz6;
reg Xdlzz6, Pflzz6, Khlzz6, Cjlzz6, Xklzz6, Pmlzz6, Holzz6, Kqlzz6, Atlzz6, Svlzz6;
reg Gylzz6, S0mzz6, L3mzz6, B6mzz6, R8mzz6, Hbmzz6, Wdmzz6, Igmzz6, Mjmzz6, Qmmzz6;
reg Lpmzz6, Ksmzz6, Jvmzz6, Iymzz6, K1nzz6, B4nzz6, V6nzz6, P9nzz6, Jcnzz6, Dfnzz6;
reg Vhnzz6, Nknzz6, Cnnzz6, Upnzz6, Ysnzz6, Cwnzz6, Rynzz6, J1ozz6, E3ozz6, W4ozz6;
reg O6ozz6, R8ozz6, Hbozz6, Zdozz6, Rfozz6, Uhozz6, Mkozz6, Bnozz6, Fqozz6, Jtozz6;
reg Zvozz6, Ryozz6, M0pzz6, E2pzz6, S3pzz6, L5pzz6, Z6pzz6, Dapzz6, Hdpzz6, Vfpzz6;
reg Nipzz6, Qlpzz6, Topzz6, Hrpzz6, Ztpzz6, Tvpzz6, Kxpzz6, Bzpzz6, D1qzz6, A4qzz6;
reg X6qzz6, M9qzz6, Dcqzz6, Xdqzz6, Ofqzz6, Diqzz6, Ukqzz6, Omqzz6, Foqzz6, Wpqzz6;
reg Yrqzz6, Quqzz6, Gwqzz6, Hyqzz6, W0rzz6, N3rzz6, C6rzz6, T8rzz6, Ibrzz6, Zdrzz6;
reg Ogrzz6, Fjrzz6, Blrzz6, Xmrzz6, Torzz6, Pqrzz6, Lsrzz6, Hurzz6, Bwrzz6, Sxrzz6;
reg H0szz6, Y2szz6, N5szz6, H7szz6, Y8szz6, Pbszz6, Eeszz6, Tgszz6, Ijszz6, Vlszz6;
reg Coszz6, Vqszz6, Nsszz6, Qvszz6, Tyszz6, H1tzz6, Z3tzz6, T5tzz6, H8tzz6, Zatzz6;
reg Tctzz6, Ketzz6, Dhtzz6, Sjtzz6, Oltzz6, Kntzz6, Gptzz6, Crtzz6, Ystzz6, Vutzz6;
reg Swtzz6, Pytzz6, M0uzz6, J2uzz6, F4uzz6, B6uzz6, Y7uzz6, V9uzz6, Sbuzz6, Pduzz6;
reg Ofuzz6, Jhuzz6, Hjuzz6, Vkuzz6, Qmuzz6, Iouzz6, Aquzz6, Dsuzz6, Vuuzz6, Lxuzz6;
reg D0vzz6, R1vzz6, L3vzz6, F5vzz6, V6vzz6, S8vzz6, Iavzz6, Ybvzz6, Odvzz6, Rgvzz6;
reg Ujvzz6, Mmvzz6, Bpvzz6, Fsvzz6, Jvvzz6, Byvzz6, Q0wzz6, U3wzz6, Y6wzz6, X9wzz6;
reg Bdwzz6, Agwzz6, Eiwzz6, Ikwzz6, Jnwzz6, Mqwzz6, Otwzz6, Rwwzz6, Tzwzz6, W2xzz6;
reg Y5xzz6, B9xzz6, Ecxzz6, Gfxzz6, Iixzz6, Hlxzz6, Loxzz6, Krxzz6, Ktxzz6, Lwxzz6;
reg Lyxzz6, M0yzz6, N2yzz6, O4yzz6, Q6yzz6, Q8yzz6, Vayzz6, Ycyzz6, Weyzz6, Ygyzz6;
reg Ckyzz6, Fnyzz6, Ipyzz6, Nryzz6, Ptyzz6, Xvyzz6, Uyyzz6, R1zzz6, V4zzz6, N7zzz6;
reg Cazzz6, Gdzzz6, Kgzzz6, Cjzzz6, Xkzzz6, Pmzzz6, Epzzz6, Iszzz6, Mvzzz6, Eyzzz6;
reg Zzzzz6, R10007, G40007, K70007, Oa0007, Sd0007, Rg0007, Cj0007, Nl0007, Yn0007;
reg Jq0007, Os0007, Ev0007, Ux0007, K01007, A31007, R51007, I81007, Ab1007, Rd1007;
reg Jg1007, Aj1007, Sl1007, Jo1007, Br1007, St1007, Kw1007, Bz1007, T12007, K42007;
reg C72007, T92007, Lc2007, Cf2007, Uh2007, Lk2007, Dn2007, Up2007, Ms2007, Dv2007;
reg Vx2007, M03007, E33007, V53007, N83007, Eb3007, Wd3007, Mg3007, Cj3007, Tl3007;
reg Jo3007, Ar3007, St3007, Jw3007, Bz3007, S14007, K44007, B74007, T94007, Jc4007;
reg Af4007, Rh4007, Ik4007, Zm4007, Qp4007, Hs4007, Yu4007, Px4007, G05007, X25007;
reg O55007, F85007, Wa5007, Nd5007, Eg5007, Vi5007, Ml5007, Do5007, Uq5007, Lt5007;
reg Cw5007, Sy5007, I16007, Y36007, O66007, E96007, Ub6007, Ke6007, Ah6007, Qj6007;
reg Gm6007, Xo6007, Or6007, Fu6007, Ww6007, Nz6007, E27007, V47007, M77007, Da7007;
reg Uc7007, Lf7007, Ci7007, Tk7007, Kn7007, Bq7007, Ss7007, Jv7007, Ay7007, R08007;
reg I38007, Z58007, P88007, Fb8007, Vd8007, Lg8007, Bj8007, Rl8007, Ho8007, Xq8007;
reg Nt8007, Dw8007, Uy8007, L19007, C49007, T69007, K99007, Bc9007, Se9007, Jh9007;
reg Ak9007, Rm9007, Ip9007, Zr9007, Qu9007, Hx9007, Yz9007, P2a007, G5a007, X7a007;
reg Oaa007, Fda007, Wfa007, Mia007, Cla007, Sna007, Iqa007, Ysa007, Ova007, Eya007;
reg U0b007, K3b007, A6b007, R8b007, Ibb007, Zdb007, Qgb007, Hjb007, Ylb007, Pob007;
reg Grb007, Xtb007, Owb007, Fzb007, W1c007, N4c007, E7c007, V9c007, Mcc007, Dfc007;
reg Uhc007, Lkc007, Cnc007, Tpc007, Jsc007, Zuc007, Pxc007, F0d007, V2d007, L5d007;
reg B8d007, Rad007, Hdd007, Xfd007, Oid007, Fld007, Wnd007, Nqd007, Etd007, Vvd007;
reg Myd007, D1e007, U3e007, L6e007, C9e007, Tbe007, Kee007, Bhe007, Sje007, Jme007;
reg Ape007, Rre007, Iue007, Zwe007, Qze007, G2f007, W4f007, M7f007, Caf007, Scf007;
reg Iff007, Yhf007, Okf007, Enf007, Vpf007, Nsf007, Fvf007, Xxf007, P0g007, H3g007;
reg Z5g007, R8g007, Jbg007, Beg007, Tgg007, Ljg007, Dmg007, Vog007, Nrg007, Fug007;
reg Xwg007, Pzg007, H2h007, Z4h007, R7h007, Jah007, Adh007, Rfh007, Iih007, Zkh007;
reg Qnh007, Hqh007, Ysh007, Pvh007, Gyh007, X0i007, P3i007, H6i007, Z8i007, Rbi007;
reg Jei007, Bhi007, Tji007, Lmi007, Dpi007, Vri007, Nui007, Fxi007, Xzi007, P2j007;
reg H5j007, Z7j007, Raj007, Jdj007, Bgj007, Tij007, Llj007, Coj007, Tqj007, Ktj007;
reg Bwj007, Syj007, J1k007, A4k007, R6k007, I9k007, Zbk007, Rek007, Jhk007, Bkk007;
reg Tmk007, Lpk007, Dsk007, Vuk007, Nxk007, F0l007, X2l007, P5l007, H8l007, Zal007;
reg Rdl007, Jgl007, Bjl007, Tll007, Lol007, Drl007, Vtl007, Nwl007, Ezl007, V1m007;
reg M4m007, D7m007, U9m007, Lcm007, Cfm007, Thm007, Kkm007, Bnm007, Tpm007, Lsm007;
reg Dvm007, Vxm007, N0n007, F3n007, X5n007, P8n007, Hbn007, Zdn007, Rgn007, Jjn007;
reg Bmn007, Ton007, Lrn007, Dun007, Vwn007, Nzn007, F2o007, X4o007, P7o007, Gao007;
reg Xco007, Ofo007, Fio007, Wko007, Nno007, Eqo007, Vso007, Nvo007, Fyo007, X0p007;
reg P3p007, H6p007, Z8p007, Rbp007, Jep007, Bhp007, Tjp007, Lmp007, Dpp007, Vrp007;
reg Nup007, Fxp007, Xzp007, P2q007, H5q007, Z7q007, Raq007, Jdq007, Agq007, Riq007;
reg Ilq007, Znq007, Qqq007, Htq007, Yvq007, Pyq007, G1r007, W3r007, N6r007, E9r007;
reg Vbr007, Mer007, Dhr007, Ujr007, Lmr007, Cpr007, Trr007, Kur007, Bxr007, Szr007;
reg J2s007, A5s007, R7s007, Ias007, Zcs007, Qfs007, His007, Yks007, Pns007, Fqs007;
reg Vss007, Lvs007, Bys007, R0t007, H3t007, X5t007, N8t007, Dbt007, Tdt007, Kgt007;
reg Bjt007, Slt007, Jot007, Art007, Rtt007, Iwt007, Zyt007, Q1u007, H4u007, Y6u007;
reg P9u007, Gcu007, Xeu007, Ohu007, Fku007, Wmu007, Npu007, Esu007, Vuu007, Mxu007;
reg C0v007, S2v007, I5v007, Y7v007, Oav007, Edv007, Ufv007, Kiv007, Alv007, Qnv007;
reg Hqv007, Ysv007, Pvv007, Gyv007, X0w007, O3w007, F6w007, W8w007, Nbw007, Eew007;
reg Vgw007, Mjw007, Dmw007, Uow007, Lrw007, Cuw007, Tww007, Kzw007, B2x007, S4x007;
reg J7x007, Z9x007, Pcx007, Ffx007, Vhx007, Lkx007, Bnx007, Rpx007, Hsx007, Xux007;
reg Nxx007, E0y007, V2y007, M5y007, D8y007, Uay007, Ldy007, Cgy007, Tiy007, Kly007;
reg Boy007, Sqy007, Jty007, Awy007, Ryy007, I1z007, Z3z007, Q6z007, H9z007, Ybz007;
reg Pez007, Ghz007, Wjz007, Mmz007, Cpz007, Srz007, Iuz007, Ywz007, Ozz007, E20107;
reg U40107, Y70107, Qa0107, Lc0107, De0107, Sg0107, Wj0107, An0107, Pp0107, Hs0107;
reg Cu0107, Uv0107, Yy0107, C21107, R41107, J71107, E91107, Wa1107, Ae1107, Eh1107;
reg Tj1107, Lm1107, Go1107, Yp1107, Ct1107, Gw1107, Ez1107, L12107, S32107, V62107;
reg U92107, Yc2107, Nf2107, Fi2107, Ak2107, Sl2107, Wo2107, As2107, Yu2107, Xx2107;
reg W03107, V33107, U63107, T93107, Sc3107, Rf3107, Sh3107, Sj3107, Yl3107, Fo3107;
reg Oq3107, Rt3107, Qw3107, Wy3107, C14107, H34107, N54107, T74107, Z94107, Fc4107;
reg Le4107, Rg4107, Xi4107, Dl4107, Jn4107, Pp4107, Vr4107, Bu4107, Ax4107, Xz4107;
reg U25107, L55107, I85107, Ka5107, Yc5107, Wf5107, Ui5107, Kl5107, En5107, Yo5107;
reg Oq5107, Is5107, Yt5107, Ov5107, Bx5107, Ry5107, I06107, Z16107, P36107, F56107;
reg V66107, L86107, Ba6107, Rb6107, Gd6107, Ve6107, Kg6107, Yh6107, Lj6107, Fl6107;
reg Zn6107, Br6107, Du6107, Bx6107, Vz6107, U27107, T57107, V87107, Xb7107, We7107;
reg Dh7107, Kj7107, Rl7107, Yn7107, Eq7107, Ks7107, Lu7107, Qw7107, Qz7107, Q28107;
reg Q58107, Q88107, Gttf07, Gwtf07, Eztf07, G2uf07, G5uf07, J8uf07, Mbuf07, Peuf07;
reg Ahuf07, Xjuf07, Umuf07, Fpuf07, Csuf07, Zuuf07, Kxuf07, H0vf07, E3vf07, B6vf07;
reg I8vf07, Mbvf07, Bevf07, Tgvf07, Oivf07, Gkvf07, Knvf07, Oqvf07, Dtvf07, Vvvf07;
reg Qxvf07, Izvf07, M2wf07, Q5wf07, F8wf07, Xawf07, Scwf07, Kewf07, Ohwf07, Skwf07;
reg Wnwf07, Lqwf07, Ltwf07, Jwwf07, Hzwf07, D2xf07, D5xf07, A8xf07, Uaxf07, Udxf07;
reg Ngxf07, Wixf07, Xkxf07, Unxf07, Bqxf07, Hsxf07, Nuxf07, Twxf07, Zyxf07, F1yf07;
reg K3yf07, P5yf07, U7yf07, Xayf07, Ndyf07, Dgyf07, Tiyf07, Jlyf07, Znyf07, Pqyf07;
reg Ftyf07, Tvyf07, Xyyf07, B2zf07, E5zf07, I8zf07, Nazf07, Sczf07, Tfzf07, Thzf07;
reg Vjzf07, Lmzf07, Fozf07, Zqzf07, Ptzf07, Owzf07, Byzf07, Yzzf07, M10g07, C30g07;
reg S40g07, H60g07, W70g07, L90g07, Ab0g07, Pc0g07, Ee0g07, Tf0g07, Zg0g07, Fi0g07;
reg Lj0g07, Rk0g07, Om0g07, Lo0g07, Iq0g07, Fs0g07, Cu0g07, Zv0g07, Wx0g07, Uz0g07;
reg S11g07, N31g07, F51g07, G71g07, V81g07, Ka1g07, Zb1g07, Od1g07, Df1g07, Pg1g07;
reg Qi1g07, Rk1g07, Mm1g07, Ap1g07, Ds1g07, Gv1g07, Uw1g07, Iy1g07, Xz1g07, L12g07;
reg C42g07, T62g07, M92g07, Fc2g07, Ye2g07, Rh2g07, Lk2g07, Fn2g07, Zp2g07, Ts2g07;
reg Nv2g07, Hy2g07, B13g07, V33g07, P63g07, J93g07, Dc3g07, Xe3g07, Rh3g07, Lk3g07;
reg Fn3g07, Zp3g07, Ts3g07, Nv3g07, Hy3g07, B14g07, V34g07, O64g07, S84g07, Ra4g07;
reg Tc4g07, Af4g07, Yh4g07, Xk4g07, Vn4g07, Tq4g07, Rt4g07, Pw4g07, Oz4g07, N25g07;
reg M55g07, L85g07, Kb5g07, Ie5g07, Gh5g07, Bk5g07, Ym5g07, Xp5g07, Ws5g07, Vv5g07;
reg Uy5g07, T16g07, W46g07, Z76g07, Xa6g07, Ae6g07, Yg6g07, Wj6g07, Xm6g07, Yp6g07;
reg Zs6g07, Gv6g07, Ky6g07, T07g07, H37g07, P57g07, R87g07, Tb7g07, Ve7g07, Xh7g07;
reg Ak7g07, Dm7g07, Go7g07, Jq7g07, Ss7g07, Bv7g07, Lx7g07, Vz7g07, V18g07, E48g07;
reg N68g07, W88g07, Fb8g07, Kd8g07, Pf8g07, Uh8g07, Zj8g07, Em8g07, Jo8g07, Oq8g07;
reg Ts8g07, Yu8g07, Dx8g07, Iz8g07, N19g07, S39g07, W59g07, A89g07, Ea9g07, Ic9g07;
reg Me9g07, Qg9g07, Ui9g07, Yk9g07, Hn9g07, Qp9g07, Sr9g07, Ut9g07, Wv9g07, Zx9g07;
reg C0ag07, F2ag07, H4ag07, J6ag07, L8ag07, Paag07, Tcag07, Xeag07, Bhag07, Gjag07;
reg Llag07, Qnag07, Vpag07, Asag07, Fuag07, Kwag07, Nyag07, Q0bg07, T2bg07, W4bg07;
reg Z6bg07, C9bg07, Fbbg07, Idbg07, Lfbg07, Phbg07, Tjbg07, Ylbg07, Dobg07, Iqbg07;
reg Nsbg07, Subg07, Xwbg07, Czbg07, H1cg07, M3cg07, R5cg07, W7cg07, Aacg07, Eccg07;
reg Iecg07, Mgcg07, Qicg07, Ukcg07, Ymcg07, Cpcg07, Grcg07, Ktcg07, Ovcg07, Nxcg07;
reg Mzcg07, P1dg07, S3dg07, V5dg07, Y7dg07, Badg07, Ecdg07, Hedg07, Kgdg07, Nidg07;
reg Qkdg07, Tmdg07, Wodg07, Zqdg07, Ctdg07, Fvdg07, Ixdg07, Lzdg07, O1eg07, R3eg07;
reg U5eg07, X7eg07, Aaeg07, Dceg07, Geeg07, Jgeg07, Mieg07, Pkeg07, Smeg07, Qpeg07;
reg Rseg07, Vueg07, Xweg07, Czeg07, H1fg07, M3fg07, R5fg07, W7fg07, Bafg07, Gcfg07;
reg Lefg07, Qgfg07, Vifg07, Alfg07, Enfg07, Ipfg07, Mrfg07, Qtfg07, Uvfg07, Yxfg07;
reg C0gg07, G2gg07, K4gg07, O6gg07, S8gg07, Pagg07, Qcgg07, Oegg07, Tggg07, Bjgg07;
reg Klgg07, Ongg07, Cqgg07, Jsgg07, Qugg07, Xwgg07, Ezgg07, B2hg07, Y4hg07, F7hg07;
reg M9hg07, Pbhg07, Sdhg07, Vfhg07, Rhhg07, Njhg07, Jlhg07, Fnhg07, Bphg07, Xqhg07;
reg Tshg07, Puhg07, Mwhg07, Jyhg07, G0ig07, D2ig07, A4ig07, X5ig07, U7ig07, R9ig07;
reg Obig07, Ldig07, Ifig07, Fhig07, Cjig07, Zkig07, Wmig07, Toig07, Qqig07, Nsig07;
reg Kuig07, Hwig07, Myig07, R0jg07, W2jg07, B5jg07, G7jg07, L9jg07, Qbjg07, Vdjg07;
reg Agjg07, Fijg07, Kkjg07, Omjg07, Sojg07, Wqjg07, Atjg07, Evjg07, Ixjg07, Mzjg07;
reg Q1kg07, U3kg07, Y5kg07, C8kg07, Cakg07, Hckg07, Mekg07, Rgkg07, Wikg07, Blkg07;
reg Gnkg07, Lpkg07, Qrkg07, Vtkg07, Awkg07, Fykg07, J0lg07, N2lg07, R4lg07, V6lg07;
reg Z8lg07, Dblg07, Hdlg07, Lflg07, Phlg07, Tjlg07, Xllg07, Bolg07, Qplg07, Hrlg07;
reg Yslg07, Zulg07, Axlg07, Ezlg07, I1mg07, H3mg07, I5mg07, J7mg07, F9mg07, Lbmg07;
reg Rdmg07, Xfmg07, Dimg07, Hkmg07, Ylmg07, Pnmg07, Epmg07, Vqmg07, Msmg07, Dumg07;
reg Vvmg07, Nxmg07, Fzmg07, X0ng07, P2ng07, H4ng07, Z5ng07, R7ng07, J9ng07, Bbng07;
reg Tcng07, Leng07, Dgng07, Vhng07, Njng07, Flng07, Xmng07, Pong07, Hqng07, Zrng07;
reg Rtng07, Jvng07, Axng07, Ryng07, I0og07, Z1og07, Q3og07, H5og07, Y6og07, P8og07;
reg Gaog07, Ncog07, Eeog07, Vfog07, Mhog07, Djog07, Ukog07, Lmog07, Coog07, Tpog07;
reg Krog07, Btog07, Tuog07, Lwog07, Dyog07, Vzog07, N1pg07, F3pg07, X4pg07, P6pg07;
reg H8pg07, Z9pg07, Rbpg07, Jdpg07, Bfpg07, Tgpg07, Lipg07, Dkpg07, Vlpg07, Nnpg07;
reg Fppg07, Xqpg07, Pspg07, Supg07, Xwpg07, Azpg07, C1qg07, G3qg07, J5qg07, N7qg07;
reg T9qg07, Ubqg07, Wdqg07, Yfqg07, Biqg07, Dkqg07, Gmqg07, Joqg07, Mqqg07, Psqg07;
reg Suqg07, Vwqg07, Yyqg07, B1rg07, E3rg07, H5rg07, K7rg07, N9rg07, Qbrg07, Tdrg07;
reg Wfrg07, Yhrg07, Akrg07, Cmrg07, Eorg07, Gqrg07, Isrg07, Kurg07, Mwrg07, Oyrg07;
reg T0sg07, Y2sg07, D5sg07, I7sg07, N9sg07, Sbsg07, Xdsg07, Cgsg07, Hisg07, Mksg07;
reg Rmsg07, Vosg07, Zqsg07, Dtsg07, Hvsg07, Lxsg07, Pzsg07, T1tg07, X3tg07, B6tg07;
reg F8tg07, Jatg07, Kctg07, Letg07, Kgtg07, Jitg07, Iktg07, Hmtg07, Hotg07, Hqtg07;
reg Hstg07, Hutg07, Hwtg07, Hytg07, G0ug07, F2ug07, E4ug07, J6ug07, O8ug07, Taug07;
reg Ycug07, Dfug07, Ihug07, Njug07, Slug07, Xnug07, Cqug07, Hsug07, Luug07, Pwug07;
reg Tyug07, X0vg07, B3vg07, F5vg07, J7vg07, N9vg07, Rbvg07, Vdvg07, Zfvg07, Aivg07;
reg Bkvg07, Cmvg07, Dovg07, Eqvg07, Fsvg07, Guvg07, Hwvg07, Iyvg07, J0wg07, K2wg07;
reg L4wg07, M6wg07, N8wg07, Nawg07, Ocwg07, Pewg07, Qgwg07, Riwg07, Skwg07, Tmwg07;
reg Towg07, Tqwg07, Tswg07, Tuwg07, Twwg07, Tywg07, T0xg07, U2xg07, S5xg07, Q8xg07;
reg Vaxg07, Adxg07, Ffxg07, Khxg07, Pjxg07, Ulxg07, Znxg07, Eqxg07, Jsxg07, Ouxg07;
reg Twxg07, Xyxg07, B1yg07, F3yg07, J5yg07, N7yg07, R9yg07, Vbyg07, Zdyg07, Dgyg07;
reg Hiyg07, Lkyg07, Nmyg07, Poyg07, Rqyg07, Tsyg07, Vuyg07, Xwyg07, Zyyg07, B1zg07;
reg E3zg07, H5zg07, K7zg07, N9zg07, Qbzg07, Tdzg07, Wfzg07, Zhzg07, Ckzg07, Fmzg07;
reg Iozg07, Lqzg07, Oszg07, Ruzg07, Uwzg07, Xyzg07, A10h07, D30h07, G50h07, J70h07;
reg L90h07, Nb0h07, Pd0h07, Rf0h07, Th0h07, Vj0h07, Xl0h07, Zn0h07, Bq0h07, Ds0h07;
reg Fu0h07, Hw0h07, Iy0h07, J01h07, K21h07, L41h07, M61h07, N81h07, Oa1h07, Hd1h07;
reg Ag1h07, Ni1h07, Ml1h07, Lo1h07, Zq1h07, St1h07, Lw1h07, Kz1h07, J22h07, F52h07;
reg C82h07, R92h07, Fb2h07, Xc2h07, Ne2h07, Dg2h07, Th2h07, Ij2h07, Xk2h07, Mm2h07;
reg Bo2h07, Qp2h07, Fr2h07, Vs2h07, Lu2h07, Bw2h07, Rx2h07, Hz2h07, X03h07, N23h07;
reg D43h07, V53h07, J73h07, B93h07, Ra3h07, Hc3h07, Xd3h07, Mf3h07, Bh3h07, Qi3h07;
reg Fk3h07, Ul3h07, Jn3h07, Zo3h07, Pq3h07, Fs3h07, Vt3h07, Lv3h07, Bx3h07, Ry3h07;
reg H04h07, Z14h07, M34h07, A54h07, Q64h07, G84h07, W94h07, Lb4h07, Ad4h07, Pe4h07;
reg Eg4h07, Th4h07, Ij4h07, Yk4h07, Om4h07, Eo4h07, Up4h07, Kr4h07, At4h07, Qu4h07;
reg Gw4h07, Ux4h07, Kz4h07, A15h07, P25h07, E45h07, T55h07, I75h07, X85h07, Ma5h07;
reg Cc5h07, Sd5h07, If5h07, Yg5h07, Oi5h07, Ek5h07, Ul5h07, In5h07, Ap5h07, Qq5h07;
reg Gs5h07, Wt5h07, Lv5h07, Ax5h07, Py5h07, E06h07, T16h07, I36h07, Y46h07, O66h07;
reg E86h07, U96h07, Kb6h07, Ad6h07, Qe6h07, Gg6h07, Yh6h07, Mj6h07, El6h07, Um6h07;
reg Ko6h07, Aq6h07, Pr6h07, Et6h07, Tu6h07, Iw6h07, Xx6h07, Mz6h07, C17h07, S27h07;
reg I47h07, Y57h07, O77h07, E97h07, Ua7h07, Kc7h07, Ce7h07, Qf7h07, Gh7h07, Wi7h07;
reg Mk7h07, Bm7h07, Qn7h07, Fp7h07, Uq7h07, Js7h07, Yt7h07, Ov7h07, Ex7h07, Uy7h07;
reg K08h07, A28h07, Q38h07, G58h07, W68h07, O88h07, Ca8h07, Ub8h07, Kd8h07, Af8h07;
reg Qg8h07, Fi8h07, Uj8h07, Jl8h07, Ym8h07, No8h07, Cq8h07, Sr8h07, It8h07, Yu8h07;
reg Ow8h07, Ey8h07, Uz8h07, K19h07, A39h07, S49h07, J69h07, A89h07, Q99h07, Gb9h07;
reg Wc9h07, Me9h07, Cg9h07, Sh9h07, Ij9h07, Yk9h07, Pm9h07, Go9h07, Xp9h07, Or9h07;
reg Ft9h07, Wu9h07, Xw9h07, Zy9h07, B1ah07, D3ah07, J5ah07, P7ah07, R9ah07, Tbah07;
reg Vdah07, Bgah07, Hiah07, Jkah07, Lmah07, Noah07, Oqah07, Msah07, Luah07, Kwah07;
reg Jyah07, I0bh07, H2bh07, G4bh07, F6bh07, E8bh07, Dabh07, Ccbh07, Bebh07, Agbh07;
reg Zhbh07, Yjbh07, Xlbh07, Wnbh07, Vpbh07, Urbh07, Ttbh07, Svbh07, Rxbh07, Qzbh07;
reg O1ch07, M3ch07, K5ch07, I7ch07, G9ch07, Ebch07, Cdch07, Afch07, Chch07, Fjch07;
reg Ilch07, Lnch07, Opch07, Rrch07, Utch07, Xvch07, Aych07, D0dh07, G2dh07, J4dh07;
reg M6dh07, P8dh07, Sadh07, Vcdh07, Yedh07, Bhdh07, Ejdh07, Hldh07, Kndh07, Npdh07;
reg Qrdh07, Stdh07, Uvdh07, Wxdh07, Yzdh07, A2eh07, C4eh07, E6eh07, G8eh07, Daeh07;
reg Bceh07, Zdeh07, Xfeh07, Vheh07, Tjeh07, Rleh07, Pneh07, Npeh07, Lreh07, Jteh07;
reg Hveh07, Fxeh07, Dzeh07, A1fh07, X2fh07, U4fh07, R6fh07, O8fh07, Lafh07, Icfh07;
reg Fefh07, Kgfh07, Qifh07, Wkfh07, Cnfh07, Apfh07, Yqfh07, Wsfh07, Yufh07, Axfh07;
reg Czfh07, H1gh07, N3gh07, T5gh07, Z7gh07, Bagh07, Ecgh07, Hegh07, Kggh07, Nigh07;
reg Qkgh07, Tmgh07, Wogh07, Zqgh07, Ctgh07, Fvgh07, Ixgh07, Lzgh07, O1hh07, R3hh07;
reg U5hh07, X7hh07, Aahh07, Dchh07, Gehh07, Jghh07, Mihh07, Pkhh07, Rmhh07, Tohh07;
reg Vqhh07, Xshh07, Zuhh07, Bxhh07, Dzhh07, F1ih07, H3ih07, J5ih07, L7ih07, N9ih07;
reg Pbih07, Rdih07, Tfih07, Vhih07, Yjih07, Bmih07, Eoih07, Hqih07, Ksih07, Nuih07;
reg Qwih07, Tyih07, W0jh07, Z2jh07, C5jh07, F7jh07, I9jh07, Lbjh07, Odjh07, Rfjh07;
reg Uhjh07, Xjjh07, Amjh07, Dojh07, Gqjh07, Jsjh07, Lujh07, Qwjh07, Wyjh07, C1kh07;
reg I3kh07, Q5kh07, C8kh07, Oakh07, Adkh07, Mfkh07, Uhkh07, Ckkh07, Ylkh07, Nnkh07;
reg Fqkh07, Xskh07, Pvkh07, Hykh07, Z0lh07, R3lh07, J6lh07, B9lh07, Tblh07, Kelh07;
reg Bhlh07, Sjlh07, Jmlh07, Aplh07, Rrlh07, Iulh07, Zwlh07, Qzlh07, Z1mh07, I4mh07;
reg Q6mh07, Y8mh07, Gbmh07, Pdmh07, Yfmh07, Rhmh07, Wjmh07, Bmmh07, Gomh07, Lqmh07;
reg Qsmh07, Vumh07, Dxmh07, Lzmh07, T1nh07, B4nh07, J6nh07, R8nh07, Zanh07, Idnh07;
reg Rfnh07, Ainh07, Jknh07, Smnh07, Bpnh07, Jrnh07, Etnh07, Zunh07, Uwnh07, Pynh07;
reg K0oh07, F2oh07, U3oh07, P5oh07, G7oh07, B9oh07, Kboh07, Idoh07, Gfoh07, Ehoh07;
reg Cjoh07, Aloh07, Ymoh07, Wooh07, Uqoh07, Ssoh07, Ruoh07, Pwoh07, Wyoh07, W0ph07;
reg U2ph07, R4ph07, T6ph07, W8ph07, Bbph07, Gdph07, Qfph07, Aiph07, Kkph07, Emph07;
reg Joph07, Hqph07, Lsph07, Vuph07, Ixph07, Pzph07, R1qh07, Z3qh07, F6qh07, D8qh07;
reg Oaqh07, Scqh07, Zeqh07, Dhqh07, Ejqh07, Zkqh07, Fnqh07, Woqh07, Uqqh07, Vsqh07;
reg Nuqh07, Lwqh07, Kyqh07, J0rh07, I2rh07, H4rh07, G6rh07, F8rh07, Earh07, Dcrh07;
reg Cerh07, Bgrh07, Airh07, Zjrh07, Ylrh07, Xnrh07, Wprh07, Vrrh07, Gxps07, Fzps07;
reg E1qs07, D3qs07, C5qs07, B7qs07, A9qs07, Zaqs07, Ycqs07, Xeqs07, Wgqs07, Viqs07;
reg Ukqs07, Tmqs07, Soqs07, Rqqs07, Qsqs07, Puqs07, Owqs07, Nyqs07, M0rs07, L2rs07;
reg K4rs07, I6rs07, G8rs07, Ears07, Ccrs07, Aers07, Yfrs07, Whrs07, Ujrs07, Dmrs07;
reg Mors07, Vqrs07, Etrs07, Nvrs07, Wxrs07, F0ss07, O2ss07, X4ss07, L7ss07, G9ss07;
reg Bbss07, Wcss07, Tess07, Ngss07, Hiss07, Bkss07, Cmss07, Aoss07, Ypss07, Vrss07;
reg Stss07, Pvss07, Mxss07, Kzss07, I1ts07, G3ts07, C5ts07, P7ts07, Cats07, Fcts07;
reg Dets07, Bgts07, Zhts07, Xjts07, Vlts07, Tnts07, Rpts07, Prts07, Ntts07, Mvts07;
reg Lxts07, Kzts07, H1us07, E3us07, D5us07, F7us07, C9us07, Ebus07, Fdus07, Gfus07;
reg Thus07, Mkus07, Fnus07, Lous07, Bqus07, Prus07, Ntus07, Mvus07, Kxus07, Xzus07;
reg Q2vs07, J5vs07, H7vs07, F9vs07, Dbvs07, Bdvs07, Zevs07, Xgvs07, Vivs07, Tkvs07;
reg Rmvs07, Povs07, Nqvs07, Lsvs07, Juvs07, Hwvs07, Uyvs07, N1ws07, G4ws07, X5ws07;
reg O7ws07, F9ws07, Waws07, Ncws07, Eews07, Wfws07, Yhws07, Qjws07, Ilws07, Lnws07;
reg Hpws07, Drws07, Atws07, Xuws07, Uwws07, Tyws07, S0xs07, R2xs07, Q4xs07, P6xs07;
reg O8xs07, Naxs07, Mcxs07, Lexs07, Kgxs07, Jixs07, Ikxs07, Hmxs07, Goxs07, Fqxs07;
reg Esxs07, Duxs07, Cwxs07, Byxs07, A0ys07, Z1ys07, Y3ys07, V6ys07, Y9ys07, Bdys07;
reg Egys07, Ijys07, Mmys07, Qpys07, Usys07, Yvys07, Czys07, G2zs07, D5zs07, M7zs07;
reg W9zs07, Gczs07, Qezs07, Ahzs07, Kjzs07, Ulzs07, Eozs07, Oqzs07, Yszs07, Hvzs07;
reg Rxzs07, B00t07, L20t07, V40t07, F70t07, O90t07, Lc0t07, Ve0t07, Sh0t07, Dk0t07;
reg Gm0t07, Lo0t07, Kr0t07, Ju0t07, Ix0t07, L01t07, M31t07, J61t07, G91t07, Lb1t07;
reg Qd1t07, Tg1t07, Qi1t07, Sk1t07, Um1t07, Wo1t07, Cr1t07, Jt1t07, Pv1t07, Nx1t07;
reg Lz1t07, N12t07, P32t07, R52t07, Z72t07, Ba2t07, Ac2t07, Ge2t07, Fg2t07, Li2t07;
reg Tk2t07, Vm2t07, Xo2t07, Er2t07, It2t07, Pv2t07, Ox2t07, Qz2t07, J23t07, K33t07;
reg J43t07, K63t07, Q83t07, Pa3t07, Pc3t07, Qe3t07, Ug3t07, Ni3t07, Kk3t07, Jm3t07;
reg Io3t07, Hq3t07, Gs3t07, Fu3t07, Ew3t07, Dy3t07, C04t07, H24t07, Q44t07, Y64t07;
reg V94t07, Sc4t07, Pf4t07, Mi4t07, Ik4t07, Zn4t07, Qr4t07, Hv4t07, Vy4t07, N25t07;
reg F65t07, X95t07, Pd5t07, Hh5t07, Tk5t07, Fo5t07, Rr5t07, Dv5t07, Py5t07, B26t07;
reg N56t07, Z86t07, Lc6t07, Xf6t07, Jj6t07, Vm6t07, Hq6t07, Tt6t07, Fx6t07, R07t07;
reg D47t07, P77t07, Bb7t07, Ne7t07, Zh7t07, Ll7t07, Xo7t07, Js7t07, Uv7t07, Gz7t07;
reg S28t07, E68t07, P98t07, Ad8t07, Lg8t07, Tj8t07, Gn8t07, Tq8t07, Gu8t07, Tx8t07;
reg K19t07, B59t07, S89t07, Gc9t07, Yf9t07, Qj9t07, In9t07, Ar9t07, Su9t07, Ey9t07;
reg Q1at07, C5at07, O8at07, Acat07, Mfat07, Yiat07, Kmat07, Wpat07, Itat07, Uwat07;
reg G0bt07, S3bt07, E7bt07, Qabt07, Cebt07, Ohbt07, Albt07, Mobt07, Yrbt07, Kvbt07;
reg Wybt07, I2ct07, U5ct07, F9ct07, Rcct07, Dgct07, Pjct07, Anct07, Lqct07, Wtct07;
reg Exct07, R0dt07, E4dt07, R7dt07, Ebdt07, Vedt07, Midt07, Dmdt07, Rpdt07, Jtdt07;
reg Bxdt07, T0et07, L4et07, D8et07, Pbet07, Bfet07, Niet07, Zlet07, Lpet07, Xset07;
reg Jwet07, Vzet07, H3ft07, T6ft07, Faft07, Rdft07, Dhft07, Pkft07, Boft07, Nrft07;
reg Zuft07, Lyft07, X1gt07, J5gt07, V8gt07, Hcgt07, Tfgt07, Fjgt07, Qmgt07, Cqgt07;
reg Otgt07, Axgt07, L0ht07, W3ht07, H7ht07, Paht07, Ceht07, Phht07, Clht07, Poht07;
reg Gsht07, Xvht07, Ozht07, C3it07, U6it07, Mait07, Eeit07, Whit07, Olit07, Apit07;
reg Msit07, Yvit07, Kzit07, W2jt07, I6jt07, U9jt07, Gdjt07, Sgjt07, Ekjt07, Qnjt07;
reg Crjt07, Oujt07, Ayjt07, M1kt07, Y4kt07, K8kt07, Wbkt07, Ifkt07, Uikt07, Gmkt07;
reg Spkt07, Etkt07, Qwkt07, B0lt07, N3lt07, Z6lt07, Lalt07, Wdlt07, Hhlt07, Sklt07;
reg Aolt07, Nrlt07, Avlt07, Nylt07, A2mt07, U3mt07, V5mt07, Q7mt07, Pamt07, Scmt07;
reg Uemt07, Rhmt07, Ilmt07, Zomt07, Qsmt07, Ewmt07, Wzmt07, O3nt07, G7nt07, Yant07;
reg Qent07, Cint07, Olnt07, Apnt07, Msnt07, Yvnt07, Kznt07, W2ot07, I6ot07, U9ot07;
reg Gdot07, Sgot07, Ekot07, Qnot07, Crot07, Ouot07, Ayot07, M1pt07, Y4pt07, K8pt07;
reg Wbpt07, Ifpt07, Uipt07, Gmpt07, Sppt07, Dtpt07, Pwpt07, B0qt07, N3qt07, Y6qt07;
reg Jaqt07, Udqt07, Chqt07, Pkqt07, Coqt07, Prqt07, Cvqt07, Zxqt07, Q1rt07, H5rt07;
reg Y8rt07, Mcrt07, Egrt07, Wjrt07, Onrt07, Grrt07, Yurt07, Kyrt07, W1st07, I5st07;
reg U8st07, Gcst07, Sfst07, Ejst07, Qmst07, Cqst07, Otst07, Axst07, M0tt07, Y3tt07;
reg K7tt07, Watt07, Iett07, Uhtt07, Gltt07, Sott07, Estt07, Qvtt07, Cztt07, O2ut07;
reg A6ut07, L9ut07, Xcut07, Jgut07, Vjut07, Gnut07, Rqut07, Cuut07, Kxut07, X0vt07;
reg K4vt07, X7vt07, Kbvt07, Hevt07, Yhvt07, Plvt07, Gpvt07, Usvt07, Mwvt07, E0wt07;
reg W3wt07, O7wt07, Gbwt07, Sewt07, Eiwt07, Qlwt07, Cpwt07, Oswt07, Awwt07, Mzwt07;
reg Y2xt07, K6xt07, W9xt07, Idxt07, Ugxt07, Gkxt07, Snxt07, Erxt07, Quxt07, Cyxt07;
reg O1yt07, A5yt07, M8yt07, Ybyt07, Kfyt07, Wiyt07, Imyt07, Tpyt07, Ftyt07, Rwyt07;
reg D0zt07, O3zt07, Z6zt07, Kazt07, Sdzt07, Fhzt07, Skzt07, Fozt07, Crzt07, Tuzt07;
reg Kyzt07, B20u07, P50u07, H90u07, Zc0u07, Rg0u07, Jk0u07, Bo0u07, Nr0u07, Zu0u07;
reg Ly0u07, X11u07, J51u07, V81u07, Hc1u07, Pf1u07, Cj1u07, Pm1u07, Cq1u07, Ot1u07;
reg Ax1u07, M02u07, Y32u07, K72u07, Wa2u07, Ie2u07, Uh2u07, Fl2u07, Ro2u07, Ds2u07;
reg Pv2u07, Az2u07, L23u07, W53u07, I93u07, Uc3u07, Gg3u07, Sj3u07, En3u07, Qq3u07;
reg Cu3u07, Ox3u07, Oz3u07, B34u07, O64u07, Ba4u07, Od4u07, Bh4u07, Ok4u07, Bo4u07;
reg Or4u07, Lt4u07, Av4u07, Pw4u07, Ey4u07, Tz4u07, I15u07, X25u07, M45u07, B65u07;
reg H85u07, Na5u07, Uc5u07, Ef5u07, Ii5u07, Pk5u07, Zm5u07, Xp5u07, Bt5u07, Iv5u07;
reg Sx5u07, W06u07, D36u07, I66u07, N96u07, Tc6u07, Zf6u07, Fj6u07, Lm6u07, Rp6u07;
reg Xs6u07, Dw6u07, Jz6u07, P27u07, V57u07, B97u07, Fc7u07, Fe7u07, Qg7u07, Qi7u07;
reg Bl7u07, Bn7u07, Mp7u07, Mr7u07, Xt7u07, Xv7u07, Iy7u07, I08u07, T28u07, T48u07;
reg E78u07, E98u07, Pb8u07, Pd8u07, Ag8u07, Bi8u07, Nk8u07, Om8u07, Ap8u07, Br8u07;
reg Nt8u07, Ov8u07, Ay8u07, B09u07, N29u07, O49u07, A79u07, B99u07, Nb9u07, Od9u07;
reg Ag9u07, Bi9u07, Nk9u07, Om9u07, Ap9u07, Br9u07, Nt9u07, Ov9u07, Ay9u07, B0au07;
reg N2au07, O4au07, A7au07, B9au07, Nbau07, Odau07, Agau07, Biau07, Nkau07, Omau07;
reg Apau07, Brau07, Ntau07, Ovau07, Ayau07, B0bu07, N2bu07, O4bu07, A7bu07, A9bu07;
reg Zabu07, Ldbu07, Sfbu07, Rhbu07, Dkbu07, Kmbu07, Jobu07, Vqbu07, Ctbu07, Bvbu07;
reg Nxbu07, Uzbu07, T1cu07, F4cu07, M6cu07, L8cu07, Xacu07, Edcu07, Dfcu07, Phcu07;
reg Ojcu07, Amcu07, Zncu07, Lqcu07, Lscu07, Yucu07, Ywcu07, Lzcu07, L1du07, Y3du07;
reg Y5du07, L8du07, Ladu07, Ycdu07, Yedu07, Lhdu07, Ljdu07, Yldu07, Yndu07, Lqdu07;
reg Lsdu07, Yudu07, Ywdu07, Lzdu07, L1eu07, Y3eu07, Y5eu07, L8eu07, Laeu07, Yceu07;
reg Yeeu07, Lheu07, Ljeu07, Yleu07, Yneu07, Lqeu07, Lseu07, Yueu07, Yweu07, Lzeu07;
reg L1fu07, Y3fu07, Y5fu07, L8fu07, Lafu07, Ycfu07, Lffu07, Mhfu07, Ljfu07, Rlfu07;
reg Rnfu07, Zpfu07, Bsfu07, Cufu07, Dwfu07, Eyfu07, D0gu07, D2gu07, L4gu07, N6gu07;
reg O9gu07, Pbgu07, Ndgu07, Ofgu07, Uhgu07, Akgu07, Imgu07, Qogu07, Uqgu07, Xsgu07;
reg Wugu07, Vwgu07, Azgu07, D1hu07, E3hu07, H5hu07, K7hu07, N9hu07, Rbhu07, Vdhu07;
reg Zfhu07, Dihu07, Hkhu07, Lmhu07, Pohu07, Tqhu07, Xshu07, Bvhu07, Fxhu07, Jzhu07;
reg N1iu07, R3iu07, V5iu07, Z7iu07, Daiu07, Hciu07, Leiu07, Pgiu07, Tiiu07, Xkiu07;
reg Fniu07, Npiu07, Vriu07, Ytiu07, Gwiu07, Oyiu07, W0ju07, E3ju07, M5ju07, U7ju07;
reg Caju07, Kcju07, Seju07, Ahju07, Ijju07, Qlju07, Ynju07, Gqju07, Osju07, Wuju07;
reg Exju07, Mzju07, T1ku07, A4ku07, J6ku07, A9ku07, Ibku07, Gdku07, Afku07, Zgku07;
reg Xiku07, Vkku07, Tmku07, Roku07, Pqku07, Nsku07, Luku07, Jwku07, Hyku07, G0lu07;
reg F2lu07, E4lu07, D6lu07, C8lu07, Ualu07, Qclu07, Pelu07, Qglu07, Qilu07, Tklu07;
reg Vmlu07, Hqlu07, Stlu07, Exlu07, P0mu07, B4mu07, M7mu07, Yamu07, Jemu07, Vhmu07;
reg Glmu07, Somu07, Dsmu07, Pvmu07, Azmu07, M2nu07, X5nu07, U7nu07, W9nu07, Mbnu07;
reg Bdnu07, Qenu07, Fgnu07, Uhnu07, Jjnu07, Yknu07, Nmnu07, Conu07, Frnu07, Wtnu07;
reg Ee9917, Ng9917, Sj9917, Jm9917, Mp9917, Vr9917, Av9917, Ix9917, Zz9917, I2a917;
reg Z4a917, C8a917, Laa917, Hda917, Dga917, Zia917, Vla917, Roa917, Nra917, Mta917;
reg Mva917, Rxa917, Vza917, Y1b917, W3b917, X6b917, A9b917, Dbb917, Gdb917, Jfb917;
reg Mhb917, Pjb917, Slb917, Vnb917, Ypb917, Bsb917, Fub917, Jwb917, Nyb917, R0c917;
reg V2c917, Z4c917, D7c917, H9c917, Lbc917, Pdc917, Tfc917, Xhc917, Bkc917, Slc917;
reg Rnc917, Mpc917, Vrc917, Muc917, Uwc917, Vyc917, N1d917, C4d917, R6d917, G9d917;
reg Vbd917, Ydd917, Dgd917, Nid917, Rkd917, Wmd917, Gpd917, Krd917, Rtd917, Wvd917;
reg Gyd917, K0e917, R2e917, W4e917, V7e917, Uae917, Sde917, Qge917, Pje917, Ome917;
reg Yoe917, Cre917, Jte917, Ove917, Yxe917, C0f917, H2f917, G5f917, F8f917, Ebf917;
reg Def917, Chf917, Bkf917, Zmf917, Wof917, Vrf917, Uuf917, Txf917, S0g917, R3g917;
reg Q6g917, P9g917, Ocg917, Nfg917, Mig917, Llg917, Kog917, Jrg917, Iug917, Hxg917;
reg F0h917, D3h917, C6h917, B9h917, Ach917, Zeh917, Yhh917, Xkh917, Wnh917, Vqh917;
reg Uth917, Twh917, Szh917, R2i917, Q5i917, P8i917, Obi917, Nei917, Mhi917, Lki917;
reg Kni917, Jqi917, Iti917, Hwi917, Gzi917, F2j917, E5j917, D8j917, Naj917, Rcj917;
reg Qfj917, Pij917, Olj917, Noj917, Lrj917, Qtj917, Vvj917, Ayj917, F0k917, G2k917;
reg J4k917, M6k917, J8k917, Bck917, Nfk917, Fjk917, Rmk917, Jqk917, Vtk917, Nxk917;
reg Z0l917, R4l917, D8l917, Vbl917, Hfl917, Zil917, Lml917, Dql917, Ptl917, Svl917;
reg Yyl917, P0m917, F2m917, V3m917, L5m917, B7m917, R8m917, Ham917, Xbm917, Ndm917;
reg Nfm917, Phm917, Ikm917, Emm917, Hom917, Lqm917, Psm917, Tum917, Xwm917, Bzm917;
reg F1n917, J3n917, O5n917, T7n917, Y9n917, Dcn917, Ien917, Ngn917, Sin917, Xkn917;
reg Ann917, Dpn917, Ern917, Btn917, Nwn917, Zzn917, L3o917, X6o917, Jao917, Vdo917;
reg Hho917, Tko917, Vmo917, Woo917, Xqo917, Yso917, Zuo917, Axo917, Bzo917, C1p917;
reg D3p917, E5p917, F7p917, H9p917, Nbp917, Udp917, Bgp917, Iip917, Pkp917, Dnp917;
reg Spp917, Bsp917, Kup917, Twp917, Czp917, L1q917, U3q917, D6q917, M8q917, Vaq917;
reg Edq917, Nfq917, Whq917, Fkq917, Omq917, Xoq917, Grq917, Ptq917, Yvq917, Hyq917;
reg Q0r917, Z2r917, I5r917, Q7r917, Y9r917, Gcr917, Oer917, Wgr917, Ejr917, Mlr917;
reg Unr917, Cqr917, Esr917, Gur917, Iwr917, Kyr917, M0s917, O2s917, Q4s917, S6s917;
reg U8s917, Was917, Ycs917, Afs917, Chs917, Ejs917, Gls917, Ins917, Lps917, Krs917;
reg Ats917, Tus917, Qws917, Nys917, K0t917, G2t917, C4t917, Y5t917, U7t917, Q9t917;
reg Mbt917, Idt917, Fft917, Cht917, Zit917, Vkt917, Tmt917, Ipt917, Xrt917, Qtt917;
reg Bwt917, Myt917, K0u917, X2u917, N5u917, D8u917, Qau917, Gdu917, Wfu917, Jiu917;
reg Zku917, Pnu917, Opu917, Mru917, Ktu917, Yvu917, Myu917, N0v917, F3v917, X5v917;
reg R7v917, J9v917, Ebv917, Rdv917, Hgv917, Xiv917, Klv917, Aov917, Qqv917, Dtv917;
reg Tvv917, Jyv917, J0w917, G2w917, G4w917, D6w917, A8w917, X9w917, Rbw917, Ndw917;
reg Jfw917, Fhw917, Bjw917, Ykw917, Smw917, Pow917, Qqw917, Rsw917, Suw917, Tww917;
reg Oyw917, O0x917, O2x917, O4x917, T6x917, E9x917, Pbx917, Mdx917, Efx917, Dhx917;
reg Cjx917, Blx917, Anx917, Zox917, Wqx917, Osx917, Jux917, Lwx917, Nyx917, P0y917;
reg S2y917, Y5y917, P7y917, F9y917, Vay917, Lcy917, Bey917, Rfy917, Hhy917, Xiy917;
reg Nky917, Pmy917, Moy917, Hqy917, Zry917, Lty917, Ovy917, Uxy917, A0z917, N2z917;
reg A5z917, N7z917, Aaz917, Ncz917, Afz917, Nhz917, Bkz917, Pmz917, Dpz917, Rrz917;
reg Fuz917, Twz917, Hzz917, V10a17, J40a17, X60a17, L90a17, Zb0a17, Ne0a17, Bh0a17;
reg Pj0a17, Dm0a17, Qo0a17, Dr0a17, Ot0a17, Bw0a17, Oy0a17, B11a17, R31a17, N61a17;
reg R91a17, Jb1a17, Xd1a17, Lg1a17, Zi1a17, Ml1a17, Po1a17, Or1a17, Nu1a17, Mx1a17;
reg L02a17, K32a17, J62a17, I92a17, Hc2a17, Gf2a17, Ki2a17, Jl2a17, Io2a17, Hr2a17;
reg Gu2a17, Fx2a17, E03a17, D33a17, C63a17, B93a17, Ac3a17, Ze3a17, Yh3a17, Xk3a17;
reg Wn3a17, Vq3a17, Ut3a17, Tw3a17, Sz3a17, R24a17, Q54a17, P84a17, Ob4a17, Ne4a17;
reg Mh4a17, Lk4a17, Kn4a17, Jq4a17, It4a17, Hw4a17, Gz4a17, F25a17, E55a17, C85a17;
reg Bb5a17, Ae5a17, Zg5a17, Yj5a17, Xm5a17, Wp5a17, Vs5a17, Uv5a17, Ty5a17, S16a17;
reg R46a17, Q76a17, Pa6a17, Od6a17, Ng6a17, Lj6a17, Jm6a17, Ip6a17, Hs6a17, Gv6a17;
reg Fy6a17, E17a17, I37a17, H67a17, G97a17, Qb7a17, Ud7a17, Bg7a17, Ei7a17, Ik7a17;
reg Gm7a17, Fo7a17, Eq7a17, Ds7a17, Cu7a17, Bw7a17, Zx7a17, Tz7a17, B28a17, A48a17;
reg O68a17, O88a17, Ma8a17, Kc8a17, Ie8a17, Gg8a17, Ei8a17, Ck8a17, Am8a17, Yn8a17;
reg Wp8a17, Nr8a17, Mt8a17, Dv8a17, Cx8a17, Kz8a17, M19a17, L39a17, I59a17, F79a17;
reg C99a17, Za9a17, Qc9a17, Ne9a17, Kg9a17, Hi9a17, Ek9a17, Bm9a17, Yn9a17, Vp9a17;
reg Sr9a17, Pt9a17, Mv9a17, Jx9a17, Gz9a17, N1aa17, U3aa17, B6aa17, Y7aa17, V9aa17;
reg Sbaa17, Pdaa17, Mfaa17, Jhaa17, Gjaa17, Dlaa17, Anaa17, Xoaa17, Uqaa17, Rsaa17;
reg Ouaa17, Lwaa17, Iyaa17, F0ba17, C2ba17, Z3ba17, W5ba17, T7ba17, Q9ba17, Nbba17;
reg Kdba17, Hfba17, Ohba17, Skba17, Pmba17, Tpba17, Rrba17, Ptba17, Pvba17, Pxba17;
reg Xzba17, F2ca17, N4ca17, K6ca17, H8ca17, Eaca17, Bcca17, Ydca17, Vfca17, Shca17;
reg Pjca17, Mlca17, Jnca17, Gpca17, Drca17, Atca17, Xuca17, Uwca17, Ryca17, O0da17;
reg L2da17, I4da17, F6da17, C8da17, Z9da17, Wbda17, Tdda17, Qfda17, Nhda17, Kjda17;
reg Hlda17, Enda17, Bpda17, Yqda17, Vsda17, Suda17, Pwda17, Myda17, J0ea17, G2ea17;
reg D4ea17, A6ea17, X7ea17, U9ea17, Rbea17, Odea17, Lfea17, Ihea17, Djea17, Blea17;
reg Zmea17, Xoea17, Xqea17, Tsea17, Wvea17, Kyea17, J1fa17, I4fa17, H7fa17, Uafa17;
reg Bdfa17, Iffa17, Phfa17, Wjfa17, Dmfa17, Kofa17, Rqfa17, Ysfa17, Mvfa17, Uxfa17;
reg C0ga17, K2ga17, S4ga17, A7ga17, I9ga17, Qbga17, Ndga17, Cfga17, Rgga17, Giga17;
reg Vjga17, Klga17, Zmga17, Ooga17, Dqga17, Jsga17, Puga17, Mwga17, Bzga17, V0ha17;
reg V2ha17, X5ha17, Z8ha17, Qbha17, Ieha17, Ahha17, Sjha17, Omha17, Gpha17, Yrha17;
reg Quha17, Mxha17, L0ia17, K3ia17, J6ia17, I9ia17, Hcia17, Gfia17, Fiia17, Elia17;
reg Ynia17, Sqia17, Ntia17, Iwia17, Dzia17, Y1ja17, T4ja17, O7ja17, Jaja17, Hdja17;
reg Fgja17, Ejja17, Mlja17, Vnja17, Sqja17, Ptja17, Mwja17, Jzja17, G2ka17, D5ka17;
reg A8ka17, Xaka17, Vdka17, Tgka17, Qjka17, Nmka17, Lpka17, Jska17, Hvka17, Fyka17;
reg D1la17, B4la17, Z6la17, X9la17, Vcla17, Tfla17, Rila17, Plla17, Nola17, Lrla17;
reg Jula17, Hxla17, F0ma17, Z2ma17, T5ma17, N8ma17, Ibma17, Dema17, Ygma17, Tjma17;
reg Omma17, Jpma17, Gsma17, Dvma17, Ayma17, X0na17, U3na17, R6na17, O9na17, Lcna17;
reg Ifna17, Fina17, Dlna17, Bona17, Zqna17, Xtna17, Vwna17, Tzna17, R2oa17, P5oa17;
reg N8oa17, Lboa17, Jeoa17, Hhoa17, Fkoa17, Dnoa17, Bqoa17, Zsoa17, Xvoa17, Vyoa17;
reg T1pa17, R4pa17, O7pa17, Oapa17, Tdpa17, Agpa17, Kipa17, Ukpa17, Enpa17, Oppa17;
reg Mspa17, Kvpa17, Pxpa17, M0qa17, O2qa17, G4qa17, I6qa17, S8qa17, Jbqa17, Aeqa17;
reg Lgqa17, Wiqa17, Hlqa17, Snqa17, Dqqa17, Osqa17, Zuqa17, Kxqa17, Vzqa17, G2ra17;
reg S4ra17, E7ra17, Q9ra17, Ccra17, Oera17, Ahra17, Mjra17, Ylra17, Kora17, Wqra17;
reg Itra17, Uvra17, Gyra17, S0sa17, E3sa17, Q5sa17, C8sa17, Oasa17, Adsa17, Mfsa17;
reg Yhsa17, Kksa17, Rnsa17, Arsa17, Tssa17, Musa17, Fwsa17, Yxsa17, Rzsa17, K1ta17;
reg D3ta17, W4ta17, P6ta17, I8ta17, Cata17, Wbta17, Qdta17, Kfta17, Ehta17, Yita17;
reg Skta17, Mmta17, Gota17, Aqta17, Trta17, Qtta17, Ivta17, Bxta17, Yyta17, Q0ua17;
reg L2ua17, H4ua17, D6ua17, Z7ua17, V9ua17, Rbua17, Ndua17, Jfua17, Fhua17, Bjua17;
reg Xkua17, Tmua17, Poua17, Lqua17, Hsua17, Duua17, Zvua17, Vxua17, Rzua17, N1va17;
reg J3va17, F5va17, B7va17, X8va17, Tava17, Pcva17, Leva17, Hgva17, Diva17, Zjva17;
reg Vlva17, Rnva17, Npva17, Jrva17, Ftva17, Bvva17, Xwva17, Tyva17, P0wa17, K2wa17;
reg F4wa17, A6wa17, V7wa17, Q9wa17, Lbwa17, Gdwa17, Bfwa17, Wgwa17, Oiwa17, Mkwa17;
reg Kmwa17, Iowa17, Fqwa17, Wrwa17, Utwa17, Svwa17, Qxwa17, Ozwa17, K1xa17, M4xa17;
reg O7xa17, Vaxa17, Cexa17, Jhxa17, Skxa17, Knxa17, Cqxa17, Nsxa17, Yuxa17, Qxxa17;
reg I0ya17, T2ya17, E5ya17, P7ya17, Aaya17, Lcya17, Dfya17, Vhya17, Gkya17, Rmya17;
reg Vpya17, Trya17, Rtya17, Ovya17, Lxya17, Izya17, F1za17, C3za17, Z4za17, W6za17;
reg T8za17, Qaza17, Ncza17, Keza17, Hgza17, Eiza17, Bkza17, Ylza17, Vnza17, Spza17;
reg Prza17, Mtza17, Jvza17, Gxza17, Dzza17, A10b17, X20b17, S40b17, Q60b17, O80b17;
reg Ma0b17, Kc0b17, He0b17, Eg0b17, Bi0b17, Yj0b17, Vl0b17, Sn0b17, Pp0b17, Mr0b17;
reg Jt0b17, Gv0b17, Dx0b17, Az0b17, X01b17, U21b17, R41b17, O61b17, L81b17, Ia1b17;
reg Fc1b17, Ce1b17, Zf1b17, Wh1b17, Tj1b17, Ql1b17, Nn1b17, Kp1b17, Hr1b17, Et1b17;
reg Bv1b17, Yw1b17, Vy1b17, S02b17, P22b17, M42b17, J62b17, G82b17, Da2b17, Ac2b17;
reg Xd2b17, Uf2b17, Rh2b17, Oj2b17, Ll2b17, In2b17, Fp2b17, Cr2b17, Zs2b17, Wu2b17;
reg Tw2b17, Qy2b17, N03b17, K23b17, H43b17, E63b17, B83b17, Y93b17, Vb3b17, Sd3b17;
reg Pf3b17, Mh3b17, Jj3b17, Gl3b17, Dn3b17, Ap3b17, Xq3b17, Us3b17, Ru3b17, Ow3b17;
reg Ly3b17, I04b17, F24b17, C44b17, Z54b17, W74b17, T94b17, Qb4b17, Nd4b17, Kf4b17;
reg Hh4b17, Ej4b17, Zk4b17, Xm4b17, Vo4b17, Tq4b17, Rs4b17, Pu4b17, Nw4b17, Uy4b17;
reg X05b17, D45b17, U55b17, K75b17, A95b17, Qa5b17, Gc5b17, Wd5b17, Mf5b17, Ch5b17;
reg Si5b17, Sk5b17, Um5b17, Ro5b17, Cr5b17, Nt5b17, Yv5b17, Jy5b17, U06b17, F36b17;
reg Q56b17, T86b17, Wb6b17, Qe6b17, Tg6b17, Zj6b17, Ql6b17, Gn6b17, Wo6b17, Mq6b17;
reg Cs6b17, St6b17, Iv6b17, Yw6b17, Oy6b17, L07b17, M37b17, Q57b17, R67b17, T77b17;
reg V87b17, W97b17, Xa7b17, Yb7b17, Zc7b17, Yg5m17, Ai5m17, Cj5m17, Ek5m17, Gl5m17;
reg Im5m17, Kn5m17, Mo5m17, Op5m17, Qq5m17, Sr5m17, Us5m17, Wt5m17, Yu5m17, Aw5m17;
reg Cx5m17, Ey5m17, Gz5m17, I06m17, K16m17, M26m17, O36m17, Q46m17, S56m17, U66m17;
reg W76m17, Y86m17, Aa6m17, Cb6m17, Ec6m17, Gd6m17, Ie6m17, Kf6m17, Mg6m17, Oh6m17;
reg Qi6m17, Sj6m17, Uk6m17, Wl6m17, Ym6m17, Ao6m17, Cp6m17, Eq6m17, Gr6m17, Is6m17;
reg Kt6m17, Mu6m17, Ov6m17, Qw6m17, Sx6m17, Uy6m17, Wz6m17, Y07m17, A27m17, B37m17;
reg Z47m17, X67m17, Y87m17, Fb7m17, Je7m17, Nh7m17, Tj7m17, Zl7m17, Fo7m17, Lq7m17;
reg Js7m17, Hu7m17, Fw7m17, Jy7m17, G08m17, N28m17, E58m17, V78m17, Ka8m17, Zc8m17;
reg Ye8m17, Ph8m17, Gk8m17, Nm8m17, Cp8m17, Br8m17, At8m17, Zu8m17, Yw8m17, Fz8m17;
reg W19m17, N49m17, C79m17, R99m17, Yb9m17, Pe9m17, Gh9m17, Vj9m17, Mm9m17, Dp9m17;
reg Or9m17, Du9m17, Ow9m17, Dz9m17, T0am17, I2am17, X3am17, M5am17, B7am17, Q8am17;
reg Faam17, Ubam17, Jdam17, Pfam17, Vham17, Sjam17, Wmam17, Toam17, Zqam17, Ntam17;
reg Tvam17, Qxam17, U0bm17, A3bm17, O5bm17, L7bm17, I9bm17, Tbbm17, Eebm17, Tgbm17;
reg Ejbm17, Plbm17, Eobm17, Pqbm17, Atbm17, Pvbm17, Aybm17, L0cm17, A3cm17, B6cm17;
reg H9cm17, Rbcm17, Pecm17, Mgcm17, Djcm17, Ulcm17, Locm17, Crcm17, Ttcm17, Kwcm17;
reg Bzcm17, S1dm17, J4dm17, B7dm17, T9dm17, Lcdm17, Dfdm17, Vhdm17, Nkdm17, Endm17;
reg Fodm17, Irdm17, Ftdm17, Jwdm17, Mydm17, D0em17, T1em17, J3em17, Z4em17, P6em17;
reg F8em17, V9em17, Lbem17, Bdem17, Dfem17, Ahem17, Ljem17, Wlem17, Loem17, Wqem17;
reg Htem17, Wvem17, Hyem17, S0fm17, H3fm17, S5fm17, D8fm17, Safm17, Tdfm17, Zgfm17;
reg Dkfm17, Rmfm17, Fpfm17, Srfm17, Dufm17, Owfm17, Dzfm17, O1gm17, Z3gm17, O6gm17;
reg Z8gm17, Kbgm17, Zdgm17, Kggm17, Vigm17, Klgm17, Oogm17, Kqgm17, Otgm17, Lvgm17;
reg Lygm17, M1hm17, O2hm17, Q3hm17, R4hm17, O6hm17, Z8hm17, Kbhm17, Zdhm17, Kghm17;
reg Vihm17, Klhm17, Vnhm17, Gqhm17, Vshm17, Gvhm17, Rxhm17, G0im17, J3im17, N6im17;
reg L8im17, Maim17, Pcim17, Vfim17, Mhim17, Cjim17, Skim17, Imim17, Ynim17, Opim17;
reg Erim17, Usim17, Kuim17, Hwim17, Syim17, D1jm17, S3jm17, D6jm17, O8jm17, Dbjm17;
reg Odjm17, Zfjm17, Oijm17, Zkjm17, Knjm17, Zpjm17, Xrjm17, Ytjm17, Ywjm17, D0km17;
reg H3km17, A5km17, T6km17, M8km17, Fakm17, Wbkm17, Pdkm17, Ifkm17, Fhkm17, Yikm17;
reg Alkm17, Xmkm17, Uokm17, Frkm17, Qtkm17, Fwkm17, Qykm17, B1lm17, Q3lm17, B6lm17;
reg M8lm17, Bblm17, Mdlm17, Xflm17, Milm17, Xklm17, Inlm17, Xplm17, Xrlm17, Vtlm17;
reg Wvlm17, Xylm17, Y1mm17, Z4mm17, E8mm17, Abmm17, Wdmm17, Sgmm17, Mjmm17, Cmmm17;
reg Xomm17, Asmm17, Vumm17, Yxmm17, T0nm17, W3nm17, R6nm17, M9nm17, Pcnm17, Kfnm17;
reg Ninm17, Ilnm17, Lonm17, Grnm17, Junm17, Exnm17, I0om17, D3om17, H6om17, L9om17;
reg Pcom17, Tfom17, Xiom17, Bmom17, Fpom17, Jsom17, Nvom17, Ryom17, V1pm17, Z4pm17;
reg D8pm17, Hbpm17, Lepm17, Phpm17, Tkpm17, Xnpm17, Brpm17, Fupm17, Jxpm17, M0qm17;
reg P3qm17, A5qm17, Y6qm17, Z8qm17, Xaqm17, Wcqm17, Veqm17, Ugqm17, Tiqm17, Skqm17;
reg Rmqm17, Qoqm17, Rqqm17, Ssqm17, Tuqm17, Uwqm17, Syqm17, T0rm17, Q2rm17, B5rm17;
reg M7rm17, Barm17, Mcrm17, Xerm17, Mhrm17, Xjrm17, Imrm17, Xorm17, Irrm17, Ttrm17;
reg Iwrm17, Tyrm17, E1sm17, T3sm17, V5sm17, N7sm17, A9sm17, Oasm17, Rdsm17, Ugsm17;
reg Ajsm17, Tksm17, Jnsm17, Dqsm17, Assm17, Uusm17, Sxsm17, Q0tm17, O3tm17, M6tm17;
reg K9tm17, Ictm17, Fftm17, Dhtm17, Ejtm17, Fltm17, Vntm17, Lqtm17, Bttm17, Svtm17;
reg Jytm17, A1um17, R3um17, I6um17, Z8um17, Qbum17, Heum17, Ygum17, Pjum17, Gmum17;
reg Xoum17, Orum17, Fuum17, Wwum17, Nzum17, E2vm17, V4vm17, M7vm17, Davm17, Ucvm17;
reg Lfvm17, Ihvm17, Gjvm17, Hlvm17, Invm17, Gpvm17, Ksvm17, Duvm17, Wvvm17, Pxvm17;
reg Izvm17, B1wm17, U2wm17, N4wm17, G6wm17, Z7wm17, W9wm17, Tbwm17, Udwm17, Vfwm17;
reg Thwm17, Rjwm17;
wire [33:0] Llwm17;
wire [33:0] Cnwm17;
wire [4:0] Towm17;
wire [33:0] Jqwm17;
wire [33:0] Dswm17;
wire [31:0] Puwm17;
wire [31:0] Dxwm17;
wire [33:0] Rzwm17;
wire [33:0] H2xm17;
wire [63:0] W4xm17;
wire [30:0] Y6xm17;
wire [30:0] A9xm17;
wire [33:0] Cbxm17;
wire [33:0] Edxm17;
wire [33:0] Gfxm17;
wire [33:0] Cixm17;
wire [33:0] Wkxm17;
wire [33:0] Snxm17;
wire [31:0] Mqxm17;
wire [33:0] Wtxm17;
wire [31:0] Gxxm17;
wire [33:0] Q0ym17;
wire [33:0] A4ym17;
wire [33:0] K7ym17;
wire [33:0] Uaym17;
wire [33:0] Ldym17;
wire [33:0] Agym17;
wire [33:0] Riym17;
wire [63:0] Glym17;
wire [5:0] Xnym17;
wire [31:0] Mqym17;
wire [33:0] Etym17;
wire [6:0] Uvym17;
wire [33:0] Jyym17;
wire [33:0] H1zm17;
wire [33:0] F4zm17;
wire [33:0] D7zm17;
wire [33:0] Z9zm17;

assign HTRANSI[0] = 1'b0;
assign HADDRI[1] = 1'b0;
assign HADDRI[0] = 1'b0;
assign HSIZES[2] = 1'b0;
assign HBURSTD[1] = 1'b0;
assign HBURSTD[2] = 1'b0;
assign HBURSTS[1] = 1'b0;
assign HBURSTS[2] = 1'b0;
assign CURRPRI[4] = 1'b0;
assign CURRPRI[3] = 1'b0;
assign CURRPRI[2] = 1'b0;
assign CURRPRI[1] = 1'b0;
assign CURRPRI[0] = 1'b0;
assign HTMDHSIZE[2] = 1'b0;
assign HTMDHPROT[3] = 1'b0;
assign HTMDHPROT[2] = 1'b0;
assign HTMDHRDATA[31] = HTMDHWDATA[31];
assign HTMDHRDATA[30] = HTMDHWDATA[30];
assign HTMDHRDATA[29] = HTMDHWDATA[29];
assign HTMDHRDATA[28] = HTMDHWDATA[28];
assign HTMDHRDATA[27] = HTMDHWDATA[27];
assign HTMDHRDATA[26] = HTMDHWDATA[26];
assign HTMDHRDATA[25] = HTMDHWDATA[25];
assign HTMDHRDATA[24] = HTMDHWDATA[24];
assign HTMDHRDATA[23] = HTMDHWDATA[23];
assign HTMDHRDATA[22] = HTMDHWDATA[22];
assign HTMDHRDATA[21] = HTMDHWDATA[21];
assign HTMDHRDATA[20] = HTMDHWDATA[20];
assign HTMDHRDATA[19] = HTMDHWDATA[19];
assign HTMDHRDATA[18] = HTMDHWDATA[18];
assign HTMDHRDATA[17] = HTMDHWDATA[17];
assign HTMDHRDATA[16] = HTMDHWDATA[16];
assign HTMDHRDATA[15] = HTMDHWDATA[15];
assign HTMDHRDATA[14] = HTMDHWDATA[14];
assign HTMDHRDATA[13] = HTMDHWDATA[13];
assign HTMDHRDATA[12] = HTMDHWDATA[12];
assign HTMDHRDATA[11] = HTMDHWDATA[11];
assign HTMDHRDATA[10] = HTMDHWDATA[10];
assign HTMDHRDATA[9] = HTMDHWDATA[9];
assign HTMDHRDATA[8] = HTMDHWDATA[8];
assign HTMDHRDATA[7] = HTMDHWDATA[7];
assign HTMDHRDATA[6] = HTMDHWDATA[6];
assign HTMDHRDATA[5] = HTMDHWDATA[5];
assign HTMDHRDATA[4] = HTMDHWDATA[4];
assign HTMDHRDATA[3] = HTMDHWDATA[3];
assign HTMDHRDATA[2] = HTMDHWDATA[2];
assign HTMDHRDATA[1] = HTMDHWDATA[1];
assign HTMDHRDATA[0] = HTMDHWDATA[0];
assign HBURSTI[2] = 1'b0;
assign HBURSTI[1] = 1'b0;
assign HBURSTI[0] = 1'b0;
assign HSIZEI[1] = 1'b1;
assign HSIZEI[0] = 1'b0;
assign HADDRI[31] = 1'b0;
assign HADDRI[30] = 1'b0;
assign HADDRI[29] = 1'b0;
assign HSIZEI[2] = 1'b0;
assign HPROTI[2] = 1'b0;
assign MEMATTRI[1] = 1'b0;
assign HPROTI[3] = 1'b1;
assign MEMATTRI[0] = 1'b1;
assign HADDRD[31] = 1'b0;
assign HADDRD[30] = 1'b0;
assign HADDRD[29] = 1'b0;
assign HSIZED[2] = 1'b0;
assign HPROTD[2] = 1'b0;
assign MEMATTRD[1] = 1'b0;
assign HPROTD[3] = 1'b1;
assign MEMATTRD[0] = 1'b1;
assign TRCENA = HTMDHBURST[0];
assign HTMDHBURST[2] = 1'b0;
assign HTMDHBURST[1] = 1'b0;
assign M4adt6 = Sj2nz6;
assign Cy9dt6 = Ik2nz6;
assign Y4adt6 = Zk2nz6;
assign Ez9dt6 = Ql2nz6;
assign L5adt6 = Im2nz6;
assign G0adt6 = Ym2nz6;
assign X5adt6 = Pn2nz6;
assign D1adt6 = Go2nz6;
assign Aabdt6 = Yo2nz6;
assign Kr97z6 = Eq2nz6;
assign Cbbdt6 = Er2nz6;
assign Cb77z6 = Hs2nz6;
assign Bcbdt6 = Et2nz6;
assign Cwadt6 = Su2nz6;
assign Dwb7z6[0] = Aw2nz6;
assign Dwb7z6[1] = Ny2nz6;
assign Dwb7z6[2] = A13nz6;
assign Dwb7z6[3] = N33nz6;
assign Dwb7z6[4] = A63nz6;
assign Dwb7z6[5] = N83nz6;
assign Ffeet6 = Ab3nz6;
assign Cr97z6 = (!Cd3nz6);
assign Evadt6 = Bf3nz6;
assign Jd47v6 = Yg3nz6;
assign Mp67v6 = Xh3nz6;
assign Gj47v6 = Vj3nz6;
assign Tah7v6 = Ul3nz6;
assign I977v6 = Un3nz6;
assign Fy67v6 = Ip3nz6;
assign Gg77v6 = Vq3nz6;
assign Dp77v6 = Ms3nz6;
assign TRACECLK = Su3nz6;
assign Tho7v6 = (!Su3nz6);
assign Ti2nz6[5] = Mw3nz6;
assign Pdc7z6[26] = Sx3nz6;
assign Kxb7z6[26] = T04nz6;
assign Fth7z6[31] = D34nz6;
assign Wlr7z6[31] = B64nz6;
assign K0wmz6[7] = P84nz6;
assign Nsvmz6[7] = Ab4nz6;
assign La6ft6 = Pd4nz6;
assign V7xmz6[7] = Jf4nz6;
assign V7xmz6[1] = Jh4nz6;
assign Pp1nz6[1] = Jj4nz6;
assign U81nz6[1] = Hl4nz6;
assign J1h7v6 = Un4nz6;
assign Af1nz6[1] = Nq4nz6;
assign Itb7z6[0] = Gt4nz6;
assign Tim7z6[0] = Yv4nz6;
assign Zec7z6[16] = My4nz6;
assign Dvc7z6[31] = L15nz6;
assign Hrb7z6[1] = R45nz6;
assign Zec7z6[15] = H65nz6;
assign Byc7z6[15] = G95nz6;
assign Zec7z6[31] = Kc5nz6;
assign Lvg7z6[3] = Jf5nz6;
assign Vi7et6 = Mi5nz6;
assign Fth7z6[0] = Kl5nz6;
assign Kxb7z6[0] = Ho5nz6;
assign D6gdt6 = Qq5nz6;
assign X9s7z6[38] = Rs5nz6;
assign Gyvmz6[6] = Ou5nz6;
assign Nsvmz6[6] = Zw5nz6;
assign V7xmz6[6] = Oz5nz6;
assign Mm1nz6[6] = O16nz6;
assign Pdc7z6[30] = M36nz6;
assign Kxb7z6[30] = N66nz6;
assign Alf7z6[31] = X86nz6;
assign Yxf7z6[0] = Vb6nz6;
assign Yxf7z6[4] = Pe6nz6;
assign Yxf7z6[8] = Jh6nz6;
assign Yxf7z6[12] = Dk6nz6;
assign Yxf7z6[16] = Ym6nz6;
assign Yxf7z6[20] = Tp6nz6;
assign Yxf7z6[24] = Os6nz6;
assign Yxf7z6[28] = Jv6nz6;
assign Yxf7z6[32] = Ey6nz6;
assign O4gdt6 = Z07nz6;
assign Tim7z6[31] = A37nz6;
assign Itb7z6[31] = P57nz6;
assign Dto7z6[1] = H87nz6;
assign Woyet6 = Z97nz6;
assign Znn7z6[1] = Oc7nz6;
assign Hjn7z6[6] = Af7nz6;
assign Tim7z6[30] = Qh7nz6;
assign Fth7z6[6] = Fk7nz6;
assign Pdc7z6[6] = Cn7nz6;
assign Kxb7z6[6] = Cq7nz6;
assign Onf7z6[31] = Ls7nz6;
assign Yxf7z6[3] = Jv7nz6;
assign Yxf7z6[7] = Dy7nz6;
assign Yxf7z6[11] = X08nz6;
assign Yxf7z6[15] = S38nz6;
assign Yxf7z6[19] = N68nz6;
assign Yxf7z6[23] = I98nz6;
assign Yxf7z6[27] = Dc8nz6;
assign Yxf7z6[31] = Ye8nz6;
assign H9gdt6 = Th8nz6;
assign X9s7z6[36] = Uj8nz6;
assign Gyvmz6[4] = Rl8nz6;
assign Nsvmz6[4] = Co8nz6;
assign V7xmz6[4] = Rq8nz6;
assign Mm1nz6[4] = Rs8nz6;
assign Pdc7z6[28] = Pu8nz6;
assign Kxb7z6[28] = Qx8nz6;
assign Fre7z6[0] = A09nz6;
assign Elgdt6 = X29nz6;
assign Onf7z6[30] = R59nz6;
assign D5f7z6[5] = P89nz6;
assign Bdf7z6[1] = Lb9nz6;
assign K1i7z6[0] = Le9nz6;
assign V5k7z6[31] = Oh9nz6;
assign Fth7z6[30] = Ik9nz6;
assign M6j7z6[63] = Gn9nz6;
assign Itbet6 = Fq9nz6;
assign M6bdt6 = Ct9nz6;
assign Oc47v6 = Av9nz6;
assign Uq97z6 = Zv9nz6;
assign Mq97z6 = Zw9nz6;
assign Eq97z6 = Zx9nz6;
assign Wp97z6 = Zy9nz6;
assign Op97z6 = Zz9nz6;
assign Gp97z6 = Z0anz6;
assign Yo97z6 = Z1anz6;
assign Qo97z6 = Z2anz6;
assign Io97z6 = Z3anz6;
assign Ao97z6 = Z4anz6;
assign Sn97z6 = A6anz6;
assign Kn97z6 = B7anz6;
assign Cn97z6 = C8anz6;
assign Um97z6 = D9anz6;
assign Mm97z6 = Eaanz6;
assign Em97z6 = Fbanz6;
assign Wl97z6 = Gcanz6;
assign Ol97z6 = Hdanz6;
assign Gl97z6 = Ieanz6;
assign Yk97z6 = Jfanz6;
assign Qk97z6 = Kganz6;
assign Ik97z6 = Lhanz6;
assign Ak97z6 = Mianz6;
assign Sj97z6 = Njanz6;
assign Kj97z6 = Okanz6;
assign Cj97z6 = Planz6;
assign Ui97z6 = Qmanz6;
assign Mi97z6 = Rnanz6;
assign Ei97z6 = Soanz6;
assign Wh97z6 = Tpanz6;
assign Oh97z6 = Uqanz6;
assign Gh97z6 = Vranz6;
assign Yg97z6 = Wsanz6;
assign Qg97z6 = Xtanz6;
assign Ig97z6 = Yuanz6;
assign Ag97z6 = Zvanz6;
assign Sf97z6 = Axanz6;
assign Kf97z6 = Byanz6;
assign Cf97z6 = Czanz6;
assign Ue97z6 = D0bnz6;
assign Me97z6 = E1bnz6;
assign Ee97z6 = F2bnz6;
assign Wd97z6 = G3bnz6;
assign Od97z6 = H4bnz6;
assign Gd97z6 = I5bnz6;
assign Yc97z6 = J6bnz6;
assign Qc97z6 = K7bnz6;
assign Ic97z6 = L8bnz6;
assign Ac97z6 = M9bnz6;
assign Sb97z6 = Nabnz6;
assign Kb97z6 = Obbnz6;
assign Cb97z6 = Pcbnz6;
assign Ua97z6 = Qdbnz6;
assign Ma97z6 = Rebnz6;
assign Ea97z6 = Sfbnz6;
assign W997z6 = Tgbnz6;
assign O997z6 = Uhbnz6;
assign G997z6 = Vibnz6;
assign Y897z6 = Wjbnz6;
assign Q897z6 = Xkbnz6;
assign I897z6 = Ylbnz6;
assign A897z6 = Zmbnz6;
assign S797z6 = Aobnz6;
assign K797z6 = Bpbnz6;
assign C797z6 = Cqbnz6;
assign Ei77z6 = Drbnz6;
assign U697z6 = Dsbnz6;
assign Jqj7z6[0] = Etbnz6;
assign Jqj7z6[72] = Fwbnz6;
assign Jqj7z6[71] = Hzbnz6;
assign Jqj7z6[70] = J2cnz6;
assign Jqj7z6[69] = L5cnz6;
assign Jqj7z6[68] = N8cnz6;
assign Jqj7z6[67] = Pbcnz6;
assign Jqj7z6[66] = Recnz6;
assign Jqj7z6[65] = Thcnz6;
assign Jqj7z6[64] = Vkcnz6;
assign Jqj7z6[63] = Xncnz6;
assign Jqj7z6[62] = Zqcnz6;
assign Jqj7z6[61] = Bucnz6;
assign Jqj7z6[60] = Dxcnz6;
assign Jqj7z6[59] = F0dnz6;
assign Jqj7z6[58] = H3dnz6;
assign Jqj7z6[57] = J6dnz6;
assign Jqj7z6[56] = L9dnz6;
assign Jqj7z6[55] = Ncdnz6;
assign Jqj7z6[54] = Pfdnz6;
assign Jqj7z6[53] = Ridnz6;
assign Jqj7z6[52] = Tldnz6;
assign Jqj7z6[51] = Vodnz6;
assign Jqj7z6[50] = Xrdnz6;
assign Jqj7z6[49] = Zudnz6;
assign Jqj7z6[48] = Bydnz6;
assign Jqj7z6[47] = D1enz6;
assign Jqj7z6[46] = F4enz6;
assign Jqj7z6[45] = H7enz6;
assign Jqj7z6[44] = Jaenz6;
assign Jqj7z6[43] = Ldenz6;
assign Jqj7z6[42] = Ngenz6;
assign Jqj7z6[41] = Pjenz6;
assign Jqj7z6[40] = Rmenz6;
assign Jqj7z6[39] = Tpenz6;
assign Jqj7z6[38] = Vsenz6;
assign Jqj7z6[37] = Xvenz6;
assign Jqj7z6[36] = Zyenz6;
assign Jqj7z6[35] = B2fnz6;
assign Jqj7z6[34] = D5fnz6;
assign Jqj7z6[33] = F8fnz6;
assign Jqj7z6[32] = Hbfnz6;
assign Jqj7z6[31] = Jefnz6;
assign Jqj7z6[30] = Lhfnz6;
assign Jqj7z6[29] = Nkfnz6;
assign Jqj7z6[28] = Pnfnz6;
assign Jqj7z6[27] = Rqfnz6;
assign Jqj7z6[26] = Ttfnz6;
assign Jqj7z6[25] = Vwfnz6;
assign Jqj7z6[24] = Xzfnz6;
assign Jqj7z6[23] = Z2gnz6;
assign Jqj7z6[22] = B6gnz6;
assign Jqj7z6[21] = D9gnz6;
assign Jqj7z6[20] = Fcgnz6;
assign Jqj7z6[19] = Hfgnz6;
assign Jqj7z6[18] = Jignz6;
assign Jqj7z6[17] = Llgnz6;
assign Jqj7z6[16] = Nognz6;
assign Jqj7z6[15] = Prgnz6;
assign Jqj7z6[14] = Rugnz6;
assign Jqj7z6[13] = Txgnz6;
assign Jqj7z6[12] = V0hnz6;
assign Jqj7z6[11] = X3hnz6;
assign Jqj7z6[10] = Z6hnz6;
assign Jqj7z6[9] = Bahnz6;
assign Jqj7z6[1] = Cdhnz6;
assign V5get6 = Dghnz6;
assign Ldh7v6 = (!Bjhnz6);
assign Kkadt6 = Elhnz6;
assign Aiadt6 = Cnhnz6;
assign Cgc7z6[2] = Hphnz6;
assign Vjddt6 = Yrhnz6;
assign Dvc7z6[10] = Tuhnz6;
assign Hrb7z6[0] = Zxhnz6;
assign Zec7z6[23] = Pzhnz6;
assign Byc7z6[23] = O2inz6;
assign Zec7z6[7] = S5inz6;
assign V1c7z6[5] = Q8inz6;
assign Nzg7z6[0] = Vainz6;
assign Nzg7z6[1] = Xdinz6;
assign Nzg7z6[2] = Zginz6;
assign Nzg7z6[3] = Bkinz6;
assign Wfxdt6 = Dninz6;
assign Sj77z6 = (!Tpinz6);
assign K73et6 = Osinz6;
assign Pl7et6 = Kvinz6;
assign M697z6 = (!Myinz6);
assign Bzi7z6[1] = O1jnz6;
assign Nneet6 = N3jnz6;
assign HALTED = S5jnz6;
assign Ldo7v6 = (!S5jnz6);
assign Z2c7v6 = Q7jnz6;
assign I1c7v6 = P9jnz6;
assign Sdh7v6 = (!Objnz6);
assign DBGRESTARTED = Qdjnz6;
assign Dgo7v6 = (!Qdjnz6);
assign Cbeet6 = Wfjnz6;
assign Opeet6 = Bijnz6;
assign Jjbdt6 = Fkjnz6;
assign Uyb7z6[2] = Gmjnz6;
assign Pdc7z6[2] = Qojnz6;
assign Kxb7z6[2] = Qrjnz6;
assign Ir7et6 = Ztjnz6;
assign Cjq7z6[0] = Fxjnz6;
assign C4s7z6[1] = Lzjnz6;
assign V1s7z6[0] = P2knz6;
assign Sywmz6[0] = D5knz6;
assign Kms7z6[0] = O7knz6;
assign V7xmz6[0] = Daknz6;
assign Nn1nz6[0] = Dcknz6;
assign Pdc7z6[24] = Beknz6;
assign Kxb7z6[24] = Chknz6;
assign Fth7z6[24] = Mjknz6;
assign Oreet6 = Kmknz6;
assign Iladt6 = Qoknz6;
assign Cgc7z6[1] = Vqknz6;
assign Nbddt6 = Mtknz6;
assign Dvc7z6[11] = Jwknz6;
assign Ccnet6 = Pzknz6;
assign Ywcdt6 = J2lnz6;
assign Pdc7z6[1] = L5lnz6;
assign Kxb7z6[1] = L8lnz6;
assign Fth7z6[1] = Ualnz6;
assign Zec7z6[0] = Rdlnz6;
assign V1c7z6[0] = Pglnz6;
assign Kxb7z6[8] = Uilnz6;
assign Fth7z6[8] = Dllnz6;
assign Pdc7z6[8] = Aolnz6;
assign Dvc7z6[8] = Arlnz6;
assign A3ddt6 = Fulnz6;
assign X7get6 = Exlnz6;
assign Byi7z6[31] = Azlnz6;
assign Fth7z6[7] = A1mnz6;
assign Pdc7z6[7] = X3mnz6;
assign Kxb7z6[7] = X6mnz6;
assign Fhc7z6[31] = G9mnz6;
assign Kxb7z6[4] = Qbmnz6;
assign Fth7z6[4] = Zdmnz6;
assign Pdc7z6[4] = Wgmnz6;
assign Dvc7z6[30] = Wjmnz6;
assign U4zet6 = Cnmnz6;
assign N7zet6 = Zpmnz6;
assign Ysn7z6[0] = Wsmnz6;
assign Ysn7z6[2] = Xvmnz6;
assign Ysn7z6[1] = Yymnz6;
assign Khoet6 = Z1nnz6;
assign Wmoet6 = X4nnz6;
assign Ihs7z6[1] = T7nnz6;
assign Ci27v6 = N9nnz6;
assign Zas7z6[2] = Gbnnz6;
assign Tl6ft6 = Wcnnz6;
assign Gyvmz6[8] = Sennz6;
assign Nsvmz6[8] = Dhnnz6;
assign Fbxmz6[1] = Sjnnz6;
assign Fbxmz6[0] = Plnnz6;
assign Mm1nz6[5] = Mnnnz6;
assign Pdc7z6[29] = Kpnnz6;
assign Kxb7z6[29] = Lsnnz6;
assign Fth7z6[29] = Vunnz6;
assign Wui7z6[13] = Txnnz6;
assign Pdc7z6[21] = Vznnz6;
assign Kxb7z6[21] = W2onz6;
assign Fth7z6[21] = G5onz6;
assign Fpo7z6[19] = E8onz6;
assign Ygh7v6 = (!U9onz6);
assign Zbpet6 = U9onz6;
assign Hryet6 = Nbonz6;
assign Qln7z6[0] = Ceonz6;
assign Wzxet6 = Sgonz6;
assign Tim7z6[24] = Ijonz6;
assign Zec7z6[8] = Xlonz6;
assign Byc7z6[8] = Voonz6;
assign Zec7z6[24] = Yronz6;
assign V1c7z6[8] = Xuonz6;
assign Kxb7z6[31] = Cxonz6;
assign Bdf7z6[0] = Mzonz6;
assign Kxb7z6[3] = M2pnz6;
assign Fth7z6[3] = V4pnz6;
assign X9s7z6[19] = S7pnz6;
assign Sywmz6[3] = P9pnz6;
assign Kms7z6[3] = Acpnz6;
assign V7xmz6[3] = Pepnz6;
assign Mm1nz6[3] = Pgpnz6;
assign Pdc7z6[27] = Nipnz6;
assign Kxb7z6[27] = Olpnz6;
assign Fth7z6[27] = Ynpnz6;
assign Kfq7z6[0] = Wqpnz6;
assign V1s7z6[2] = Etpnz6;
assign Sywmz6[2] = Svpnz6;
assign Kms7z6[2] = Dypnz6;
assign V7xmz6[2] = S0qnz6;
assign Mm1nz6[2] = S2qnz6;
assign Pdc7z6[18] = Q4qnz6;
assign Kxb7z6[18] = R7qnz6;
assign Fth7z6[18] = Baqnz6;
assign Z3j7z6[10] = Zcqnz6;
assign Fhcet6 = Xfqnz6;
assign P2j7z6[1] = Viqnz6;
assign M6j7z6[5] = Zkqnz6;
assign P2j7z6[0] = Ynqnz6;
assign Z3j7z6[13] = Cqqnz6;
assign P2j7z6[4] = Atqnz6;
assign M6j7z6[15] = Evqnz6;
assign P2j7z6[2] = Dyqnz6;
assign M6j7z6[55] = H0rnz6;
assign P2j7z6[3] = G3rnz6;
assign Sgcdt6 = K5rnz6;
assign Pdc7z6[25] = O8rnz6;
assign Kxb7z6[25] = Pbrnz6;
assign Fth7z6[25] = Zdrnz6;
assign Wui7z6[9] = Xgrnz6;
assign Pdc7z6[17] = Yirnz6;
assign Kxb7z6[17] = Zlrnz6;
assign Fth7z6[17] = Jornz6;
assign Cjq7z6[1] = Hrrnz6;
assign Cjq7z6[7] = Ntrnz6;
assign Pdc7z6[23] = Tvrnz6;
assign Kxb7z6[23] = Uyrnz6;
assign Fth7z6[23] = E1snz6;
assign Xch7v6 = (!C4snz6);
assign Lfp7z6[1] = F6snz6;
assign Eo2ft6 = F8snz6;
assign Lybdt6 = Hasnz6;
assign Fccdt6 = Fcsnz6;
assign T8ddt6 = Jesnz6;
assign Ztcdt6 = Hhsnz6;
assign Ujnet6 = Kksnz6;
assign Crcdt6 = Xmsnz6;
assign Aocdt6 = Ypsnz6;
assign Kqm7z6[2] = Etsnz6;
assign Zec7z6[13] = Ewsnz6;
assign Byc7z6[13] = Dzsnz6;
assign Zec7z6[29] = H2tnz6;
assign V1c7z6[15] = G5tnz6;
assign Kxb7z6[22] = M7tnz6;
assign Fth7z6[22] = W9tnz6;
assign Xu67v6 = Uctnz6;
assign Uu0nz6[4] = Oetnz6;
assign Rr0nz6[0] = Mgtnz6;
assign Ocd7v6 = Kitnz6;
assign Hw0nz6[2] = Jktnz6;
assign E5d7v6 = Hmtnz6;
assign Hw0nz6[1] = Fotnz6;
assign Rr0nz6[1] = Dqtnz6;
assign Ak67z6 = Bstnz6;
assign Bv1nz6[0] = Wttnz6;
assign Ja1nz6[2] = Uvtnz6;
assign Fwg7v6 = Hytnz6;
assign Fg1nz6[2] = A1unz6;
assign Ja1nz6[1] = T3unz6;
assign Qtg7v6 = G6unz6;
assign Fg1nz6[1] = Z8unz6;
assign Zs1nz6[0] = Sbunz6;
assign Au1nz6[0] = Qdunz6;
assign Yr1nz6[0] = Ofunz6;
assign Yr1nz6[1] = Mhunz6;
assign Pdc7z6[9] = Kjunz6;
assign Kxb7z6[9] = Kmunz6;
assign Fth7z6[9] = Tounz6;
assign Wui7z6[25] = Qrunz6;
assign M43et6 = Stunz6;
assign Jqj7z6[4] = Uwunz6;
assign Jqj7z6[6] = Vzunz6;
assign Oecet6 = W2vnz6;
assign P2j7z6[6] = U5vnz6;
assign P2j7z6[5] = Y7vnz6;
assign Tnzdt6 = Cavnz6;
assign Cgc7z6[0] = Ccvnz6;
assign Cgc7z6[3] = Tevnz6;
assign Fsc7z6[0] = Khvnz6;
assign W8h7v6 = (!Pkvnz6);
assign Inadt6 = Smvnz6;
assign Fjadt6 = Rovnz6;
assign Mmddt6 = Prvnz6;
assign E697z6 = (!Stvnz6);
assign V5ddt6 = Wvvnz6;
assign Pkbet6 = Yyvnz6;
assign Fhc7z6[30] = D1wnz6;
assign Lsfdt6 = N3wnz6;
assign Wui7z6[27] = O5wnz6;
assign Pdc7z6[19] = Q7wnz6;
assign Kxb7z6[19] = Rawnz6;
assign Fth7z6[19] = Bdwnz6;
assign Ipymz6[0] = Zfwnz6;
assign Gm77v6 = Fiwnz6;
assign Pdc7z6[11] = Lkwnz6;
assign vis_psp_o[11] = Mnwnz6;
assign Fhc7z6[11] = Eqwnz6;
assign Kxb7z6[20] = Oswnz6;
assign Fth7z6[20] = Yuwnz6;
assign Fpo7z6[10] = Wxwnz6;
assign Fth7z6[12] = Mzwnz6;
assign Pdc7z6[12] = K2xnz6;
assign Kxb7z6[12] = L5xnz6;
assign Pdq7z6[0] = V7xnz6;
assign Pdq7z6[6] = Baxnz6;
assign Pdc7z6[14] = Hcxnz6;
assign Kxb7z6[14] = Ifxnz6;
assign Fth7z6[14] = Shxnz6;
assign Hhq7z6[6] = Qkxnz6;
assign Hhq7z6[5] = Wmxnz6;
assign S7gdt6 = Cpxnz6;
assign Wui7z6[29] = Drxnz6;
assign Pdc7z6[13] = Ftxnz6;
assign Kxb7z6[13] = Gwxnz6;
assign Fth7z6[13] = Qyxnz6;
assign Pk1nz6[5] = O1ynz6;
assign Td2nz6[0] = L3ynz6;
assign Vuf7v6 = J5ynz6;
assign W3e7v6 = E7ynz6;
assign Thg7v6 = Y8ynz6;
assign Imh7v6 = Ebynz6;
assign W597z6 = (!Kdynz6);
assign We6ft6 = Gfynz6;
assign Qb6ft6 = Chynz6;
assign Vis7z6[5] = Yiynz6;
assign P7s7z6[29] = Xkynz6;
assign E46ft6 = Rmynz6;
assign Nu27v6 = Hoynz6;
assign Iuvmz6[5] = Gqynz6;
assign Iuvmz6[6] = Gsynz6;
assign Iuvmz6[7] = Guynz6;
assign Iuvmz6[8] = Gwynz6;
assign Iuvmz6[4] = Gyynz6;
assign Y4wmz6[0] = G0znz6;
assign Gyvmz6[7] = Y2znz6;
assign Y4wmz6[1] = J5znz6;
assign K0wmz6[4] = B8znz6;
assign K0wmz6[6] = Maznz6;
assign K0wmz6[8] = Xcznz6;
assign Bewmz6[0] = Ifznz6;
assign Bewmz6[1] = Aiznz6;
assign J7wmz6[8] = Skznz6;
assign Ly37v6 = Dnznz6;
assign Fth7z6[15] = Kpznz6;
assign Pdc7z6[15] = Isznz6;
assign Kxb7z6[15] = Jvznz6;
assign Z3j7z6[7] = Txznz6;
assign Z3j7z6[15] = R00oz6;
assign Moj7z6[2] = P30oz6;
assign Zgadt6 = T50oz6;
assign W9edt6 = T70oz6;
assign Mfe7z6[3] = Ba0oz6;
assign Ohe7z6[7] = Ec0oz6;
assign Mfe7z6[7] = Ge0oz6;
assign H3adt6 = Jg0oz6;
assign Wfo7v6 = (!Jg0oz6);
assign Q087v6 = Ki0oz6;
assign W577v6 = Ek0oz6;
assign Gdc7v6 = Em0oz6;
assign Hqb7v6 = Io0oz6;
assign Jsb7v6 = Sq0oz6;
assign Tkb7v6 = Qs0oz6;
assign Bhb7v6 = Wu0oz6;
assign Ifb7v6 = Xw0oz6;
assign Bq0nz6[6] = Yy0oz6;
assign Kj67z6 = V01oz6;
assign Au1nz6[6] = Q21oz6;
assign Zs1nz6[6] = O41oz6;
assign Ohe7z6[6] = M61oz6;
assign Mfe7z6[6] = O81oz6;
assign Yl2et6 = Ra1oz6;
assign Dqr8v6 = (!Md1oz6);
assign Oaadt6 = Eg1oz6;
assign Hhq7z6[4] = Ji1oz6;
assign Qmb7z6[4] = Pk1oz6;
assign Nob7z6[4] = Ln1oz6;
assign D4b7v6 = Qp1oz6;
assign Jjh7v6 = (!Or1oz6);
assign O777v6 = Zt1oz6;
assign Xw67v6 = Wv1oz6;
assign Lzb7v6 = Jx1oz6;
assign Tf87v6 = Oz1oz6;
assign B41nz6[1] = H12oz6;
assign B41nz6[0] = H32oz6;
assign Zwzmz6[7] = H52oz6;
assign Sj67z6 = E72oz6;
assign Au1nz6[7] = Z82oz6;
assign Zs1nz6[7] = Xa2oz6;
assign Ppb7z6[7] = Vc2oz6;
assign Z7edt6 = Df2oz6;
assign Tkbdt6 = Eh2oz6;
assign Fsc7z6[1] = Gj2oz6;
assign Pxg7z6[0] = Lm2oz6;
assign P4c7z6[0] = Ip2oz6;
assign E8h7z6[0] = Fs2oz6;
assign vis_r3_o[0] = Cv2oz6;
assign vis_r3_o[30] = Sx2oz6;
assign vis_r3_o[11] = J03oz6;
assign vis_r3_o[1] = A33oz6;
assign E3c7z6[1] = Q53oz6;
assign Kxb7z6[10] = Z73oz6;
assign Fth7z6[10] = Ja3oz6;
assign O597z6 = (!Hd3oz6);
assign Dkm7z6[1] = Tg3oz6;
assign S7n7z6[0] = Sj3oz6;
assign Pdc7z6[16] = Lm3oz6;
assign Kxb7z6[16] = Mp3oz6;
assign Fth7z6[16] = Wr3oz6;
assign U9p7z6[24] = Uu3oz6;
assign Lfp7z6[0] = Ww3oz6;
assign Fgzmz6[0] = Wy3oz6;
assign Lczmz6[0] = A14oz6;
assign Lczmz6[1] = J34oz6;
assign Lczmz6[2] = S54oz6;
assign Lczmz6[3] = B84oz6;
assign Bq0nz6[3] = Ka4oz6;
assign Mi67z6 = Hc4oz6;
assign Au1nz6[3] = Ce4oz6;
assign Zs1nz6[3] = Ag4oz6;
assign Ohe7z6[5] = Yh4oz6;
assign Mfe7z6[5] = Ak4oz6;
assign Xkr8v6 = (!Dm4oz6);
assign Wzcdt6 = Vo4oz6;
assign P6d7z6[0] = Ds4oz6;
assign Vbh7v6 = (!Gv4oz6);
assign L9d7z6[1] = Ky4oz6;
assign O977z6 = (!O15oz6);
assign A877z6 = (!R45oz6);
assign W177z6 = (!V75oz6);
assign I077z6 = (!Za5oz6);
assign P6d7z6[1] = Ce5oz6;
assign Abh7v6 = (!Fh5oz6);
assign L9d7z6[3] = Jk5oz6;
assign Ea77z6 = (!Nn5oz6);
assign Q877z6 = (!Qq5oz6);
assign M277z6 = (!Ut5oz6);
assign Y077z6 = (!Yw5oz6);
assign P6d7z6[2] = B06oz6;
assign Zec7z6[14] = E36oz6;
assign Uicdt6 = D66oz6;
assign Yfadt6 = A96oz6;
assign Bqbdt6 = Db6oz6;
assign Lpc7z6[1] = Hd6oz6;
assign G597z6 = (!Ig6oz6);
assign Pmc7z6[2] = Jj6oz6;
assign Pmc7z6[1] = Mm6oz6;
assign Ohe7z6[1] = Pp6oz6;
assign L2gdt6 = Rr6oz6;
assign vis_r3_o[5] = Yt6oz6;
assign vis_psp_o[5] = Ow6oz6;
assign Fhc7z6[5] = Fz6oz6;
assign Bdf7z6[3] = O17oz6;
assign Bdf7z6[2] = O47oz6;
assign D5f7z6[3] = O77oz6;
assign D5f7z6[4] = Ka7oz6;
assign Zhbdt6 = Gd7oz6;
assign L9d7z6[5] = Hf7oz6;
assign Pacdt6 = Li7oz6;
assign Bfd7z6[1] = Kl7oz6;
assign Gcd7z6[1] = No7oz6;
assign Byc7z6[19] = Pr7oz6;
assign Zec7z6[3] = Tu7oz6;
assign Byc7z6[3] = Rx7oz6;
assign Zec7z6[19] = U08oz6;
assign Ohe7z6[4] = T38oz6;
assign N0gdt6 = V58oz6;
assign Mfe7z6[4] = X78oz6;
assign Hir8v6 = (!Aa8oz6);
assign Cubdt6 = Sc8oz6;
assign D6c7z6[3] = Sf8oz6;
assign J2cdt6 = Ui8oz6;
assign N1m7z6[4] = Xk8oz6;
assign K6adt6 = Ko8oz6;
assign Ven7z6[1] = Hr8oz6;
assign Tim7z6[9] = Vt8oz6;
assign K377z6 = (!Jw8oz6);
assign U277z6 = (!Mz8oz6);
assign Zec7z6[25] = P29oz6;
assign Byc7z6[25] = O59oz6;
assign Zec7z6[9] = S89oz6;
assign V1c7z6[3] = Qb9oz6;
assign Nnr8v6 = (!Vd9oz6);
assign Kgbdt6 = Ng9oz6;
assign Ke2ft6 = Qj9oz6;
assign H8c7v6 = Ql9oz6;
assign Uib7v6 = Nn9oz6;
assign Rmb7v6 = Up9oz6;
assign Jezmz6[7] = Zr9oz6;
assign Fed7v6 = Gu9oz6;
assign Ft0nz6[4] = Gw9oz6;
assign Ft0nz6[1] = Gy9oz6;
assign Ft0nz6[0] = G0aoz6;
assign Ei67z6 = G2aoz6;
assign Au1nz6[2] = B4aoz6;
assign Zs1nz6[2] = Z5aoz6;
assign Ohe7z6[3] = X7aoz6;
assign Wui7z6[26] = Z9aoz6;
assign Qmb7z6[2] = Bcaoz6;
assign Nob7z6[2] = Xeaoz6;
assign G5j7z6[48] = Chaoz6;
assign M6j7z6[48] = Bkaoz6;
assign Qmb7z6[8] = Anaoz6;
assign Nob7z6[8] = Wpaoz6;
assign G5j7z6[60] = Bsaoz6;
assign M6j7z6[60] = Avaoz6;
assign Itb7z6[28] = Zxaoz6;
assign Tim7z6[28] = R0boz6;
assign K777z6 = (!G3boz6);
assign U677z6 = (!K6boz6);
assign Zec7z6[12] = O9boz6;
assign Byc7z6[12] = Ncboz6;
assign Zec7z6[28] = Rfboz6;
assign Ecc7z6[12] = Qiboz6;
assign Dzget6 = Plboz6;
assign Senet6 = Foboz6;
assign Oe2et6 = Zqboz6;
assign Ldbdt6 = Qtboz6;
assign Ihnet6 = Jwboz6;
assign Ifo7v6 = (!Wyboz6);
assign Byi7z6[30] = Y1coz6;
assign Itb7z6[30] = Y3coz6;
assign Coxmz6[30] = Q6coz6;
assign L5ymz6[33] = L8coz6;
assign L5ymz6[32] = Eacoz6;
assign L5ymz6[31] = Xbcoz6;
assign L5ymz6[30] = Qdcoz6;
assign L5ymz6[29] = Jfcoz6;
assign L5ymz6[28] = Chcoz6;
assign L5ymz6[27] = Vicoz6;
assign L5ymz6[26] = Okcoz6;
assign L5ymz6[25] = Hmcoz6;
assign Tfxmz6[10] = Aocoz6;
assign Hnxmz6[10] = Cqcoz6;
assign Njxmz6[10] = Xrcoz6;
assign Ab57v6 = Aucoz6;
assign Hf57v6 = Pvcoz6;
assign Ii57v6 = Fxcoz6;
assign Tq57v6 = Vycoz6;
assign SWDOEN = J0doz6;
assign Ifh7v6 = (!J0doz6);
assign B1ymz6[0] = X1doz6;
assign B1ymz6[1] = T3doz6;
assign B1ymz6[2] = P5doz6;
assign B1ymz6[3] = L7doz6;
assign B1ymz6[4] = H9doz6;
assign B1ymz6[5] = Dbdoz6;
assign Fqxmz6[5] = Zcdoz6;
assign Fqxmz6[3] = Vedoz6;
assign Fqxmz6[2] = Rgdoz6;
assign Fqxmz6[1] = Nidoz6;
assign Fqxmz6[4] = Jkdoz6;
assign Fqxmz6[0] = Fmdoz6;
assign R9ymz6[2] = Bodoz6;
assign R9ymz6[0] = Updoz6;
assign R9ymz6[3] = Nrdoz6;
assign R9ymz6[1] = Gtdoz6;
assign nTDOEN = (!Zudoz6);
assign G8ymz6[3] = Nwdoz6;
assign G8ymz6[2] = Fydoz6;
assign G8ymz6[1] = Xzdoz6;
assign G8ymz6[0] = P1eoz6;
assign W6ymz6[0] = H3eoz6;
assign W6ymz6[1] = Y4eoz6;
assign W6ymz6[2] = P6eoz6;
assign W6ymz6[3] = G8eoz6;
assign V357v6 = X9eoz6;
assign Ud57v6 = Nbeoz6;
assign Cxxmz6[7] = Edeoz6;
assign Omxmz6[7] = Veeoz6;
assign U3o7z6[11] = Ngeoz6;
assign Coxmz6[11] = Djeoz6;
assign L5ymz6[14] = Ykeoz6;
assign L5ymz6[13] = Rmeoz6;
assign L5ymz6[12] = Koeoz6;
assign L5ymz6[11] = Dqeoz6;
assign L5ymz6[10] = Wreoz6;
assign L5ymz6[9] = Pteoz6;
assign L5ymz6[8] = Hveoz6;
assign L5ymz6[7] = Zweoz6;
assign F267v6 = Ryeoz6;
assign Aixmz6[4] = I0foz6;
assign Aixmz6[5] = M2foz6;
assign Aixmz6[6] = Q4foz6;
assign Aixmz6[7] = U6foz6;
assign Aixmz6[8] = Y8foz6;
assign Aixmz6[9] = Cbfoz6;
assign Aixmz6[10] = Gdfoz6;
assign Aixmz6[11] = Lffoz6;
assign Aixmz6[22] = Qhfoz6;
assign Aixmz6[23] = Vjfoz6;
assign Aixmz6[24] = Amfoz6;
assign Aixmz6[25] = Fofoz6;
assign Aixmz6[26] = Kqfoz6;
assign Aixmz6[27] = Psfoz6;
assign Aixmz6[28] = Uufoz6;
assign Aixmz6[29] = Zwfoz6;
assign Aixmz6[30] = Ezfoz6;
assign Qs67z6 = (!J1goz6);
assign S367v6 = V2goz6;
assign Bmh7v6 = K4goz6;
assign Oh67z6 = (!A6goz6);
assign Ye47v6 = X7goz6;
assign Up47v6 = V9goz6;
assign Un67v6 = Nbgoz6;
assign Ek47v6 = Jdgoz6;
assign Is67z6 = (!Gfgoz6);
assign Wh77z6 = (!Sggoz6);
assign Uu57v6 = Ligoz6;
assign Hw57v6 = Ckgoz6;
assign Ulh7v6 = Rlgoz6;
assign Gh67z6 = (!Jngoz6);
assign Ee47v6 = Ipgoz6;
assign Hnxmz6[0] = Irgoz6;
assign Njxmz6[0] = Ctgoz6;
assign Cxxmz6[12] = Evgoz6;
assign Cxxmz6[11] = Wwgoz6;
assign Ikxmz6[3] = Oygoz6;
assign Dbymz6[1] = P0hoz6;
assign Dbymz6[0] = A2hoz6;
assign Fvzet6 = L3hoz6;
assign F5o7z6[7] = Z5hoz6;
assign Gco7z6[6] = P8hoz6;
assign Io47v6 = Abhoz6;
assign H557v6 = Uchoz6;
assign Pm57v6 = Jehoz6;
assign Cxxmz6[31] = Wfhoz6;
assign Omxmz6[31] = Ohhoz6;
assign Cxxmz6[30] = Cjhoz6;
assign Omxmz6[30] = Ukhoz6;
assign Sl47v6 = Imhoz6;
assign R1adt6 = Dohoz6;
assign A9bdt6 = Sphoz6;
assign D9h7v6 = (!Wqhoz6);
assign Gr67v6 = Urhoz6;
assign Ii47v6 = Sthoz6;
assign L5ymz6[34] = Rvhoz6;
assign Aixmz6[31] = Kxhoz6;
assign U3o7z6[31] = Pzhoz6;
assign Fvb7z6[31] = F2ioz6;
assign C1o7z6[1] = X4ioz6;
assign Vveet6 = W7ioz6;
assign A0fet6 = Faioz6;
assign Qteet6 = Mcioz6;
assign Y497z6 = (!Veioz6);
assign Qboet6 = Xhioz6;
assign U8oet6 = Xkioz6;
assign Wbxdt6 = Xnioz6;
assign W13et6 = Arioz6;
assign No7et6 = Utioz6;
assign Kih7z6[1] = Twioz6;
assign Kih7z6[0] = Pzioz6;
assign D6c7z6[2] = L2joz6;
assign Yg77z6 = (!N5joz6);
assign Thbet6 = F8joz6;
assign X4eet6 = Fbjoz6;
assign Lcadt6 = Jdjoz6;
assign Ohe7z6[2] = Cgjoz6;
assign vis_psp_o[30] = Eijoz6;
assign vis_psp_o[8] = Wkjoz6;
assign Fhc7z6[8] = Nnjoz6;
assign Fuadt6 = Wpjoz6;
assign Uebdt6 = Yrjoz6;
assign vis_pc_o[31] = Yujoz6;
assign vis_pc_o[1] = Fxjoz6;
assign vis_pc_o[2] = Lzjoz6;
assign vis_pc_o[3] = R1koz6;
assign vis_pc_o[4] = X3koz6;
assign vis_pc_o[5] = D6koz6;
assign vis_pc_o[6] = J8koz6;
assign vis_pc_o[7] = Pakoz6;
assign vis_pc_o[8] = Vckoz6;
assign vis_pc_o[9] = Bfkoz6;
assign vis_pc_o[10] = Hhkoz6;
assign vis_pc_o[11] = Ojkoz6;
assign vis_pc_o[12] = Vlkoz6;
assign vis_pc_o[13] = Cokoz6;
assign vis_pc_o[14] = Jqkoz6;
assign vis_pc_o[15] = Qskoz6;
assign vis_pc_o[16] = Xukoz6;
assign vis_pc_o[17] = Exkoz6;
assign vis_pc_o[18] = Lzkoz6;
assign vis_pc_o[19] = S1loz6;
assign vis_pc_o[20] = Z3loz6;
assign vis_pc_o[21] = G6loz6;
assign vis_pc_o[22] = N8loz6;
assign vis_pc_o[23] = Ualoz6;
assign vis_pc_o[24] = Bdloz6;
assign vis_pc_o[25] = Ifloz6;
assign vis_pc_o[26] = Phloz6;
assign Fhc7z6[26] = Wjloz6;
assign Fth7z6[26] = Gmloz6;
assign Tim7z6[2] = Eploz6;
assign Uu67z6 = (!Srloz6);
assign Eu67z6 = (!Vuloz6);
assign Zec7z6[18] = Yxloz6;
assign Byc7z6[18] = X0moz6;
assign Zec7z6[2] = B4moz6;
assign Pxg7z6[1] = Z6moz6;
assign P4c7z6[1] = W9moz6;
assign Xz7et6 = Tcmoz6;
assign Toi7z6[2] = Ufmoz6;
assign Aqadt6 = Dimoz6;
assign Esadt6 = Kkmoz6;
assign Zjb7z6[9] = Mmmoz6;
assign Dradt6 = Gpmoz6;
assign O6cet6 = Krmoz6;
assign O9adt6 = Ptmoz6;
assign P8adt6 = Tvmoz6;
assign Frzet6 = Wxmoz6;
assign Oeo7z6[2] = J0noz6;
assign R0bdt6 = W2noz6;
assign Cp47v6 = G5noz6;
assign S657v6 = Y6noz6;
assign Cxxmz6[4] = N8noz6;
assign Omxmz6[4] = Eanoz6;
assign F5o7z6[4] = Wbnoz6;
assign Ugo7z6[1] = Menoz6;
assign Itb7z6[17] = Dhnoz6;
assign Tim7z6[17] = Vjnoz6;
assign Wt67z6 = (!Kmnoz6);
assign Gt67z6 = (!Opnoz6);
assign Zec7z6[1] = Ssnoz6;
assign Byc7z6[1] = Qvnoz6;
assign Zec7z6[17] = Tynoz6;
assign Qyddt6 = S1ooz6;
assign Y3fet6 = S3ooz6;
assign Geddt6 = R5ooz6;
assign Edh7z6[1] = O8ooz6;
assign S7n7z6[1] = Kbooz6;
assign Tim7z6[29] = Deooz6;
assign Itb7z6[29] = Sgooz6;
assign Coxmz6[29] = Kjooz6;
assign Cxxmz6[29] = Flooz6;
assign Cxxmz6[28] = Xmooz6;
assign Omxmz6[28] = Poooz6;
assign Qm47v6 = Dqooz6;
assign Lc57v6 = Yrooz6;
assign M257v6 = Ltooz6;
assign On47v6 = Yuooz6;
assign Coxmz6[0] = Twooz6;
assign Krxmz6[0] = Nyooz6;
assign Cxxmz6[0] = E0poz6;
assign Fy47v6 = V1poz6;
assign Uzxmz6[2] = O3poz6;
assign D857v6 = C5poz6;
assign Krxmz6[29] = U6poz6;
assign Krxmz6[11] = M8poz6;
assign Krxmz6[30] = Eapoz6;
assign Krxmz6[6] = Wbpoz6;
assign Cxxmz6[6] = Ndpoz6;
assign Omxmz6[6] = Efpoz6;
assign F5o7z6[6] = Wgpoz6;
assign Oeo7z6[0] = Mjpoz6;
assign Blzet6 = Zlpoz6;
assign T21ft6 = Nopoz6;
assign Hgzet6 = Drpoz6;
assign Dnh7v6 = (!Ntpoz6);
assign F51ft6 = Fwpoz6;
assign Zdh7v6 = (!Yypoz6);
assign L3bdt6 = L1qoz6;
assign Fvb7z6[11] = A4qoz6;
assign Ugo7z6[0] = S6qoz6;
assign Itb7z6[1] = J9qoz6;
assign Coxmz6[1] = Bcqoz6;
assign Krxmz6[1] = Vdqoz6;
assign Cxxmz6[1] = Mfqoz6;
assign Ulxmz6[1] = Dhqoz6;
assign Pl0ft6 = Fjqoz6;
assign Hub7z6[0] = Zlqoz6;
assign U3o7z6[10] = Qoqoz6;
assign Fvb7z6[10] = Grqoz6;
assign Coxmz6[10] = Ytqoz6;
assign Krxmz6[10] = Tvqoz6;
assign Cxxmz6[10] = Lxqoz6;
assign Cxxmz6[9] = Dzqoz6;
assign Fuxmz6[1] = U0roz6;
assign Uzxmz6[4] = K2roz6;
assign Uzxmz6[3] = Y3roz6;
assign Uzxmz6[0] = M5roz6;
assign Uzxmz6[1] = A7roz6;
assign Cl57v6 = O8roz6;
assign Yn57v6 = Earoz6;
assign Ovxmz6[0] = Ubroz6;
assign Ds57v6 = Pdroz6;
assign Kp57v6 = Bfroz6;
assign Tg57v6 = Ogroz6;
assign Yg67z6 = (!Hiroz6);
assign Ulxmz6[4] = Ujroz6;
assign Ulxmz6[6] = Wlroz6;
assign Ulxmz6[7] = Ynroz6;
assign Ulxmz6[9] = Aqroz6;
assign Ulxmz6[10] = Csroz6;
assign Ulxmz6[11] = Furoz6;
assign Ulxmz6[12] = Iwroz6;
assign Ulxmz6[28] = Lyroz6;
assign U3o7z6[28] = O0soz6;
assign Fvb7z6[28] = E3soz6;
assign Ulxmz6[29] = W5soz6;
assign U3o7z6[29] = Z7soz6;
assign Fvb7z6[29] = Pasoz6;
assign Ulxmz6[30] = Hdsoz6;
assign U3o7z6[30] = Kfsoz6;
assign Fvb7z6[30] = Aisoz6;
assign Ulxmz6[31] = Sksoz6;
assign Ulxmz6[0] = Vmsoz6;
assign Usxmz6[0] = Xosoz6;
assign Usxmz6[1] = Pqsoz6;
assign E157v6 = Hssoz6;
assign Yt47v6 = Ttsoz6;
assign Cxxmz6[2] = Ivsoz6;
assign Ulxmz6[2] = Zwsoz6;
assign Blxmz6[0] = Bzsoz6;
assign Hnxmz6[11] = E1toz6;
assign Njxmz6[11] = Z2toz6;
assign Cxxmz6[23] = C5toz6;
assign Ulxmz6[23] = U6toz6;
assign U3o7z6[23] = X8toz6;
assign Fvb7z6[23] = Nbtoz6;
assign Cxxmz6[22] = Fetoz6;
assign Ulxmz6[22] = Xftoz6;
assign U3o7z6[22] = Aitoz6;
assign Fvb7z6[22] = Qktoz6;
assign Cxxmz6[21] = Odazz6;
assign Ulxmz6[21] = Gfazz6;
assign Njxmz6[9] = Jhazz6;
assign Hnxmz6[9] = Ljazz6;
assign Tfxmz6[9] = Flazz6;
assign L5ymz6[24] = Gnazz6;
assign Aixmz6[21] = Zoazz6;
assign U3o7z6[21] = Erazz6;
assign Fvb7z6[21] = Utazz6;
assign L5ymz6[23] = Mwazz6;
assign Aixmz6[20] = Fyazz6;
assign Tfxmz6[8] = K0bzz6;
assign Hnxmz6[8] = L2bzz6;
assign Njxmz6[8] = F4bzz6;
assign Cxxmz6[20] = H6bzz6;
assign Ulxmz6[20] = Z7bzz6;
assign U3o7z6[20] = Cabzz6;
assign Fvb7z6[20] = Scbzz6;
assign Cxxmz6[19] = Kfbzz6;
assign Ulxmz6[19] = Chbzz6;
assign Njxmz6[7] = Fjbzz6;
assign Hnxmz6[7] = Hlbzz6;
assign Tfxmz6[7] = Bnbzz6;
assign L5ymz6[22] = Cpbzz6;
assign Aixmz6[19] = Vqbzz6;
assign U3o7z6[19] = Atbzz6;
assign Fvb7z6[19] = Qvbzz6;
assign L5ymz6[21] = Iybzz6;
assign Aixmz6[18] = B0czz6;
assign Tfxmz6[6] = G2czz6;
assign Hnxmz6[6] = H4czz6;
assign Njxmz6[6] = B6czz6;
assign Cxxmz6[18] = D8czz6;
assign Ulxmz6[18] = V9czz6;
assign U3o7z6[18] = Ybczz6;
assign Fvb7z6[18] = Oeczz6;
assign Cxxmz6[17] = Ghczz6;
assign Ulxmz6[17] = Yiczz6;
assign Njxmz6[5] = Blczz6;
assign Hnxmz6[5] = Dnczz6;
assign Tfxmz6[5] = Xoczz6;
assign L5ymz6[20] = Yqczz6;
assign Aixmz6[17] = Rsczz6;
assign U3o7z6[17] = Wuczz6;
assign Fvb7z6[17] = Mxczz6;
assign L5ymz6[19] = E0dzz6;
assign Aixmz6[16] = X1dzz6;
assign Tfxmz6[4] = C4dzz6;
assign Hnxmz6[4] = D6dzz6;
assign Njxmz6[4] = X7dzz6;
assign Cxxmz6[16] = Z9dzz6;
assign Ulxmz6[16] = Rbdzz6;
assign U3o7z6[16] = Uddzz6;
assign Fvb7z6[16] = Kgdzz6;
assign Cxxmz6[15] = Cjdzz6;
assign Ulxmz6[15] = Ukdzz6;
assign Njxmz6[3] = Xmdzz6;
assign Hnxmz6[3] = Zodzz6;
assign Tfxmz6[3] = Tqdzz6;
assign L5ymz6[18] = Usdzz6;
assign Aixmz6[15] = Nudzz6;
assign U3o7z6[15] = Swdzz6;
assign Fvb7z6[15] = Izdzz6;
assign L5ymz6[17] = A2ezz6;
assign Aixmz6[14] = T3ezz6;
assign Tfxmz6[2] = Y5ezz6;
assign Hnxmz6[2] = Z7ezz6;
assign Njxmz6[2] = T9ezz6;
assign Cxxmz6[14] = Vbezz6;
assign Ulxmz6[14] = Ndezz6;
assign U3o7z6[14] = Qfezz6;
assign Fvb7z6[14] = Giezz6;
assign Cxxmz6[13] = Ykezz6;
assign Ulxmz6[13] = Qmezz6;
assign Njxmz6[1] = Toezz6;
assign Hnxmz6[1] = Vqezz6;
assign Tfxmz6[1] = Psezz6;
assign L5ymz6[16] = Quezz6;
assign Aixmz6[13] = Jwezz6;
assign U3o7z6[13] = Oyezz6;
assign Fvb7z6[13] = E1fzz6;
assign L5ymz6[15] = W3fzz6;
assign Aixmz6[12] = P5fzz6;
assign U3o7z6[12] = U7fzz6;
assign Fvb7z6[12] = Kafzz6;
assign Klo7z6[0] = Cdfzz6;
assign Q497z6 = (!Yefzz6);
assign Lq0ft6 = Vhfzz6;
assign Ejo7z6[0] = Pkfzz6;
assign Ejo7z6[1] = Cnfzz6;
assign Xczet6 = Ppfzz6;
assign U71ft6 = Dsfzz6;
assign Ua77z6 = (!Wufzz6);
assign Ma77z6 = (!Jxfzz6);
assign K4bdt6 = Xzfzz6;
assign O3uet6 = P2gzz6;
assign I2yet6 = P5gzz6;
assign Rnm7z6[2] = D8gzz6;
assign Rnm7z6[1] = Dbgzz6;
assign Rnm7z6[0] = Degzz6;
assign I497z6 = (!Dhgzz6);
assign Dkm7z6[0] = Dkgzz6;
assign Knh7v6 = (!Cngzz6);
assign Qln7z6[1] = Wpgzz6;
assign Ygo7v6 = (!Msgzz6);
assign X0oet6 = Jvgzz6;
assign Meoet6 = Bygzz6;
assign Kqm7z6[0] = D1hzz6;
assign Kqm7z6[1] = D4hzz6;
assign Sz67z6 = (!D7hzz6);
assign Cz67z6 = (!Gahzz6);
assign Zec7z6[22] = Jdhzz6;
assign Byc7z6[22] = Ighzz6;
assign Zec7z6[6] = Mjhzz6;
assign I0c7z6[0] = Kmhzz6;
assign Edh7z6[0] = Tohzz6;
assign Ven7z6[0] = Prhzz6;
assign Tim7z6[3] = Duhzz6;
assign Itb7z6[3] = Rwhzz6;
assign Coxmz6[3] = Jzhzz6;
assign Krxmz6[3] = D1izz6;
assign Cxxmz6[3] = U2izz6;
assign Ulxmz6[3] = L4izz6;
assign Blxmz6[1] = N6izz6;
assign Omxmz6[3] = Q8izz6;
assign Omxmz6[2] = Haizz6;
assign R957v6 = Ybizz6;
assign L5ymz6[6] = Ldizz6;
assign Aixmz6[3] = Dfizz6;
assign L5ymz6[5] = Hhizz6;
assign Aixmz6[2] = Ziizz6;
assign L5ymz6[4] = Dlizz6;
assign Aixmz6[1] = Vmizz6;
assign L5ymz6[3] = Zoizz6;
assign Aixmz6[0] = Rqizz6;
assign L5ymz6[2] = Vsizz6;
assign Uixmz6[3] = Nuizz6;
assign F5o7z6[3] = Ewizz6;
assign L5ymz6[1] = Uyizz6;
assign Uixmz6[2] = M0jzz6;
assign Cozet6 = D2jzz6;
assign Zn0ft6 = X4jzz6;
assign K6uet6 = N7jzz6;
assign O7o7z6[2] = Fajzz6;
assign Oeo7z6[1] = Zcjzz6;
assign Ppzet6 = Mfjzz6;
assign Ov0ft6 = Bijzz6;
assign L1bdt6 = Rkjzz6;
assign Ekoet6 = Bnjzz6;
assign Xnnet6 = Xpjzz6;
assign Styet6 = Osjzz6;
assign Znn7z6[0] = Fvjzz6;
assign Tszet6 = Rxjzz6;
assign Hub7z6[1] = H0kzz6;
assign F5o7z6[2] = Y2kzz6;
assign L5ymz6[0] = O5kzz6;
assign Hhxmz6[0] = G7kzz6;
assign Hhxmz6[1] = I9kzz6;
assign Ogxmz6[0] = Kbkzz6;
assign Ogxmz6[1] = Ndkzz6;
assign Ogxmz6[2] = Qfkzz6;
assign Ogxmz6[3] = Thkzz6;
assign Qf47v6 = Wjkzz6;
assign Mg47v6 = Plkzz6;
assign Kh47v6 = Knkzz6;
assign Ez57v6 = Fpkzz6;
assign Tfxmz6[11] = Xqkzz6;
assign S067v6 = Zskzz6;
assign Uixmz6[25] = Qukzz6;
assign Uixmz6[26] = Gwkzz6;
assign Uixmz6[27] = Wxkzz6;
assign Uixmz6[28] = Mzkzz6;
assign Uixmz6[29] = C1lzz6;
assign Uixmz6[30] = S2lzz6;
assign Uixmz6[31] = I4lzz6;
assign Uixmz6[4] = Y5lzz6;
assign Uixmz6[5] = S7lzz6;
assign F5o7z6[5] = M9lzz6;
assign Coxmz6[17] = Cclzz6;
assign Krxmz6[17] = Xdlzz6;
assign Coxmz6[28] = Pflzz6;
assign Krxmz6[28] = Khlzz6;
assign Coxmz6[25] = Cjlzz6;
assign Krxmz6[25] = Xklzz6;
assign Cxxmz6[25] = Pmlzz6;
assign Ulxmz6[25] = Holzz6;
assign U3o7z6[25] = Kqlzz6;
assign Fvb7z6[25] = Atlzz6;
assign Ven7z6[2] = Svlzz6;
assign Znn7z6[2] = Gylzz6;
assign Gmnet6 = S0mzz6;
assign Aym7z6[1] = L3mzz6;
assign Aym7z6[2] = B6mzz6;
assign Aym7z6[3] = R8mzz6;
assign Sjyet6 = Hbmzz6;
assign Znn7z6[3] = Wdmzz6;
assign Ueh7v6 = (!Igmzz6);
assign G977z6 = (!Mjmzz6);
assign Gazet6 = Qmmzz6;
assign Kyn7z6[1] = Lpmzz6;
assign Kyn7z6[0] = Ksmzz6;
assign Kyn7z6[2] = Jvmzz6;
assign D6c7z6[0] = Iymzz6;
assign Ewyet6 = K1nzz6;
assign Dtm7z6[3] = B4nzz6;
assign Dtm7z6[1] = V6nzz6;
assign Dtm7z6[0] = P9nzz6;
assign Dtm7z6[2] = Jcnzz6;
assign Itb7z6[2] = Dfnzz6;
assign Itb7z6[9] = Vhnzz6;
assign Tim7z6[25] = Nknzz6;
assign Itb7z6[25] = Cnnzz6;
assign S377z6 = (!Upnzz6);
assign C377z6 = (!Ysnzz6);
assign Tim7z6[27] = Cwnzz6;
assign Itb7z6[27] = Rynzz6;
assign Coxmz6[27] = J1ozz6;
assign Krxmz6[27] = E3ozz6;
assign Cxxmz6[27] = W4ozz6;
assign Ulxmz6[27] = O6ozz6;
assign U3o7z6[27] = R8ozz6;
assign Fvb7z6[27] = Hbozz6;
assign Cxxmz6[26] = Zdozz6;
assign Ulxmz6[26] = Rfozz6;
assign Itb7z6[26] = Uhozz6;
assign Tim7z6[26] = Mkozz6;
assign Y477z6 = (!Bnozz6);
assign I477z6 = (!Fqozz6);
assign U3o7z6[26] = Jtozz6;
assign Fvb7z6[26] = Zvozz6;
assign Coxmz6[26] = Ryozz6;
assign Krxmz6[26] = M0pzz6;
assign Omxmz6[26] = E2pzz6;
assign Wk47v6 = S3pzz6;
assign Omxmz6[27] = L5pzz6;
assign E677z6 = (!Z6pzz6);
assign O577z6 = (!Dapzz6);
assign Tim7z6[4] = Hdpzz6;
assign Itb7z6[4] = Vfpzz6;
assign Gx67z6 = (!Nipzz6);
assign Qw67z6 = (!Qlpzz6);
assign Tim7z6[5] = Topzz6;
assign Itb7z6[5] = Hrpzz6;
assign Coxmz6[5] = Ztpzz6;
assign Krxmz6[5] = Tvpzz6;
assign Cxxmz6[5] = Kxpzz6;
assign Ulxmz6[5] = Bzpzz6;
assign Gco7z6[5] = D1qzz6;
assign Gco7z6[4] = A4qzz6;
assign U3o7z6[9] = X6qzz6;
assign Fvb7z6[9] = M9qzz6;
assign Coxmz6[9] = Dcqzz6;
assign Krxmz6[9] = Xdqzz6;
assign U3o7z6[8] = Ofqzz6;
assign Fvb7z6[8] = Diqzz6;
assign Coxmz6[8] = Ukqzz6;
assign Krxmz6[8] = Omqzz6;
assign Cxxmz6[8] = Foqzz6;
assign Ulxmz6[8] = Wpqzz6;
assign Itb7z6[8] = Yrqzz6;
assign Fuxmz6[0] = Quqzz6;
assign Ikxmz6[0] = Gwqzz6;
assign U3o7z6[7] = Hyqzz6;
assign Fvb7z6[7] = W0rzz6;
assign U3o7z6[6] = N3rzz6;
assign Fvb7z6[6] = C6rzz6;
assign U3o7z6[5] = T8rzz6;
assign Fvb7z6[5] = Ibrzz6;
assign U3o7z6[4] = Zdrzz6;
assign Fvb7z6[4] = Ogrzz6;
assign Klo7z6[6] = Fjrzz6;
assign Klo7z6[4] = Blrzz6;
assign Klo7z6[5] = Xmrzz6;
assign Klo7z6[3] = Torzz6;
assign Klo7z6[2] = Pqrzz6;
assign Klo7z6[1] = Lsrzz6;
assign Coxmz6[4] = Hurzz6;
assign Krxmz6[4] = Bwrzz6;
assign Y9o7z6[3] = Sxrzz6;
assign Fvb7z6[3] = H0szz6;
assign Y9o7z6[2] = Y2szz6;
assign Coxmz6[2] = N5szz6;
assign Krxmz6[2] = H7szz6;
assign Fvb7z6[2] = Y8szz6;
assign Y9o7z6[1] = Pbszz6;
assign Y9o7z6[0] = Eeszz6;
assign Bizet6 = Tgszz6;
assign K01ft6 = Ijszz6;
assign Mezet6 = Vlszz6;
assign Wmh7v6 = (!Coszz6);
assign Omxmz6[5] = Vqszz6;
assign My67z6 = (!Nsszz6);
assign Wx67z6 = (!Qvszz6);
assign Tim7z6[6] = Tyszz6;
assign Itb7z6[6] = H1tzz6;
assign Coxmz6[6] = Z3tzz6;
assign Tim7z6[7] = T5tzz6;
assign Itb7z6[7] = H8tzz6;
assign Coxmz6[7] = Zatzz6;
assign Krxmz6[7] = Tctzz6;
assign Qmzet6 = Ketzz6;
assign K2bdt6 = Dhtzz6;
assign Pjb7z6[3] = Sjtzz6;
assign Pjb7z6[4] = Oltzz6;
assign Pjb7z6[6] = Kntzz6;
assign Pjb7z6[7] = Gptzz6;
assign Pjb7z6[9] = Crtzz6;
assign Pjb7z6[13] = Ystzz6;
assign Pjb7z6[14] = Vutzz6;
assign Pjb7z6[15] = Swtzz6;
assign Pjb7z6[16] = Pytzz6;
assign Pjb7z6[17] = M0uzz6;
assign Pjb7z6[5] = J2uzz6;
assign Pjb7z6[8] = F4uzz6;
assign Pjb7z6[10] = B6uzz6;
assign Pjb7z6[11] = Y7uzz6;
assign Pjb7z6[18] = V9uzz6;
assign Pjb7z6[19] = Sbuzz6;
assign D16ft6 = Pduzz6;
assign K2adt6 = Ofuzz6;
assign A497z6 = (!Jhuzz6);
assign Omxmz6[25] = Hjuzz6;
assign Coxmz6[24] = Vkuzz6;
assign Krxmz6[24] = Qmuzz6;
assign Cxxmz6[24] = Iouzz6;
assign Ulxmz6[24] = Aquzz6;
assign Itb7z6[24] = Dsuzz6;
assign U3o7z6[24] = Vuuzz6;
assign Fvb7z6[24] = Lxuzz6;
assign S397z6 = (!D0vzz6);
assign Uixmz6[6] = R1vzz6;
assign Uixmz6[7] = L3vzz6;
assign Uixmz6[24] = F5vzz6;
assign Oh77z6 = (!V6vzz6);
assign Q2ymz6[1] = S8vzz6;
assign Q2ymz6[0] = Iavzz6;
assign Sx57v6 = Ybvzz6;
assign Aw67z6 = (!Odvzz6);
assign Kv67z6 = (!Rgvzz6);
assign Itb7z6[10] = Ujvzz6;
assign Tim7z6[10] = Mmvzz6;
assign Q477z6 = (!Bpvzz6);
assign A477z6 = (!Fsvzz6);
assign Itb7z6[11] = Jvvzz6;
assign Tim7z6[11] = Byvzz6;
assign W577z6 = (!Q0wzz6);
assign G577z6 = (!U3wzz6);
assign Zec7z6[27] = Y6wzz6;
assign Byc7z6[27] = X9wzz6;
assign Zec7z6[11] = Bdwzz6;
assign Qwddt6 = Agwzz6;
assign K397z6 = (!Eiwzz6);
assign Lpc7z6[0] = Ikwzz6;
assign Bfd7z6[3] = Jnwzz6;
assign Gcd7z6[3] = Mqwzz6;
assign Bfd7z6[5] = Otwzz6;
assign Gcd7z6[5] = Rwwzz6;
assign Bfd7z6[0] = Tzwzz6;
assign Gcd7z6[0] = W2xzz6;
assign Bfd7z6[2] = Y5xzz6;
assign Bfd7z6[4] = B9xzz6;
assign Gcd7z6[4] = Ecxzz6;
assign Gcd7z6[2] = Gfxzz6;
assign Zec7z6[26] = Iixzz6;
assign Byc7z6[26] = Hlxzz6;
assign Zec7z6[10] = Loxzz6;
assign F4edt6 = Krxzz6;
assign Jqj7z6[5] = Ktxzz6;
assign Xsddt6 = Lwxzz6;
assign Geh7v6 = (!Lyxzz6);
assign Ffadt6 = M0yzz6;
assign Tuddt6 = N2yzz6;
assign S6cdt6 = O4yzz6;
assign Uobdt6 = Q6yzz6;
assign M5e7z6[1] = Q8yzz6;
assign Knbdt6 = Vayzz6;
assign W9c7v6 = Ycyzz6;
assign N6c7v6 = Weyzz6;
assign Byc7z6[10] = Ygyzz6;
assign Pmc7z6[0] = Ckyzz6;
assign I5cdt6 = Fnyzz6;
assign K7e7z6[1] = Ipyzz6;
assign B6edt6 = Nryzz6;
assign T3cdt6 = Ptyzz6;
assign Xnh7z6[1] = Xvyzz6;
assign Xnh7z6[0] = Uyyzz6;
assign Byc7z6[11] = R1zzz6;
assign Itb7z6[12] = V4zzz6;
assign Tim7z6[12] = N7zzz6;
assign C777z6 = (!Cazzz6);
assign M677z6 = (!Gdzzz6);
assign Itb7z6[13] = Kgzzz6;
assign Coxmz6[13] = Cjzzz6;
assign Krxmz6[13] = Xkzzz6;
assign Tim7z6[13] = Pmzzz6;
assign I877z6 = (!Epzzz6);
assign S777z6 = (!Iszzz6);
assign Itb7z6[14] = Mvzzz6;
assign Coxmz6[14] = Eyzzz6;
assign Krxmz6[14] = Zzzzz6;
assign Tim7z6[14] = R10007;
assign Byc7z6[14] = G40007;
assign Bfh7v6 = (!K70007);
assign Y877z6 = (!Oa0007);
assign Zec7z6[30] = Sd0007;
assign Ide7z6[0] = Rg0007;
assign Ide7z6[3] = Cj0007;
assign Ide7z6[2] = Nl0007;
assign Ide7z6[1] = Yn0007;
assign K7e7z6[0] = Jq0007;
assign vis_r3_o[3] = Os0007;
assign vis_r3_o[6] = Ev0007;
assign vis_r3_o[7] = Ux0007;
assign vis_r3_o[9] = K01007;
assign vis_psp_o[9] = A31007;
assign vis_r3_o[12] = R51007;
assign vis_psp_o[12] = I81007;
assign vis_r3_o[13] = Ab1007;
assign vis_psp_o[13] = Rd1007;
assign vis_r3_o[14] = Jg1007;
assign vis_psp_o[14] = Aj1007;
assign vis_r3_o[16] = Sl1007;
assign vis_psp_o[16] = Jo1007;
assign vis_r3_o[17] = Br1007;
assign vis_psp_o[17] = St1007;
assign vis_r3_o[19] = Kw1007;
assign vis_psp_o[19] = Bz1007;
assign vis_r3_o[20] = T12007;
assign vis_psp_o[20] = K42007;
assign vis_r3_o[21] = C72007;
assign vis_psp_o[21] = T92007;
assign vis_r3_o[22] = Lc2007;
assign vis_psp_o[22] = Cf2007;
assign vis_r3_o[23] = Uh2007;
assign vis_psp_o[23] = Lk2007;
assign vis_r3_o[24] = Dn2007;
assign vis_psp_o[24] = Up2007;
assign vis_r3_o[25] = Ms2007;
assign vis_psp_o[25] = Dv2007;
assign vis_r3_o[10] = Vx2007;
assign vis_psp_o[10] = M03007;
assign vis_r3_o[18] = E33007;
assign vis_psp_o[18] = V53007;
assign vis_r3_o[26] = N83007;
assign vis_psp_o[26] = Eb3007;
assign vis_r3_o[4] = Wd3007;
assign vis_r3_o[2] = Mg3007;
assign vis_psp_o[2] = Cj3007;
assign vis_r3_o[8] = Tl3007;
assign vis_r3_o[27] = Jo3007;
assign vis_psp_o[27] = Ar3007;
assign vis_r3_o[15] = St3007;
assign vis_psp_o[15] = Jw3007;
assign vis_r3_o[29] = Bz3007;
assign vis_psp_o[29] = S14007;
assign vis_r3_o[28] = K44007;
assign vis_psp_o[28] = B74007;
assign vis_r1_o[0] = T94007;
assign vis_r1_o[30] = Jc4007;
assign vis_r1_o[29] = Af4007;
assign vis_r1_o[28] = Rh4007;
assign vis_r1_o[27] = Ik4007;
assign vis_r1_o[26] = Zm4007;
assign vis_r1_o[25] = Qp4007;
assign vis_r1_o[24] = Hs4007;
assign vis_r1_o[23] = Yu4007;
assign vis_r1_o[22] = Px4007;
assign vis_r1_o[21] = G05007;
assign vis_r1_o[20] = X25007;
assign vis_r1_o[19] = O55007;
assign vis_r1_o[18] = F85007;
assign vis_r1_o[17] = Wa5007;
assign vis_r1_o[16] = Nd5007;
assign vis_r1_o[15] = Eg5007;
assign vis_r1_o[14] = Vi5007;
assign vis_r1_o[13] = Ml5007;
assign vis_r1_o[12] = Do5007;
assign vis_r1_o[11] = Uq5007;
assign vis_r1_o[10] = Lt5007;
assign vis_r1_o[9] = Cw5007;
assign vis_r1_o[8] = Sy5007;
assign vis_r1_o[7] = I16007;
assign vis_r1_o[6] = Y36007;
assign vis_r1_o[5] = O66007;
assign vis_r1_o[4] = E96007;
assign vis_r1_o[3] = Ub6007;
assign vis_r1_o[2] = Ke6007;
assign vis_r1_o[1] = Ah6007;
assign vis_r5_o[0] = Qj6007;
assign vis_r5_o[30] = Gm6007;
assign vis_r5_o[29] = Xo6007;
assign vis_r5_o[28] = Or6007;
assign vis_r5_o[27] = Fu6007;
assign vis_r5_o[26] = Ww6007;
assign vis_r5_o[25] = Nz6007;
assign vis_r5_o[24] = E27007;
assign vis_r5_o[23] = V47007;
assign vis_r5_o[22] = M77007;
assign vis_r5_o[21] = Da7007;
assign vis_r5_o[20] = Uc7007;
assign vis_r5_o[19] = Lf7007;
assign vis_r5_o[18] = Ci7007;
assign vis_r5_o[17] = Tk7007;
assign vis_r5_o[16] = Kn7007;
assign vis_r5_o[15] = Bq7007;
assign vis_r5_o[14] = Ss7007;
assign vis_r5_o[13] = Jv7007;
assign vis_r5_o[12] = Ay7007;
assign vis_r5_o[11] = R08007;
assign vis_r5_o[10] = I38007;
assign vis_r5_o[9] = Z58007;
assign vis_r5_o[8] = P88007;
assign vis_r5_o[7] = Fb8007;
assign vis_r5_o[6] = Vd8007;
assign vis_r5_o[5] = Lg8007;
assign vis_r5_o[4] = Bj8007;
assign vis_r5_o[3] = Rl8007;
assign vis_r5_o[2] = Ho8007;
assign vis_r5_o[1] = Xq8007;
assign vis_r7_o[0] = Nt8007;
assign vis_r7_o[30] = Dw8007;
assign vis_r7_o[29] = Uy8007;
assign vis_r7_o[28] = L19007;
assign vis_r7_o[27] = C49007;
assign vis_r7_o[26] = T69007;
assign vis_r7_o[25] = K99007;
assign vis_r7_o[24] = Bc9007;
assign vis_r7_o[23] = Se9007;
assign vis_r7_o[22] = Jh9007;
assign vis_r7_o[21] = Ak9007;
assign vis_r7_o[20] = Rm9007;
assign vis_r7_o[19] = Ip9007;
assign vis_r7_o[18] = Zr9007;
assign vis_r7_o[17] = Qu9007;
assign vis_r7_o[16] = Hx9007;
assign vis_r7_o[15] = Yz9007;
assign vis_r7_o[14] = P2a007;
assign vis_r7_o[13] = G5a007;
assign vis_r7_o[12] = X7a007;
assign vis_r7_o[11] = Oaa007;
assign vis_r7_o[10] = Fda007;
assign vis_r7_o[9] = Wfa007;
assign vis_r7_o[8] = Mia007;
assign vis_r7_o[7] = Cla007;
assign vis_r7_o[6] = Sna007;
assign vis_r7_o[5] = Iqa007;
assign vis_r7_o[4] = Ysa007;
assign vis_r7_o[3] = Ova007;
assign vis_r7_o[2] = Eya007;
assign vis_r7_o[1] = U0b007;
assign vis_r8_o[0] = K3b007;
assign vis_r8_o[30] = A6b007;
assign vis_r8_o[29] = R8b007;
assign vis_r8_o[28] = Ibb007;
assign vis_r8_o[27] = Zdb007;
assign vis_r8_o[26] = Qgb007;
assign vis_r8_o[25] = Hjb007;
assign vis_r8_o[24] = Ylb007;
assign vis_r8_o[23] = Pob007;
assign vis_r8_o[22] = Grb007;
assign vis_r8_o[21] = Xtb007;
assign vis_r8_o[20] = Owb007;
assign vis_r8_o[19] = Fzb007;
assign vis_r8_o[18] = W1c007;
assign vis_r8_o[17] = N4c007;
assign vis_r8_o[16] = E7c007;
assign vis_r8_o[15] = V9c007;
assign vis_r8_o[14] = Mcc007;
assign vis_r8_o[13] = Dfc007;
assign vis_r8_o[12] = Uhc007;
assign vis_r8_o[11] = Lkc007;
assign vis_r8_o[10] = Cnc007;
assign vis_r8_o[9] = Tpc007;
assign vis_r8_o[8] = Jsc007;
assign vis_r8_o[7] = Zuc007;
assign vis_r8_o[6] = Pxc007;
assign vis_r8_o[5] = F0d007;
assign vis_r8_o[4] = V2d007;
assign vis_r8_o[3] = L5d007;
assign vis_r8_o[2] = B8d007;
assign vis_r8_o[1] = Rad007;
assign vis_r9_o[0] = Hdd007;
assign vis_r9_o[30] = Xfd007;
assign vis_r9_o[29] = Oid007;
assign vis_r9_o[28] = Fld007;
assign vis_r9_o[27] = Wnd007;
assign vis_r9_o[26] = Nqd007;
assign vis_r9_o[25] = Etd007;
assign vis_r9_o[24] = Vvd007;
assign vis_r9_o[23] = Myd007;
assign vis_r9_o[22] = D1e007;
assign vis_r9_o[21] = U3e007;
assign vis_r9_o[20] = L6e007;
assign vis_r9_o[19] = C9e007;
assign vis_r9_o[18] = Tbe007;
assign vis_r9_o[17] = Kee007;
assign vis_r9_o[16] = Bhe007;
assign vis_r9_o[15] = Sje007;
assign vis_r9_o[14] = Jme007;
assign vis_r9_o[13] = Ape007;
assign vis_r9_o[12] = Rre007;
assign vis_r9_o[11] = Iue007;
assign vis_r9_o[10] = Zwe007;
assign vis_r9_o[9] = Qze007;
assign vis_r9_o[8] = G2f007;
assign vis_r9_o[7] = W4f007;
assign vis_r9_o[6] = M7f007;
assign vis_r9_o[5] = Caf007;
assign vis_r9_o[4] = Scf007;
assign vis_r9_o[3] = Iff007;
assign vis_r9_o[2] = Yhf007;
assign vis_r9_o[1] = Okf007;
assign vis_r10_o[0] = Enf007;
assign vis_r10_o[30] = Vpf007;
assign vis_r10_o[29] = Nsf007;
assign vis_r10_o[28] = Fvf007;
assign vis_r10_o[27] = Xxf007;
assign vis_r10_o[26] = P0g007;
assign vis_r10_o[25] = H3g007;
assign vis_r10_o[24] = Z5g007;
assign vis_r10_o[23] = R8g007;
assign vis_r10_o[22] = Jbg007;
assign vis_r10_o[21] = Beg007;
assign vis_r10_o[20] = Tgg007;
assign vis_r10_o[19] = Ljg007;
assign vis_r10_o[18] = Dmg007;
assign vis_r10_o[17] = Vog007;
assign vis_r10_o[16] = Nrg007;
assign vis_r10_o[15] = Fug007;
assign vis_r10_o[14] = Xwg007;
assign vis_r10_o[13] = Pzg007;
assign vis_r10_o[12] = H2h007;
assign vis_r10_o[11] = Z4h007;
assign vis_r10_o[10] = R7h007;
assign vis_r10_o[9] = Jah007;
assign vis_r10_o[8] = Adh007;
assign vis_r10_o[7] = Rfh007;
assign vis_r10_o[6] = Iih007;
assign vis_r10_o[5] = Zkh007;
assign vis_r10_o[4] = Qnh007;
assign vis_r10_o[3] = Hqh007;
assign vis_r10_o[2] = Ysh007;
assign vis_r10_o[1] = Pvh007;
assign vis_r11_o[0] = Gyh007;
assign vis_r11_o[30] = X0i007;
assign vis_r11_o[29] = P3i007;
assign vis_r11_o[28] = H6i007;
assign vis_r11_o[27] = Z8i007;
assign vis_r11_o[26] = Rbi007;
assign vis_r11_o[25] = Jei007;
assign vis_r11_o[24] = Bhi007;
assign vis_r11_o[23] = Tji007;
assign vis_r11_o[22] = Lmi007;
assign vis_r11_o[21] = Dpi007;
assign vis_r11_o[20] = Vri007;
assign vis_r11_o[19] = Nui007;
assign vis_r11_o[18] = Fxi007;
assign vis_r11_o[17] = Xzi007;
assign vis_r11_o[16] = P2j007;
assign vis_r11_o[15] = H5j007;
assign vis_r11_o[14] = Z7j007;
assign vis_r11_o[13] = Raj007;
assign vis_r11_o[12] = Jdj007;
assign vis_r11_o[11] = Bgj007;
assign vis_r11_o[10] = Tij007;
assign vis_r11_o[9] = Llj007;
assign vis_r11_o[8] = Coj007;
assign vis_r11_o[7] = Tqj007;
assign vis_r11_o[6] = Ktj007;
assign vis_r11_o[5] = Bwj007;
assign vis_r11_o[4] = Syj007;
assign vis_r11_o[3] = J1k007;
assign vis_r11_o[2] = A4k007;
assign vis_r11_o[1] = R6k007;
assign vis_r12_o[0] = I9k007;
assign vis_r12_o[30] = Zbk007;
assign vis_r12_o[29] = Rek007;
assign vis_r12_o[28] = Jhk007;
assign vis_r12_o[27] = Bkk007;
assign vis_r12_o[26] = Tmk007;
assign vis_r12_o[25] = Lpk007;
assign vis_r12_o[24] = Dsk007;
assign vis_r12_o[23] = Vuk007;
assign vis_r12_o[22] = Nxk007;
assign vis_r12_o[21] = F0l007;
assign vis_r12_o[20] = X2l007;
assign vis_r12_o[19] = P5l007;
assign vis_r12_o[18] = H8l007;
assign vis_r12_o[17] = Zal007;
assign vis_r12_o[16] = Rdl007;
assign vis_r12_o[15] = Jgl007;
assign vis_r12_o[14] = Bjl007;
assign vis_r12_o[13] = Tll007;
assign vis_r12_o[12] = Lol007;
assign vis_r12_o[11] = Drl007;
assign vis_r12_o[10] = Vtl007;
assign vis_r12_o[9] = Nwl007;
assign vis_r12_o[8] = Ezl007;
assign vis_r12_o[7] = V1m007;
assign vis_r12_o[6] = M4m007;
assign vis_r12_o[5] = D7m007;
assign vis_r12_o[4] = U9m007;
assign vis_r12_o[3] = Lcm007;
assign vis_r12_o[2] = Cfm007;
assign vis_r12_o[1] = Thm007;
assign vis_msp_o[2] = Kkm007;
assign vis_msp_o[30] = Bnm007;
assign vis_msp_o[29] = Tpm007;
assign vis_msp_o[28] = Lsm007;
assign vis_msp_o[27] = Dvm007;
assign vis_msp_o[26] = Vxm007;
assign vis_msp_o[25] = N0n007;
assign vis_msp_o[24] = F3n007;
assign vis_msp_o[23] = X5n007;
assign vis_msp_o[22] = P8n007;
assign vis_msp_o[21] = Hbn007;
assign vis_msp_o[20] = Zdn007;
assign vis_msp_o[19] = Rgn007;
assign vis_msp_o[18] = Jjn007;
assign vis_msp_o[17] = Bmn007;
assign vis_msp_o[16] = Ton007;
assign vis_msp_o[15] = Lrn007;
assign vis_msp_o[14] = Dun007;
assign vis_msp_o[13] = Vwn007;
assign vis_msp_o[12] = Nzn007;
assign vis_msp_o[11] = F2o007;
assign vis_msp_o[10] = X4o007;
assign vis_msp_o[9] = P7o007;
assign vis_msp_o[8] = Gao007;
assign vis_msp_o[7] = Xco007;
assign vis_msp_o[6] = Ofo007;
assign vis_msp_o[5] = Fio007;
assign vis_msp_o[4] = Wko007;
assign vis_msp_o[3] = Nno007;
assign Pic7z6[0] = Eqo007;
assign Pic7z6[30] = Vso007;
assign Pic7z6[29] = Nvo007;
assign Pic7z6[28] = Fyo007;
assign Pic7z6[27] = X0p007;
assign Pic7z6[26] = P3p007;
assign Pic7z6[25] = H6p007;
assign Pic7z6[24] = Z8p007;
assign Pic7z6[23] = Rbp007;
assign Pic7z6[22] = Jep007;
assign Pic7z6[21] = Bhp007;
assign Pic7z6[20] = Tjp007;
assign Pic7z6[19] = Lmp007;
assign Pic7z6[18] = Dpp007;
assign Pic7z6[17] = Vrp007;
assign Pic7z6[16] = Nup007;
assign Pic7z6[15] = Fxp007;
assign Pic7z6[14] = Xzp007;
assign Pic7z6[13] = P2q007;
assign Pic7z6[12] = H5q007;
assign Pic7z6[11] = Z7q007;
assign Pic7z6[10] = Raq007;
assign Pic7z6[9] = Jdq007;
assign Pic7z6[8] = Agq007;
assign Pic7z6[7] = Riq007;
assign Pic7z6[6] = Ilq007;
assign Pic7z6[5] = Znq007;
assign Pic7z6[4] = Qqq007;
assign Pic7z6[3] = Htq007;
assign Pic7z6[2] = Yvq007;
assign Pic7z6[1] = Pyq007;
assign vis_r2_o[0] = G1r007;
assign vis_r2_o[30] = W3r007;
assign vis_r2_o[29] = N6r007;
assign vis_r2_o[28] = E9r007;
assign vis_r2_o[27] = Vbr007;
assign vis_r2_o[26] = Mer007;
assign vis_r2_o[25] = Dhr007;
assign vis_r2_o[24] = Ujr007;
assign vis_r2_o[23] = Lmr007;
assign vis_r2_o[22] = Cpr007;
assign vis_r2_o[21] = Trr007;
assign vis_r2_o[20] = Kur007;
assign vis_r2_o[19] = Bxr007;
assign vis_r2_o[18] = Szr007;
assign vis_r2_o[17] = J2s007;
assign vis_r2_o[16] = A5s007;
assign vis_r2_o[15] = R7s007;
assign vis_r2_o[14] = Ias007;
assign vis_r2_o[13] = Zcs007;
assign vis_r2_o[12] = Qfs007;
assign vis_r2_o[11] = His007;
assign vis_r2_o[10] = Yks007;
assign vis_r2_o[9] = Pns007;
assign vis_r2_o[8] = Fqs007;
assign vis_r2_o[7] = Vss007;
assign vis_r2_o[6] = Lvs007;
assign vis_r2_o[5] = Bys007;
assign vis_r2_o[4] = R0t007;
assign vis_r2_o[3] = H3t007;
assign vis_r2_o[2] = X5t007;
assign vis_r2_o[1] = N8t007;
assign vis_r4_o[0] = Dbt007;
assign vis_r4_o[30] = Tdt007;
assign vis_r4_o[29] = Kgt007;
assign vis_r4_o[28] = Bjt007;
assign vis_r4_o[27] = Slt007;
assign vis_r4_o[26] = Jot007;
assign vis_r4_o[25] = Art007;
assign vis_r4_o[24] = Rtt007;
assign vis_r4_o[23] = Iwt007;
assign vis_r4_o[22] = Zyt007;
assign vis_r4_o[21] = Q1u007;
assign vis_r4_o[20] = H4u007;
assign vis_r4_o[19] = Y6u007;
assign vis_r4_o[18] = P9u007;
assign vis_r4_o[17] = Gcu007;
assign vis_r4_o[16] = Xeu007;
assign vis_r4_o[15] = Ohu007;
assign vis_r4_o[14] = Fku007;
assign vis_r4_o[13] = Wmu007;
assign vis_r4_o[12] = Npu007;
assign vis_r4_o[11] = Esu007;
assign vis_r4_o[10] = Vuu007;
assign vis_r4_o[9] = Mxu007;
assign vis_r4_o[8] = C0v007;
assign vis_r4_o[7] = S2v007;
assign vis_r4_o[6] = I5v007;
assign vis_r4_o[5] = Y7v007;
assign vis_r4_o[4] = Oav007;
assign vis_r4_o[3] = Edv007;
assign vis_r4_o[2] = Ufv007;
assign vis_r4_o[1] = Kiv007;
assign vis_r6_o[0] = Alv007;
assign vis_r6_o[30] = Qnv007;
assign vis_r6_o[29] = Hqv007;
assign vis_r6_o[28] = Ysv007;
assign vis_r6_o[27] = Pvv007;
assign vis_r6_o[26] = Gyv007;
assign vis_r6_o[25] = X0w007;
assign vis_r6_o[24] = O3w007;
assign vis_r6_o[23] = F6w007;
assign vis_r6_o[22] = W8w007;
assign vis_r6_o[21] = Nbw007;
assign vis_r6_o[20] = Eew007;
assign vis_r6_o[19] = Vgw007;
assign vis_r6_o[18] = Mjw007;
assign vis_r6_o[17] = Dmw007;
assign vis_r6_o[16] = Uow007;
assign vis_r6_o[15] = Lrw007;
assign vis_r6_o[14] = Cuw007;
assign vis_r6_o[13] = Tww007;
assign vis_r6_o[12] = Kzw007;
assign vis_r6_o[11] = B2x007;
assign vis_r6_o[10] = S4x007;
assign vis_r6_o[9] = J7x007;
assign vis_r6_o[8] = Z9x007;
assign vis_r6_o[7] = Pcx007;
assign vis_r6_o[6] = Ffx007;
assign vis_r6_o[5] = Vhx007;
assign vis_r6_o[4] = Lkx007;
assign vis_r6_o[3] = Bnx007;
assign vis_r6_o[2] = Rpx007;
assign vis_r6_o[1] = Hsx007;
assign vis_r0_o[0] = Xux007;
assign vis_r0_o[30] = Nxx007;
assign vis_r0_o[29] = E0y007;
assign vis_r0_o[28] = V2y007;
assign vis_r0_o[27] = M5y007;
assign vis_r0_o[26] = D8y007;
assign vis_r0_o[25] = Uay007;
assign vis_r0_o[24] = Ldy007;
assign vis_r0_o[23] = Cgy007;
assign vis_r0_o[22] = Tiy007;
assign vis_r0_o[21] = Kly007;
assign vis_r0_o[20] = Boy007;
assign vis_r0_o[19] = Sqy007;
assign vis_r0_o[18] = Jty007;
assign vis_r0_o[17] = Awy007;
assign vis_r0_o[16] = Ryy007;
assign vis_r0_o[15] = I1z007;
assign vis_r0_o[14] = Z3z007;
assign vis_r0_o[13] = Q6z007;
assign vis_r0_o[12] = H9z007;
assign vis_r0_o[11] = Ybz007;
assign vis_r0_o[10] = Pez007;
assign vis_r0_o[9] = Ghz007;
assign vis_r0_o[8] = Wjz007;
assign vis_r0_o[7] = Mmz007;
assign vis_r0_o[6] = Cpz007;
assign vis_r0_o[5] = Srz007;
assign vis_r0_o[4] = Iuz007;
assign vis_r0_o[3] = Ywz007;
assign vis_r0_o[2] = Ozz007;
assign vis_r0_o[1] = E20107;
assign Byc7z6[30] = U40107;
assign Itb7z6[15] = Y70107;
assign Coxmz6[15] = Qa0107;
assign Krxmz6[15] = Lc0107;
assign Tim7z6[15] = De0107;
assign Hbh7v6 = (!Sg0107);
assign Obh7v6 = (!Wj0107);
assign Tim7z6[23] = An0107;
assign Itb7z6[23] = Pp0107;
assign Coxmz6[23] = Hs0107;
assign Krxmz6[23] = Cu0107;
assign G177z6 = (!Uv0107);
assign Q077z6 = (!Yy0107);
assign Tim7z6[22] = C21107;
assign Itb7z6[22] = R41107;
assign Coxmz6[22] = J71107;
assign Krxmz6[22] = E91107;
assign A077z6 = (!Wa1107);
assign Kz67z6 = (!Ae1107);
assign Tim7z6[21] = Eh1107;
assign Itb7z6[21] = Tj1107;
assign Coxmz6[21] = Lm1107;
assign Krxmz6[21] = Go1107;
assign Uy67z6 = (!Yp1107);
assign Ey67z6 = (!Ct1107);
assign Zec7z6[5] = Gw1107;
assign I9e7z6[1] = Ez1107;
assign I9e7z6[2] = L12107;
assign Byc7z6[5] = S32107;
assign Zec7z6[21] = V62107;
assign Byc7z6[21] = U92107;
assign Tim7z6[20] = Yc2107;
assign Itb7z6[20] = Nf2107;
assign Coxmz6[20] = Fi2107;
assign Krxmz6[20] = Ak2107;
assign Ox67z6 = (!Sl2107);
assign Yw67z6 = (!Wo2107);
assign Zec7z6[4] = As2107;
assign Vjc7z6[1] = Yu2107;
assign Vjc7z6[2] = Xx2107;
assign Vjc7z6[3] = W03107;
assign Vjc7z6[4] = V33107;
assign Vjc7z6[5] = U63107;
assign Vjc7z6[6] = T93107;
assign Vjc7z6[31] = Sc3107;
assign Usbdt6 = Rf3107;
assign M0edt6 = Sh3107;
assign Ic77z6 = (!Sj3107);
assign I9e7z6[0] = Yl3107;
assign Sb77z6 = (!Fo3107);
assign Byc7z6[4] = Oq3107;
assign Zec7z6[20] = Rt3107;
assign V1c7z6[24] = Qw3107;
assign V1c7z6[16] = Wy3107;
assign V1c7z6[9] = C14107;
assign V1c7z6[25] = H34107;
assign V1c7z6[17] = N54107;
assign V1c7z6[10] = T74107;
assign V1c7z6[26] = Z94107;
assign V1c7z6[18] = Fc4107;
assign V1c7z6[11] = Le4107;
assign V1c7z6[19] = Rg4107;
assign V1c7z6[21] = Xi4107;
assign V1c7z6[13] = Dl4107;
assign V1c7z6[22] = Jn4107;
assign V1c7z6[14] = Pp4107;
assign V1c7z6[23] = Vr4107;
assign Ecc7z6[13] = Bu4107;
assign P4c7z6[2] = Ax4107;
assign E8h7z6[2] = Xz4107;
assign Pbadt6 = U25107;
assign Xnh7z6[2] = L55107;
assign Ozbdt6 = I85107;
assign E1uet6 = Ka5107;
assign Ecc7z6[3] = Yc5107;
assign Ecc7z6[6] = Wf5107;
assign Bh2et6 = Ui5107;
assign Ihs7z6[2] = Kl5107;
assign Ihs7z6[3] = En5107;
assign Cch7v6 = (!Yo5107);
assign Ihs7z6[0] = Oq5107;
assign Tn27v6 = Is5107;
assign Zfs7z6[8] = Yt5107;
assign C397z6 = (!Ov5107);
assign Zas7z6[0] = Bx5107;
assign Zfs7z6[11] = Ry5107;
assign Zfs7z6[10] = I06107;
assign Zfs7z6[9] = Z16107;
assign Zfs7z6[7] = P36107;
assign Mm27v6 = F56107;
assign Ap27v6 = V66107;
assign Hq27v6 = L86107;
assign Zas7z6[1] = Ba6107;
assign Z4p7z6[1] = Rb6107;
assign Z4p7z6[2] = Gd6107;
assign Z4p7z6[3] = Ve6107;
assign Z4p7z6[4] = Kg6107;
assign Z4p7z6[5] = Yh6107;
assign W2adt6 = Lj6107;
assign Ow2et6 = Fl6107;
assign Wkb7z6[2] = Zn6107;
assign Gd77z6 = (!Br6107);
assign Ecc7z6[9] = Du6107;
assign Whxdt6 = Bx6107;
assign Ecc7z6[10] = Vz6107;
assign Ecc7z6[11] = U27107;
assign U6i7z6[1] = T57107;
assign U6i7z6[0] = V87107;
assign Ecc7z6[14] = Xb7107;
assign Ibe7z6[4] = We7107;
assign Ibe7z6[1] = Dh7107;
assign Ibe7z6[0] = Kj7107;
assign M3e7z6[1] = Rl7107;
assign V1c7z6[12] = Yn7107;
assign V1c7z6[20] = Eq7107;
assign I2edt6 = Ks7107;
assign M5e7z6[0] = Lu7107;
assign Q1h7z6[0] = Qw7107;
assign Q1h7z6[1] = Qz7107;
assign Q1h7z6[2] = Q28107;
assign Q1h7z6[3] = Q58107;
assign Q1h7z6[4] = Q88107;
assign Q1h7z6[5] = Gttf07;
assign Ecc7z6[5] = Gwtf07;
assign Q9xdt6 = Eztf07;
assign P58et6 = G2uf07;
assign Lvg7z6[0] = G5uf07;
assign Lvg7z6[1] = J8uf07;
assign Lvg7z6[2] = Mbuf07;
assign Z8c7z6[0] = Peuf07;
assign Ntg7z6[0] = Ahuf07;
assign O5h7z6[0] = Xjuf07;
assign Z8c7z6[3] = Umuf07;
assign Ntg7z6[3] = Fpuf07;
assign O5h7z6[3] = Csuf07;
assign Z8c7z6[1] = Zuuf07;
assign Ntg7z6[1] = Kxuf07;
assign O5h7z6[1] = H0vf07;
assign Pxg7z6[3] = E3vf07;
assign M3e7z6[0] = B6vf07;
assign Byc7z6[20] = I8vf07;
assign Tim7z6[19] = Mbvf07;
assign Itb7z6[19] = Bevf07;
assign Coxmz6[19] = Tgvf07;
assign Krxmz6[19] = Oivf07;
assign Iw67z6 = (!Gkvf07);
assign Sv67z6 = (!Knvf07);
assign Tim7z6[18] = Oqvf07;
assign Itb7z6[18] = Dtvf07;
assign Coxmz6[18] = Vvvf07;
assign Krxmz6[18] = Qxvf07;
assign Cv67z6 = (!Izvf07);
assign Mu67z6 = (!M2wf07);
assign Tim7z6[16] = Q5wf07;
assign Itb7z6[16] = F8wf07;
assign Coxmz6[16] = Xawf07;
assign Krxmz6[16] = Scwf07;
assign Byc7z6[16] = Kewf07;
assign W977z6 = (!Ohwf07);
assign Neh7v6 = (!Skwf07);
assign K9h7v6 = (!Wnwf07);
assign Xjh7v6 = (!Lqwf07);
assign Tfh7z6[1] = Ltwf07;
assign Tfh7z6[0] = Jwwf07;
assign Ez2et6 = Hzwf07;
assign R3h7z6[0] = D2xf07;
assign Zdxdt6 = D5xf07;
assign S7xdt6 = A8xf07;
assign R3h7z6[1] = Uaxf07;
assign Gg7et6 = Udxf07;
assign I0c7z6[1] = Ngxf07;
assign Mrbdt6 = Wixf07;
assign Vt2et6 = Xkxf07;
assign Lwfdt6 = Unxf07;
assign V1c7z6[27] = Bqxf07;
assign V1c7z6[28] = Hsxf07;
assign V1c7z6[29] = Nuxf07;
assign V1c7z6[30] = Twxf07;
assign V1c7z6[31] = Zyxf07;
assign V1c7z6[1] = F1yf07;
assign V1c7z6[7] = K3yf07;
assign V1c7z6[6] = P5yf07;
assign Byc7z6[6] = U7yf07;
assign J5n7z6[0] = Xayf07;
assign X9yet6 = Ndyf07;
assign Icyet6 = Dgyf07;
assign T2zet6 = Tiyf07;
assign S0zet6 = Jlyf07;
assign Ryyet6 = Znyf07;
assign Hjn7z6[5] = Pqyf07;
assign Teyet6 = Ftyf07;
assign L9d7z6[4] = Tvyf07;
assign L9d7z6[0] = Xyyf07;
assign Ieadt6 = B2zf07;
assign L9d7z6[2] = E5zf07;
assign Tlb7z6[0] = I8zf07;
assign Wkb7z6[0] = Nazf07;
assign Jqj7z6[2] = Sczf07;
assign Qg77z6 = Tfzf07;
assign Ig77z6 = Thzf07;
assign I6oet6 = Vjzf07;
assign Ja1ft6 = Lmzf07;
assign Orget6 = Fozf07;
assign Euget6 = Zqzf07;
assign C1o7z6[0] = Ptzf07;
assign D02ft6 = Owzf07;
assign Pjb7z6[12] = Byzf07;
assign L877v6 = Yzzf07;
assign Xfymz6[11] = M10g07;
assign Xfymz6[10] = C30g07;
assign Xfymz6[9] = S40g07;
assign Xfymz6[8] = H60g07;
assign Xfymz6[7] = W70g07;
assign Xfymz6[6] = L90g07;
assign Xfymz6[5] = Ab0g07;
assign Xfymz6[4] = Pc0g07;
assign Xfymz6[3] = Ee0g07;
assign Ti2nz6[4] = Tf0g07;
assign Ti2nz6[3] = Zg0g07;
assign Ti2nz6[2] = Fi0g07;
assign Ti2nz6[1] = Lj0g07;
assign J02nz6[3] = Rk0g07;
assign J02nz6[4] = Om0g07;
assign J02nz6[5] = Lo0g07;
assign J02nz6[6] = Iq0g07;
assign J02nz6[7] = Fs0g07;
assign J02nz6[8] = Cu0g07;
assign J02nz6[9] = Zv0g07;
assign J02nz6[10] = Wx0g07;
assign J02nz6[11] = Uz0g07;
assign Coxmz6[12] = S11g07;
assign Krxmz6[12] = N31g07;
assign Tfxmz6[0] = F51g07;
assign Myxmz6[0] = G71g07;
assign Myxmz6[1] = V81g07;
assign Myxmz6[2] = Ka1g07;
assign Myxmz6[3] = Zb1g07;
assign Myxmz6[4] = Od1g07;
assign Uj57v6 = Df1g07;
assign Ikxmz6[1] = Pg1g07;
assign Ikxmz6[2] = Qi1g07;
assign Ovxmz6[1] = Rk1g07;
assign Tim7z6[1] = Mm1g07;
assign Ot67z6 = (!Ap1g07);
assign Ys67z6 = (!Ds1g07);
assign SWDO = Gv1g07;
assign Uz47v6 = Uw1g07;
assign CDBGPWRUPREQ = Iy1g07;
assign Omxmz6[29] = Xz1g07;
assign Qwget6 = L12g07;
assign P1het6 = C42g07;
assign V5k7z6[6] = T62g07;
assign V5k7z6[7] = M92g07;
assign V5k7z6[8] = Fc2g07;
assign V5k7z6[9] = Ye2g07;
assign V5k7z6[10] = Rh2g07;
assign V5k7z6[11] = Lk2g07;
assign V5k7z6[12] = Fn2g07;
assign V5k7z6[13] = Zp2g07;
assign V5k7z6[14] = Ts2g07;
assign V5k7z6[15] = Nv2g07;
assign V5k7z6[16] = Hy2g07;
assign Ui77z6 = (!B13g07);
assign V5k7z6[18] = V33g07;
assign V5k7z6[19] = P63g07;
assign Cj77z6 = (!J93g07);
assign V5k7z6[21] = Dc3g07;
assign V5k7z6[22] = Xe3g07;
assign Kj77z6 = (!Rh3g07);
assign V5k7z6[24] = Lk3g07;
assign V5k7z6[25] = Fn3g07;
assign U297z6 = (!Zp3g07);
assign V5k7z6[27] = Ts3g07;
assign V5k7z6[28] = Nv3g07;
assign V5k7z6[29] = Hy3g07;
assign V5k7z6[30] = B14g07;
assign V5k7z6[5] = V34g07;
assign Gw2ft6 = O64g07;
assign D2fet6 = S84g07;
assign Mah7v6 = (!Ra4g07);
assign Ibe7z6[3] = Tc4g07;
assign Dte7z6[3] = Af4g07;
assign Dte7z6[16] = Yh4g07;
assign Dte7z6[4] = Xk4g07;
assign Dte7z6[5] = Vn4g07;
assign Dte7z6[6] = Tq4g07;
assign Dte7z6[9] = Rt4g07;
assign Dte7z6[10] = Pw4g07;
assign Dte7z6[11] = Oz4g07;
assign Dte7z6[12] = N25g07;
assign Dte7z6[18] = M55g07;
assign Dte7z6[20] = L85g07;
assign Dte7z6[2] = Kb5g07;
assign Dte7z6[0] = Ie5g07;
assign Ehgdt6 = Gh5g07;
assign Djgdt6 = Bk5g07;
assign Dte7z6[19] = Ym5g07;
assign Dte7z6[17] = Xp5g07;
assign Dte7z6[15] = Ws5g07;
assign Dte7z6[14] = Vv5g07;
assign Dte7z6[13] = Uy5g07;
assign Oac7z6[3] = T16g07;
assign Oac7z6[1] = W46g07;
assign Ubhdt6 = Z76g07;
assign Oac7z6[0] = Xa6g07;
assign Dte7z6[7] = Ae6g07;
assign Dte7z6[1] = Yg6g07;
assign Xwe7z6[0] = Wj6g07;
assign Xwe7z6[3] = Xm6g07;
assign Xwe7z6[1] = Yp6g07;
assign Ibe7z6[2] = Zs6g07;
assign Byc7z6[17] = Gv6g07;
assign Rjzet6 = Ky6g07;
assign Ay0ft6 = T07g07;
assign Kb77z6 = (!H37g07);
assign Zjb7z6[8] = P57g07;
assign Tlb7z6[3] = R87g07;
assign Tlb7z6[4] = Tb7g07;
assign Tlb7z6[1] = Ve7g07;
assign Bqi7z6[0] = Xh7g07;
assign Bqi7z6[1] = Ak7g07;
assign Bqi7z6[2] = Dm7g07;
assign Bqi7z6[3] = Go7g07;
assign Toi7z6[5] = Jq7g07;
assign Toi7z6[8] = Ss7g07;
assign Toi7z6[10] = Bv7g07;
assign Toi7z6[11] = Lx7g07;
assign Lxbet6 = Vz7g07;
assign Awbet6 = V18g07;
assign Toi7z6[9] = E48g07;
assign Toi7z6[7] = N68g07;
assign Toi7z6[6] = W88g07;
assign H1j7z6[23] = Fb8g07;
assign H1j7z6[22] = Kd8g07;
assign H1j7z6[21] = Pf8g07;
assign H1j7z6[20] = Uh8g07;
assign H1j7z6[19] = Zj8g07;
assign H1j7z6[18] = Em8g07;
assign H1j7z6[17] = Jo8g07;
assign H1j7z6[15] = Oq8g07;
assign H1j7z6[14] = Ts8g07;
assign H1j7z6[13] = Yu8g07;
assign H1j7z6[12] = Dx8g07;
assign H1j7z6[11] = Iz8g07;
assign H1j7z6[10] = N19g07;
assign H1j7z6[9] = S39g07;
assign H1j7z6[0] = W59g07;
assign H1j7z6[7] = A89g07;
assign H1j7z6[6] = Ea9g07;
assign H1j7z6[5] = Ic9g07;
assign H1j7z6[4] = Me9g07;
assign H1j7z6[3] = Qg9g07;
assign H1j7z6[1] = Ui9g07;
assign Toi7z6[4] = Yk9g07;
assign Toi7z6[3] = Hn9g07;
assign T7j7z6[0] = Qp9g07;
assign T7j7z6[2] = Sr9g07;
assign T7j7z6[1] = Ut9g07;
assign Z8j7z6[0] = Wv9g07;
assign Z8j7z6[2] = Zx9g07;
assign Z8j7z6[1] = C0ag07;
assign Nbj7z6[0] = F2ag07;
assign Nbj7z6[2] = H4ag07;
assign Nbj7z6[1] = J6ag07;
assign Lgj7z6[96] = L8ag07;
assign Lgj7z6[97] = Paag07;
assign Lgj7z6[98] = Tcag07;
assign Lgj7z6[99] = Xeag07;
assign Lgj7z6[100] = Bhag07;
assign Lgj7z6[101] = Gjag07;
assign Lgj7z6[102] = Llag07;
assign Lgj7z6[103] = Qnag07;
assign Lgj7z6[105] = Vpag07;
assign Lgj7z6[106] = Asag07;
assign Lgj7z6[107] = Fuag07;
assign Lgj7z6[0] = Kwag07;
assign Lgj7z6[1] = Nyag07;
assign Lgj7z6[2] = Q0bg07;
assign Lgj7z6[3] = T2bg07;
assign Lgj7z6[4] = W4bg07;
assign Lgj7z6[5] = Z6bg07;
assign Lgj7z6[6] = C9bg07;
assign Lgj7z6[7] = Fbbg07;
assign Lgj7z6[9] = Idbg07;
assign Lgj7z6[10] = Lfbg07;
assign Lgj7z6[11] = Phbg07;
assign Lgj7z6[108] = Tjbg07;
assign Lgj7z6[109] = Ylbg07;
assign Lgj7z6[110] = Dobg07;
assign Lgj7z6[111] = Iqbg07;
assign Lgj7z6[112] = Nsbg07;
assign Lgj7z6[113] = Subg07;
assign Lgj7z6[114] = Xwbg07;
assign Lgj7z6[115] = Czbg07;
assign Lgj7z6[117] = H1cg07;
assign Lgj7z6[118] = M3cg07;
assign Lgj7z6[119] = R5cg07;
assign Lgj7z6[12] = W7cg07;
assign Lgj7z6[13] = Aacg07;
assign Lgj7z6[14] = Eccg07;
assign Lgj7z6[15] = Iecg07;
assign Lgj7z6[16] = Mgcg07;
assign Lgj7z6[17] = Qicg07;
assign Lgj7z6[18] = Ukcg07;
assign Lgj7z6[19] = Ymcg07;
assign Lgj7z6[21] = Cpcg07;
assign Lgj7z6[22] = Grcg07;
assign Lgj7z6[23] = Ktcg07;
assign Micet6 = Ovcg07;
assign Sjcet6 = Nxcg07;
assign Ohj7z6[32] = Mzcg07;
assign Ohj7z6[33] = P1dg07;
assign Ohj7z6[35] = S3dg07;
assign Ohj7z6[36] = V5dg07;
assign Ohj7z6[37] = Y7dg07;
assign Ohj7z6[38] = Badg07;
assign Ohj7z6[39] = Ecdg07;
assign Ohj7z6[41] = Hedg07;
assign Ohj7z6[42] = Kgdg07;
assign Ohj7z6[43] = Nidg07;
assign Ohj7z6[44] = Qkdg07;
assign Ohj7z6[45] = Tmdg07;
assign Ohj7z6[46] = Wodg07;
assign Ohj7z6[47] = Zqdg07;
assign Ohj7z6[56] = Ctdg07;
assign Ohj7z6[57] = Fvdg07;
assign Ohj7z6[58] = Ixdg07;
assign Ohj7z6[59] = Lzdg07;
assign Ohj7z6[60] = O1eg07;
assign Ohj7z6[61] = R3eg07;
assign Ohj7z6[62] = U5eg07;
assign Ohj7z6[63] = X7eg07;
assign Ohj7z6[49] = Aaeg07;
assign Ohj7z6[50] = Dceg07;
assign Ohj7z6[51] = Geeg07;
assign Ohj7z6[52] = Jgeg07;
assign Ohj7z6[53] = Mieg07;
assign Ohj7z6[54] = Pkeg07;
assign Hdcet6 = Smeg07;
assign Jqj7z6[7] = Qpeg07;
assign D5cet6 = Rseg07;
assign L2cet6 = Vueg07;
assign Lgj7z6[155] = Xweg07;
assign Lgj7z6[154] = Czeg07;
assign Lgj7z6[153] = H1fg07;
assign Lgj7z6[151] = M3fg07;
assign Lgj7z6[150] = R5fg07;
assign Lgj7z6[149] = W7fg07;
assign Lgj7z6[148] = Bafg07;
assign Lgj7z6[147] = Gcfg07;
assign Lgj7z6[146] = Lefg07;
assign Lgj7z6[145] = Qgfg07;
assign Lgj7z6[144] = Vifg07;
assign Lgj7z6[59] = Alfg07;
assign Lgj7z6[58] = Enfg07;
assign Lgj7z6[57] = Ipfg07;
assign Lgj7z6[55] = Mrfg07;
assign Lgj7z6[54] = Qtfg07;
assign Lgj7z6[53] = Uvfg07;
assign Lgj7z6[52] = Yxfg07;
assign Lgj7z6[51] = C0gg07;
assign Lgj7z6[50] = G2gg07;
assign Lgj7z6[49] = K4gg07;
assign Lgj7z6[48] = O6gg07;
assign A8cet6 = S8gg07;
assign E9cet6 = Pagg07;
assign Bxi7z6[1] = Qcgg07;
assign Mleet6 = Oegg07;
assign Ijeet6 = Tggg07;
assign Dheet6 = Bjgg07;
assign X6eet6 = Klgg07;
assign Kdadt6 = Ongg07;
assign Qij7z6[6] = Cqgg07;
assign Qij7z6[5] = Jsgg07;
assign Qij7z6[4] = Qugg07;
assign Qij7z6[3] = Xwgg07;
assign P4c7z6[3] = Ezgg07;
assign E8h7z6[3] = B2hg07;
assign Qij7z6[1] = Y4hg07;
assign Qij7z6[0] = F7hg07;
assign Gaj7z6[0] = M9hg07;
assign Gaj7z6[2] = Pbhg07;
assign Gaj7z6[1] = Sdhg07;
assign Bwi7z6[0] = Vfhg07;
assign Bwi7z6[1] = Rhhg07;
assign Bwi7z6[3] = Njhg07;
assign Bwi7z6[4] = Jlhg07;
assign Bwi7z6[5] = Fnhg07;
assign Bwi7z6[6] = Bphg07;
assign Bwi7z6[7] = Xqhg07;
assign Bwi7z6[9] = Tshg07;
assign Bwi7z6[10] = Puhg07;
assign Bwi7z6[11] = Mwhg07;
assign Bwi7z6[12] = Jyhg07;
assign Bwi7z6[13] = G0ig07;
assign Bwi7z6[14] = D2ig07;
assign Bwi7z6[15] = A4ig07;
assign Bwi7z6[17] = X5ig07;
assign Bwi7z6[18] = U7ig07;
assign Bwi7z6[19] = R9ig07;
assign Bwi7z6[20] = Obig07;
assign Bwi7z6[21] = Ldig07;
assign Bwi7z6[22] = Ifig07;
assign Bwi7z6[24] = Fhig07;
assign Bwi7z6[25] = Cjig07;
assign Bwi7z6[26] = Zkig07;
assign Bwi7z6[27] = Wmig07;
assign Bwi7z6[28] = Toig07;
assign Bwi7z6[29] = Qqig07;
assign Bwi7z6[30] = Nsig07;
assign Bwi7z6[31] = Kuig07;
assign Lgj7z6[180] = Hwig07;
assign Lgj7z6[181] = Myig07;
assign Lgj7z6[182] = R0jg07;
assign Lgj7z6[183] = W2jg07;
assign Lgj7z6[184] = B5jg07;
assign Lgj7z6[185] = G7jg07;
assign Lgj7z6[186] = L9jg07;
assign Lgj7z6[187] = Qbjg07;
assign Lgj7z6[189] = Vdjg07;
assign Lgj7z6[190] = Agjg07;
assign Lgj7z6[191] = Fijg07;
assign Lgj7z6[84] = Kkjg07;
assign Lgj7z6[85] = Omjg07;
assign Lgj7z6[86] = Sojg07;
assign Lgj7z6[87] = Wqjg07;
assign Lgj7z6[88] = Atjg07;
assign Lgj7z6[89] = Evjg07;
assign Lgj7z6[90] = Ixjg07;
assign Lgj7z6[91] = Mzjg07;
assign Lgj7z6[93] = Q1kg07;
assign Lgj7z6[94] = U3kg07;
assign Lgj7z6[95] = Y5kg07;
assign Byi7z6[1] = C8kg07;
assign Lgj7z6[132] = Cakg07;
assign Lgj7z6[133] = Hckg07;
assign Lgj7z6[134] = Mekg07;
assign Lgj7z6[135] = Rgkg07;
assign Lgj7z6[136] = Wikg07;
assign Lgj7z6[137] = Blkg07;
assign Lgj7z6[138] = Gnkg07;
assign Lgj7z6[139] = Lpkg07;
assign Lgj7z6[141] = Qrkg07;
assign Lgj7z6[142] = Vtkg07;
assign Lgj7z6[143] = Awkg07;
assign Lgj7z6[36] = Fykg07;
assign Lgj7z6[37] = J0lg07;
assign Lgj7z6[38] = N2lg07;
assign Lgj7z6[39] = R4lg07;
assign Lgj7z6[40] = V6lg07;
assign Lgj7z6[41] = Z8lg07;
assign Lgj7z6[42] = Dblg07;
assign Lgj7z6[43] = Hdlg07;
assign Lgj7z6[45] = Lflg07;
assign Lgj7z6[46] = Phlg07;
assign Lgj7z6[47] = Tjlg07;
assign HTMDHBURST[0] = Xllg07;
assign HTMDHREADY = Bolg07;
assign HTMDHRESP[1] = Qplg07;
assign HTMDHRESP[0] = Hrlg07;
assign Nmq7z6[6] = Yslg07;
assign Nmq7z6[4] = Zulg07;
assign Af4ft6 = Axlg07;
assign Ah4ft6 = Ezlg07;
assign M297z6 = (!I1mg07);
assign Nmq7z6[5] = H3mg07;
assign Nmq7z6[3] = I5mg07;
assign Aj4ft6 = J7mg07;
assign Bbp7z6[0] = F9mg07;
assign Bbp7z6[1] = Lbmg07;
assign Ncp7z6[0] = Rdmg07;
assign Ncp7z6[1] = Xfmg07;
assign L42ft6 = Dimg07;
assign HTMDHPROT[0] = Hkmg07;
assign Nlh7v6 = (!Hkmg07);
assign HTMDHADDR[0] = Ylmg07;
assign Pfh7v6 = (!Ylmg07);
assign HTMDHWRITE = Pnmg07;
assign Cjh7v6 = (!Pnmg07);
assign HTMDHPROT[1] = Epmg07;
assign HTMDHSIZE[1] = Vqmg07;
assign Wfh7v6 = (!Vqmg07);
assign HTMDHSIZE[0] = Msmg07;
assign Kgh7v6 = (!Msmg07);
assign HTMDHADDR[31] = Dumg07;
assign HTMDHADDR[30] = Vvmg07;
assign HTMDHADDR[29] = Nxmg07;
assign HTMDHADDR[28] = Fzmg07;
assign HTMDHADDR[27] = X0ng07;
assign HTMDHADDR[26] = P2ng07;
assign HTMDHADDR[25] = H4ng07;
assign HTMDHADDR[24] = Z5ng07;
assign HTMDHADDR[23] = R7ng07;
assign HTMDHADDR[22] = J9ng07;
assign HTMDHADDR[21] = Bbng07;
assign HTMDHADDR[20] = Tcng07;
assign HTMDHADDR[19] = Leng07;
assign HTMDHADDR[18] = Dgng07;
assign HTMDHADDR[17] = Vhng07;
assign HTMDHADDR[16] = Njng07;
assign HTMDHADDR[15] = Flng07;
assign HTMDHADDR[14] = Xmng07;
assign HTMDHADDR[13] = Pong07;
assign HTMDHADDR[12] = Hqng07;
assign HTMDHADDR[11] = Zrng07;
assign HTMDHADDR[10] = Rtng07;
assign HTMDHADDR[9] = Jvng07;
assign HTMDHADDR[8] = Axng07;
assign HTMDHADDR[7] = Ryng07;
assign HTMDHADDR[6] = I0og07;
assign HTMDHADDR[5] = Z1og07;
assign HTMDHADDR[4] = Q3og07;
assign HTMDHADDR[3] = H5og07;
assign HTMDHADDR[2] = Y6og07;
assign HTMDHADDR[1] = P8og07;
assign Rgh7v6 = (!P8og07);
assign Ea2ft6 = Gaog07;
assign Jexmz6[0] = Ncog07;
assign Jexmz6[1] = Eeog07;
assign Jexmz6[2] = Vfog07;
assign Jexmz6[3] = Mhog07;
assign Jexmz6[4] = Djog07;
assign Jexmz6[5] = Ukog07;
assign Jexmz6[6] = Lmog07;
assign Jexmz6[7] = Coog07;
assign Jexmz6[8] = Tpog07;
assign Jexmz6[9] = Krog07;
assign Jexmz6[10] = Btog07;
assign Jexmz6[11] = Tuog07;
assign Jexmz6[12] = Lwog07;
assign Jexmz6[13] = Dyog07;
assign Jexmz6[14] = Vzog07;
assign Jexmz6[15] = N1pg07;
assign Jexmz6[16] = F3pg07;
assign Jexmz6[17] = X4pg07;
assign Jexmz6[18] = P6pg07;
assign Jexmz6[19] = H8pg07;
assign Jexmz6[20] = Z9pg07;
assign Jexmz6[21] = Rbpg07;
assign Jexmz6[22] = Jdpg07;
assign Jexmz6[23] = Bfpg07;
assign Jexmz6[24] = Tgpg07;
assign Jexmz6[25] = Lipg07;
assign Jexmz6[26] = Dkpg07;
assign Jexmz6[27] = Vlpg07;
assign Jexmz6[29] = Nnpg07;
assign Jexmz6[30] = Fppg07;
assign Jexmz6[31] = Xqpg07;
assign X0eet6 = Pspg07;
assign W2eet6 = Supg07;
assign Yydet6 = Xwpg07;
assign Brdet6 = Azpg07;
assign Zsdet6 = C1qg07;
assign Zudet6 = G3qg07;
assign Ywdet6 = J5qg07;
assign Zodet6 = N7qg07;
assign Nybet6 = T9qg07;
assign Vzbet6 = Ubqg07;
assign Qti7z6[7] = Wdqg07;
assign Pnb7z6[15] = Yfqg07;
assign Qti7z6[9] = Biqg07;
assign Pnb7z6[10] = Dkqg07;
assign Pnb7z6[11] = Gmqg07;
assign Pnb7z6[12] = Joqg07;
assign Pnb7z6[13] = Mqqg07;
assign Pnb7z6[14] = Psqg07;
assign Pnb7z6[17] = Suqg07;
assign Pnb7z6[20] = Vwqg07;
assign Pnb7z6[21] = Yyqg07;
assign Pnb7z6[31] = B1rg07;
assign Pnb7z6[25] = E3rg07;
assign Pnb7z6[26] = H5rg07;
assign Pnb7z6[27] = K7rg07;
assign Pnb7z6[28] = N9rg07;
assign Pnb7z6[29] = Qbrg07;
assign Pnb7z6[30] = Tdrg07;
assign Tcj7z6[0] = Wfrg07;
assign Tcj7z6[2] = Yhrg07;
assign Tcj7z6[1] = Akrg07;
assign Ffj7z6[0] = Cmrg07;
assign Ffj7z6[2] = Eorg07;
assign Ffj7z6[1] = Gqrg07;
assign Zdj7z6[0] = Isrg07;
assign Zdj7z6[2] = Kurg07;
assign Zdj7z6[1] = Mwrg07;
assign Lgj7z6[168] = Oyrg07;
assign Lgj7z6[169] = T0sg07;
assign Lgj7z6[170] = Y2sg07;
assign Lgj7z6[171] = D5sg07;
assign Lgj7z6[172] = I7sg07;
assign Lgj7z6[173] = N9sg07;
assign Lgj7z6[174] = Sbsg07;
assign Lgj7z6[175] = Xdsg07;
assign Lgj7z6[177] = Cgsg07;
assign Lgj7z6[178] = Hisg07;
assign Lgj7z6[179] = Mksg07;
assign Lgj7z6[72] = Rmsg07;
assign Lgj7z6[73] = Vosg07;
assign Lgj7z6[74] = Zqsg07;
assign Lgj7z6[75] = Dtsg07;
assign Lgj7z6[76] = Hvsg07;
assign Lgj7z6[77] = Lxsg07;
assign Lgj7z6[78] = Pzsg07;
assign Lgj7z6[79] = T1tg07;
assign Lgj7z6[81] = X3tg07;
assign Lgj7z6[82] = B6tg07;
assign Lgj7z6[83] = F8tg07;
assign Doadt6 = Jatg07;
assign O7adt6 = Kctg07;
assign Bzi7z6[7] = Letg07;
assign Bzi7z6[9] = Kgtg07;
assign Bzi7z6[10] = Jitg07;
assign Bzi7z6[11] = Iktg07;
assign Bzi7z6[12] = Hmtg07;
assign Bzi7z6[15] = Hotg07;
assign Bzi7z6[17] = Hqtg07;
assign Bzi7z6[18] = Hstg07;
assign Bzi7z6[19] = Hutg07;
assign Bzi7z6[25] = Hwtg07;
assign Bzi7z6[3] = Hytg07;
assign Bzi7z6[4] = G0ug07;
assign Bzi7z6[0] = F2ug07;
assign Lgj7z6[120] = E4ug07;
assign Lgj7z6[121] = J6ug07;
assign Lgj7z6[122] = O8ug07;
assign Lgj7z6[123] = Taug07;
assign Lgj7z6[124] = Ycug07;
assign Lgj7z6[125] = Dfug07;
assign Lgj7z6[126] = Ihug07;
assign Lgj7z6[127] = Njug07;
assign Lgj7z6[129] = Slug07;
assign Lgj7z6[130] = Xnug07;
assign Lgj7z6[131] = Cqug07;
assign Lgj7z6[35] = Hsug07;
assign Lgj7z6[34] = Luug07;
assign Lgj7z6[33] = Pwug07;
assign Lgj7z6[31] = Tyug07;
assign Lgj7z6[30] = X0vg07;
assign Lgj7z6[29] = B3vg07;
assign Lgj7z6[28] = F5vg07;
assign Lgj7z6[27] = J7vg07;
assign Lgj7z6[26] = N9vg07;
assign Lgj7z6[25] = Rbvg07;
assign Lgj7z6[24] = Vdvg07;
assign Dri7z6[17] = Zfvg07;
assign Dri7z6[18] = Aivg07;
assign Dri7z6[19] = Bkvg07;
assign Dri7z6[20] = Cmvg07;
assign Dri7z6[21] = Dovg07;
assign Dri7z6[22] = Eqvg07;
assign Dri7z6[24] = Fsvg07;
assign Dri7z6[25] = Guvg07;
assign Dri7z6[26] = Hwvg07;
assign Dri7z6[27] = Iyvg07;
assign Dri7z6[28] = J0wg07;
assign Dri7z6[29] = K2wg07;
assign Dri7z6[30] = L4wg07;
assign Dri7z6[31] = M6wg07;
assign Dri7z6[9] = N8wg07;
assign Dri7z6[10] = Nawg07;
assign Dri7z6[11] = Ocwg07;
assign Dri7z6[12] = Pewg07;
assign Dri7z6[13] = Qgwg07;
assign Dri7z6[14] = Riwg07;
assign Dri7z6[15] = Skwg07;
assign Dri7z6[7] = Tmwg07;
assign Dri7z6[6] = Towg07;
assign Dri7z6[5] = Tqwg07;
assign Dri7z6[4] = Tswg07;
assign Dri7z6[3] = Tuwg07;
assign Dri7z6[1] = Twwg07;
assign Dri7z6[0] = Tywg07;
assign Dtadt6 = T0xg07;
assign Ku7et6 = U2xg07;
assign R9h7v6 = (!S5xg07);
assign Lgj7z6[156] = Q8xg07;
assign Lgj7z6[157] = Vaxg07;
assign Lgj7z6[158] = Adxg07;
assign Lgj7z6[159] = Ffxg07;
assign Lgj7z6[160] = Khxg07;
assign Lgj7z6[161] = Pjxg07;
assign Lgj7z6[162] = Ulxg07;
assign Lgj7z6[163] = Znxg07;
assign Lgj7z6[165] = Eqxg07;
assign Lgj7z6[166] = Jsxg07;
assign Lgj7z6[167] = Ouxg07;
assign Lgj7z6[71] = Twxg07;
assign Lgj7z6[70] = Xyxg07;
assign Lgj7z6[69] = B1yg07;
assign Lgj7z6[67] = F3yg07;
assign Lgj7z6[66] = J5yg07;
assign Lgj7z6[65] = N7yg07;
assign Lgj7z6[64] = R9yg07;
assign Lgj7z6[63] = Vbyg07;
assign Lgj7z6[62] = Zdyg07;
assign Lgj7z6[61] = Dgyg07;
assign Lgj7z6[60] = Hiyg07;
assign Ohj7z6[0] = Lkyg07;
assign Ohj7z6[1] = Nmyg07;
assign Ohj7z6[3] = Poyg07;
assign Ohj7z6[4] = Rqyg07;
assign Ohj7z6[5] = Tsyg07;
assign Ohj7z6[6] = Vuyg07;
assign Ohj7z6[7] = Xwyg07;
assign Ohj7z6[9] = Zyyg07;
assign Ohj7z6[10] = B1zg07;
assign Ohj7z6[11] = E3zg07;
assign Ohj7z6[12] = H5zg07;
assign Ohj7z6[13] = K7zg07;
assign Ohj7z6[14] = N9zg07;
assign Ohj7z6[15] = Qbzg07;
assign Ohj7z6[17] = Tdzg07;
assign Ohj7z6[18] = Wfzg07;
assign Ohj7z6[19] = Zhzg07;
assign Ohj7z6[20] = Ckzg07;
assign Ohj7z6[21] = Fmzg07;
assign Ohj7z6[22] = Iozg07;
assign Ohj7z6[24] = Lqzg07;
assign Ohj7z6[25] = Oszg07;
assign Ohj7z6[26] = Ruzg07;
assign Ohj7z6[27] = Uwzg07;
assign Ohj7z6[28] = Xyzg07;
assign Ohj7z6[29] = A10h07;
assign Ohj7z6[30] = D30h07;
assign Ohj7z6[31] = G50h07;
assign Wui7z6[30] = J70h07;
assign Wui7z6[28] = L90h07;
assign Wui7z6[31] = Nb0h07;
assign Wui7z6[20] = Pd0h07;
assign Wui7z6[19] = Rf0h07;
assign Wui7z6[18] = Th0h07;
assign Wui7z6[17] = Vj0h07;
assign Wui7z6[14] = Xl0h07;
assign Wui7z6[12] = Zn0h07;
assign Wui7z6[11] = Bq0h07;
assign Wui7z6[10] = Ds0h07;
assign Wui7z6[15] = Fu0h07;
assign Wui7z6[0] = Hw0h07;
assign Wui7z6[6] = Iy0h07;
assign Wui7z6[5] = J01h07;
assign Wui7z6[4] = K21h07;
assign Wui7z6[3] = L41h07;
assign Wui7z6[1] = M61h07;
assign Wui7z6[7] = N81h07;
assign Dtj7z6[2] = Oa1h07;
assign Dtj7z6[5] = Hd1h07;
assign Rmget6 = Ag1h07;
assign Pvj7z6[0] = Ni1h07;
assign Pvj7z6[3] = Ml1h07;
assign Hkget6 = Lo1h07;
assign Dtj7z6[4] = Zq1h07;
assign Dtj7z6[3] = St1h07;
assign Pvj7z6[2] = Lw1h07;
assign Pvj7z6[1] = Kz1h07;
assign Phget6 = J22h07;
assign Weget6 = F52h07;
assign Z4p7z6[0] = C82h07;
assign Hq1ft6 = R92h07;
assign I1p7z6[1] = Fb2h07;
assign A0p7z6[18] = Xc2h07;
assign A0p7z6[15] = Ne2h07;
assign A0p7z6[10] = Dg2h07;
assign A0p7z6[9] = Th2h07;
assign A0p7z6[8] = Ij2h07;
assign A0p7z6[5] = Xk2h07;
assign A0p7z6[4] = Mm2h07;
assign A0p7z6[1] = Bo2h07;
assign A0p7z6[7] = Qp2h07;
assign A0p7z6[11] = Fr2h07;
assign A0p7z6[12] = Vs2h07;
assign A0p7z6[13] = Lu2h07;
assign A0p7z6[19] = Bw2h07;
assign A0p7z6[23] = Rx2h07;
assign A0p7z6[24] = Hz2h07;
assign A0p7z6[25] = X03h07;
assign A0p7z6[26] = N23h07;
assign I1p7z6[0] = D43h07;
assign Iv1ft6 = V53h07;
assign Tx1ft6 = J73h07;
assign W3p7z6[20] = B93h07;
assign W3p7z6[17] = Ra3h07;
assign W3p7z6[12] = Hc3h07;
assign W3p7z6[11] = Xd3h07;
assign W3p7z6[10] = Mf3h07;
assign W3p7z6[7] = Bh3h07;
assign W3p7z6[6] = Qi3h07;
assign W3p7z6[3] = Fk3h07;
assign W3p7z6[9] = Ul3h07;
assign W3p7z6[13] = Jn3h07;
assign W3p7z6[14] = Zo3h07;
assign W3p7z6[15] = Pq3h07;
assign W3p7z6[21] = Fs3h07;
assign W3p7z6[25] = Vt3h07;
assign W3p7z6[26] = Lv3h07;
assign W3p7z6[27] = Bx3h07;
assign W3p7z6[28] = Ry3h07;
assign Nw1ft6 = H04h07;
assign Zy1ft6 = Z14h07;
assign Tk1ft6 = M34h07;
assign Nqo7z6[18] = A54h07;
assign Nqo7z6[15] = Q64h07;
assign Nqo7z6[10] = G84h07;
assign Nqo7z6[9] = W94h07;
assign Nqo7z6[8] = Lb4h07;
assign Nqo7z6[5] = Ad4h07;
assign Nqo7z6[4] = Pe4h07;
assign Nqo7z6[1] = Eg4h07;
assign Nqo7z6[7] = Th4h07;
assign Nqo7z6[11] = Ij4h07;
assign Nqo7z6[12] = Yk4h07;
assign Nqo7z6[13] = Om4h07;
assign Nqo7z6[19] = Eo4h07;
assign Nqo7z6[23] = Up4h07;
assign Nqo7z6[24] = Kr4h07;
assign Nqo7z6[25] = At4h07;
assign Nqo7z6[26] = Qu4h07;
assign Jj1ft6 = Gw4h07;
assign Fpo7z6[18] = Ux4h07;
assign Fpo7z6[15] = Kz4h07;
assign Fpo7z6[9] = A15h07;
assign Fpo7z6[8] = P25h07;
assign Fpo7z6[5] = E45h07;
assign Fpo7z6[4] = T55h07;
assign Fpo7z6[1] = I75h07;
assign Fpo7z6[7] = X85h07;
assign Fpo7z6[11] = Ma5h07;
assign Fpo7z6[12] = Cc5h07;
assign Fpo7z6[13] = Sd5h07;
assign Fpo7z6[23] = If5h07;
assign Fpo7z6[24] = Yg5h07;
assign Fpo7z6[25] = Oi5h07;
assign Fpo7z6[26] = Ek5h07;
assign Rr1ft6 = Ul5h07;
assign Cu1ft6 = In5h07;
assign T2p7z6[20] = Ap5h07;
assign T2p7z6[17] = Qq5h07;
assign T2p7z6[12] = Gs5h07;
assign T2p7z6[11] = Wt5h07;
assign T2p7z6[10] = Lv5h07;
assign T2p7z6[7] = Ax5h07;
assign T2p7z6[6] = Py5h07;
assign T2p7z6[3] = E06h07;
assign T2p7z6[9] = T16h07;
assign T2p7z6[13] = I36h07;
assign T2p7z6[14] = Y46h07;
assign T2p7z6[15] = O66h07;
assign T2p7z6[21] = E86h07;
assign T2p7z6[25] = U96h07;
assign T2p7z6[26] = Kb6h07;
assign T2p7z6[27] = Ad6h07;
assign T2p7z6[28] = Qe6h07;
assign Ws1ft6 = Gg6h07;
assign Nn1ft6 = Yh6h07;
assign Wvo7z6[1] = Mj6h07;
assign Ouo7z6[18] = El6h07;
assign Ouo7z6[15] = Um6h07;
assign Ouo7z6[10] = Ko6h07;
assign Ouo7z6[9] = Aq6h07;
assign Ouo7z6[8] = Pr6h07;
assign Ouo7z6[5] = Et6h07;
assign Ouo7z6[4] = Tu6h07;
assign Ouo7z6[1] = Iw6h07;
assign Ouo7z6[7] = Xx6h07;
assign Ouo7z6[11] = Mz6h07;
assign Ouo7z6[12] = C17h07;
assign Ouo7z6[13] = S27h07;
assign Ouo7z6[19] = I47h07;
assign Ouo7z6[23] = Y57h07;
assign Ouo7z6[24] = O77h07;
assign Ouo7z6[25] = E97h07;
assign Ouo7z6[26] = Ua7h07;
assign Wvo7z6[0] = Kc7h07;
assign Dm1ft6 = Ce7h07;
assign Vro7z6[18] = Qf7h07;
assign Vro7z6[15] = Gh7h07;
assign Vro7z6[10] = Wi7h07;
assign Vro7z6[9] = Mk7h07;
assign Vro7z6[8] = Bm7h07;
assign Vro7z6[5] = Qn7h07;
assign Vro7z6[4] = Fp7h07;
assign Vro7z6[1] = Uq7h07;
assign Vro7z6[7] = Js7h07;
assign Vro7z6[11] = Yt7h07;
assign Vro7z6[12] = Ov7h07;
assign Vro7z6[13] = Ex7h07;
assign Vro7z6[19] = Uy7h07;
assign Vro7z6[23] = K08h07;
assign Vro7z6[24] = A28h07;
assign Vro7z6[25] = Q38h07;
assign Vro7z6[26] = G58h07;
assign Dto7z6[0] = W68h07;
assign Xo1ft6 = O88h07;
assign Pyo7z6[1] = Ca8h07;
assign Hxo7z6[18] = Ub8h07;
assign Hxo7z6[15] = Kd8h07;
assign Hxo7z6[10] = Af8h07;
assign Hxo7z6[9] = Qg8h07;
assign Hxo7z6[8] = Fi8h07;
assign Hxo7z6[5] = Uj8h07;
assign Hxo7z6[4] = Jl8h07;
assign Hxo7z6[1] = Ym8h07;
assign Hxo7z6[7] = No8h07;
assign Hxo7z6[11] = Cq8h07;
assign Hxo7z6[12] = Sr8h07;
assign Hxo7z6[13] = It8h07;
assign Hxo7z6[19] = Yu8h07;
assign Hxo7z6[23] = Ow8h07;
assign Hxo7z6[24] = Ey8h07;
assign Hxo7z6[25] = Uz8h07;
assign Hxo7z6[26] = K19h07;
assign Pyo7z6[0] = A39h07;
assign Goset6 = S49h07;
assign Juset6 = J69h07;
assign O4tet6 = A89h07;
assign P6tet6 = Q99h07;
assign Q8tet6 = Gb9h07;
assign Tetet6 = Wc9h07;
assign Ugtet6 = Me9h07;
assign Ratet6 = Cg9h07;
assign N2tet6 = Sh9h07;
assign M0tet6 = Ij9h07;
assign Lyset6 = Yk9h07;
assign Fmset6 = Pm9h07;
assign Beset6 = Go9h07;
assign Acset6 = Xp9h07;
assign Z9set6 = Or9h07;
assign Sr97z6 = (!Ft9h07);
assign Y7set6 = Ft9h07;
assign E297z6 = (!Wu9h07);
assign Rip7z6[0] = Xw9h07;
assign Rip7z6[3] = Zy9h07;
assign Rip7z6[1] = B1ah07;
assign Pdq7z6[3] = D3ah07;
assign Pdq7z6[1] = J5ah07;
assign G0q7z6[0] = P7ah07;
assign G0q7z6[3] = R9ah07;
assign G0q7z6[1] = Tbah07;
assign Cjq7z6[3] = Vdah07;
assign W22ft6 = Bgah07;
assign I7p7z6[3] = Hiah07;
assign I7p7z6[1] = Jkah07;
assign I7p7z6[0] = Lmah07;
assign M12ft6 = Noah07;
assign E6p7z6[0] = Oqah07;
assign E6p7z6[31] = Msah07;
assign E6p7z6[30] = Luah07;
assign E6p7z6[29] = Kwah07;
assign E6p7z6[28] = Jyah07;
assign E6p7z6[27] = I0bh07;
assign E6p7z6[26] = H2bh07;
assign E6p7z6[25] = G4bh07;
assign E6p7z6[24] = F6bh07;
assign E6p7z6[23] = E8bh07;
assign E6p7z6[22] = Dabh07;
assign E6p7z6[21] = Ccbh07;
assign E6p7z6[20] = Bebh07;
assign E6p7z6[19] = Agbh07;
assign E6p7z6[18] = Zhbh07;
assign E6p7z6[17] = Yjbh07;
assign E6p7z6[16] = Xlbh07;
assign E6p7z6[15] = Wnbh07;
assign E6p7z6[14] = Vpbh07;
assign E6p7z6[13] = Urbh07;
assign E6p7z6[12] = Ttbh07;
assign E6p7z6[11] = Svbh07;
assign E6p7z6[10] = Rxbh07;
assign E6p7z6[9] = Qzbh07;
assign E6p7z6[8] = O1ch07;
assign E6p7z6[7] = M3ch07;
assign E6p7z6[6] = K5ch07;
assign E6p7z6[5] = I7ch07;
assign E6p7z6[4] = G9ch07;
assign E6p7z6[3] = Ebch07;
assign E6p7z6[1] = Cdch07;
assign Bqp7z6[0] = Afch07;
assign Bqp7z6[31] = Chch07;
assign Bqp7z6[30] = Fjch07;
assign Bqp7z6[29] = Ilch07;
assign Bqp7z6[28] = Lnch07;
assign Bqp7z6[27] = Opch07;
assign Bqp7z6[26] = Rrch07;
assign Bqp7z6[25] = Utch07;
assign Bqp7z6[24] = Xvch07;
assign Bqp7z6[23] = Aych07;
assign Bqp7z6[22] = D0dh07;
assign Bqp7z6[21] = G2dh07;
assign Bqp7z6[20] = J4dh07;
assign Bqp7z6[19] = M6dh07;
assign Bqp7z6[18] = P8dh07;
assign Bqp7z6[17] = Sadh07;
assign Bqp7z6[16] = Vcdh07;
assign Bqp7z6[15] = Yedh07;
assign Bqp7z6[14] = Bhdh07;
assign Bqp7z6[13] = Ejdh07;
assign Bqp7z6[12] = Hldh07;
assign Bqp7z6[11] = Kndh07;
assign Bqp7z6[10] = Npdh07;
assign Bqp7z6[9] = Qrdh07;
assign Bqp7z6[8] = Stdh07;
assign Bqp7z6[7] = Uvdh07;
assign Bqp7z6[6] = Wxdh07;
assign Bqp7z6[5] = Yzdh07;
assign Bqp7z6[4] = A2eh07;
assign Bqp7z6[3] = C4eh07;
assign Bqp7z6[1] = E6eh07;
assign Qb4ft6 = G8eh07;
assign Xkq7z6[22] = Daeh07;
assign Xkq7z6[21] = Bceh07;
assign Xkq7z6[20] = Zdeh07;
assign Xkq7z6[19] = Xfeh07;
assign Xkq7z6[18] = Vheh07;
assign Xkq7z6[17] = Tjeh07;
assign Xkq7z6[16] = Rleh07;
assign Xkq7z6[15] = Pneh07;
assign Xkq7z6[14] = Npeh07;
assign Xkq7z6[13] = Lreh07;
assign Xkq7z6[12] = Jteh07;
assign W5q7z6[1] = Hveh07;
assign W5q7z6[0] = Fxeh07;
assign Id4ft6 = Dzeh07;
assign X9q7z6[3] = A1fh07;
assign X9q7z6[2] = X2fh07;
assign X9q7z6[1] = U4fh07;
assign X9q7z6[0] = R6fh07;
assign Y7q7z6[3] = O8fh07;
assign Y7q7z6[2] = Lafh07;
assign Y7q7z6[0] = Icfh07;
assign Dm2ft6 = Fefh07;
assign Hmp7z6[3] = Kgfh07;
assign Hmp7z6[1] = Qifh07;
assign Hmp7z6[0] = Wkfh07;
assign Q8p7z6[0] = Cnfh07;
assign Q8p7z6[3] = Apfh07;
assign Q8p7z6[1] = Yqfh07;
assign Gop7z6[0] = Wsfh07;
assign Gop7z6[3] = Yufh07;
assign Gop7z6[1] = Axfh07;
assign Ei2ft6 = Czfh07;
assign Sgp7z6[3] = H1gh07;
assign Sgp7z6[1] = N3gh07;
assign Sgp7z6[0] = T5gh07;
assign B2q7z6[0] = Z7gh07;
assign B2q7z6[31] = Bagh07;
assign B2q7z6[30] = Ecgh07;
assign B2q7z6[29] = Hegh07;
assign B2q7z6[28] = Kggh07;
assign B2q7z6[27] = Nigh07;
assign B2q7z6[26] = Qkgh07;
assign B2q7z6[25] = Tmgh07;
assign B2q7z6[24] = Wogh07;
assign B2q7z6[23] = Zqgh07;
assign B2q7z6[22] = Ctgh07;
assign B2q7z6[21] = Fvgh07;
assign B2q7z6[20] = Ixgh07;
assign B2q7z6[19] = Lzgh07;
assign B2q7z6[18] = O1hh07;
assign B2q7z6[17] = R3hh07;
assign B2q7z6[16] = U5hh07;
assign B2q7z6[15] = X7hh07;
assign B2q7z6[14] = Aahh07;
assign B2q7z6[13] = Dchh07;
assign B2q7z6[12] = Gehh07;
assign B2q7z6[11] = Jghh07;
assign B2q7z6[10] = Mihh07;
assign B2q7z6[9] = Pkhh07;
assign B2q7z6[8] = Rmhh07;
assign B2q7z6[7] = Tohh07;
assign B2q7z6[6] = Vqhh07;
assign B2q7z6[5] = Xshh07;
assign B2q7z6[4] = Zuhh07;
assign B2q7z6[3] = Bxhh07;
assign B2q7z6[1] = Dzhh07;
assign Mkp7z6[1] = F1ih07;
assign Mkp7z6[3] = H3ih07;
assign Mkp7z6[4] = J5ih07;
assign Mkp7z6[5] = L7ih07;
assign Mkp7z6[6] = N9ih07;
assign Mkp7z6[7] = Pbih07;
assign Mkp7z6[8] = Rdih07;
assign Mkp7z6[9] = Tfih07;
assign Mkp7z6[10] = Vhih07;
assign Mkp7z6[11] = Yjih07;
assign Mkp7z6[12] = Bmih07;
assign Mkp7z6[13] = Eoih07;
assign Mkp7z6[14] = Hqih07;
assign Mkp7z6[15] = Ksih07;
assign Mkp7z6[16] = Nuih07;
assign Mkp7z6[17] = Qwih07;
assign Mkp7z6[18] = Tyih07;
assign Mkp7z6[19] = W0jh07;
assign Mkp7z6[20] = Z2jh07;
assign Mkp7z6[21] = C5jh07;
assign Mkp7z6[22] = F7jh07;
assign Mkp7z6[23] = I9jh07;
assign Mkp7z6[24] = Lbjh07;
assign Mkp7z6[25] = Odjh07;
assign Mkp7z6[26] = Rfjh07;
assign Mkp7z6[27] = Uhjh07;
assign Mkp7z6[28] = Xjjh07;
assign Mkp7z6[29] = Amjh07;
assign Mkp7z6[30] = Dojh07;
assign Mkp7z6[31] = Gqjh07;
assign Mkp7z6[0] = Jsjh07;
assign Gs2ft6 = Lujh07;
assign Hyp7z6[3] = Qwjh07;
assign Hyp7z6[1] = Wyjh07;
assign Hyp7z6[0] = C1kh07;
assign Gwp7z6[1] = I3kh07;
assign Bup7z6[0] = Q5kh07;
assign Bup7z6[1] = C8kh07;
assign Wrp7z6[0] = Oakh07;
assign Wrp7z6[1] = Adkh07;
assign Cq2ft6 = Mfkh07;
assign Gwp7z6[0] = Uhkh07;
assign Pjb7z6[2] = Ckkh07;
assign Xfymz6[2] = Ylkh07;
assign Unymz6[9] = Nnkh07;
assign Unymz6[4] = Fqkh07;
assign Unymz6[6] = Xskh07;
assign Unymz6[7] = Pvkh07;
assign Unymz6[0] = Hykh07;
assign Unymz6[1] = Z0lh07;
assign Unymz6[2] = R3lh07;
assign Unymz6[3] = J6lh07;
assign Unymz6[8] = B9lh07;
assign Ojymz6[9] = Tblh07;
assign Ojymz6[4] = Kelh07;
assign Ojymz6[6] = Bhlh07;
assign Ojymz6[7] = Sjlh07;
assign Ojymz6[0] = Jmlh07;
assign Ojymz6[1] = Aplh07;
assign Ojymz6[2] = Rrlh07;
assign Ojymz6[3] = Iulh07;
assign Ojymz6[8] = Zwlh07;
assign Kmymz6[1] = Qzlh07;
assign Kmymz6[3] = Z1mh07;
assign Blymz6[1] = I4mh07;
assign Blymz6[2] = Q6mh07;
assign Blymz6[3] = Y8mh07;
assign Kmymz6[0] = Gbmh07;
assign At67v6 = Pdmh07;
assign W197z6 = Yfmh07;
assign Wd77z6 = Rhmh07;
assign Cf77z6 = Wjmh07;
assign Kf77z6 = Bmmh07;
assign Sf77z6 = Gomh07;
assign Ag77z6 = Lqmh07;
assign Gh77z6 = Qsmh07;
assign Biymz6[1] = Vumh07;
assign Biymz6[3] = Dxmh07;
assign Biymz6[4] = Lzmh07;
assign Biymz6[5] = T1nh07;
assign Biymz6[6] = B4nh07;
assign Biymz6[7] = J6nh07;
assign Biymz6[9] = R8nh07;
assign Biymz6[10] = Zanh07;
assign Biymz6[11] = Idnh07;
assign Biymz6[12] = Rfnh07;
assign Biymz6[13] = Ainh07;
assign Biymz6[14] = Jknh07;
assign Biymz6[15] = Smnh07;
assign Biymz6[0] = Bpnh07;
assign Feymz6[0] = Jrnh07;
assign Feymz6[1] = Etnh07;
assign Feymz6[2] = Zunh07;
assign Feymz6[3] = Uwnh07;
assign Bfymz6[1] = Pynh07;
assign Bfymz6[2] = K0oh07;
assign Ue77z6 = F2oh07;
assign Jke7v6 = U3oh07;
assign C477v6 = P5oh07;
assign Qc77v6 = G7oh07;
assign Bj77v6 = B9oh07;
assign H71nz6[0] = Kboh07;
assign H71nz6[1] = Idoh07;
assign H71nz6[2] = Gfoh07;
assign H71nz6[3] = Ehoh07;
assign H71nz6[4] = Cjoh07;
assign H71nz6[5] = Aloh07;
assign H71nz6[6] = Ymoh07;
assign H71nz6[7] = Wooh07;
assign H71nz6[8] = Uqoh07;
assign Kkd7v6 = Ssoh07;
assign A377v6 = Ruoh07;
assign Uw77v6 = Pwoh07;
assign W177v6 = Wyoh07;
assign Vv67v6 = W0ph07;
assign Wy67v6 = U2ph07;
assign Qobet6 = R4ph07;
assign O197z6 = (!T6ph07);
assign ETMINTSTAT[1] = W8ph07;
assign Zkh7v6 = (!W8ph07);
assign ETMINTSTAT[0] = Bbph07;
assign Skh7v6 = (!Bbph07);
assign Tjr7z6[6] = Gdph07;
assign Tjr7z6[1] = Qfph07;
assign Tjr7z6[0] = Aiph07;
assign Sr67z6 = (!Kkph07);
assign ETMINTSTAT[2] = Emph07;
assign Glh7v6 = (!Emph07);
assign Soa7v6 = Joph07;
assign Yhzmz6[4] = Hqph07;
assign Thh7v6 = (!Lsph07);
assign Yc77z6 = (!Vuph07);
assign I9b7v6 = Ixph07;
assign Mbc7v6 = Pzph07;
assign Qvb7v6 = R1qh07;
assign G197z6 = (!Z3qh07);
assign Bba7v6 = F6qh07;
assign Tjr7z6[10] = D8qh07;
assign Zxymz6[8] = Oaqh07;
assign Pazmz6[8] = Scqh07;
assign Qmbet6 = Zeqh07;
assign Ie77v6 = Dhqh07;
assign X477v6 = Ejqh07;
assign Ipymz6[1] = Zkqh07;
assign Spc7v6 = Fnqh07;
assign Y097z6 = (!Woqh07);
assign Edh7v6 = (!Uqqh07);
assign Xz67v6 = Vsqh07;
assign Gnzmz6[0] = Nuqh07;
assign Ync7v6 = Lwqh07;
assign Emc7v6 = Kyqh07;
assign Kkc7v6 = J0rh07;
assign Qic7v6 = I2rh07;
assign Wgc7v6 = H4rh07;
assign Cfc7v6 = G6rh07;
assign Gnzmz6[46] = F8rh07;
assign Gnzmz6[45] = Earh07;
assign Gnzmz6[44] = Dcrh07;
assign Gnzmz6[43] = Cerh07;
assign Gnzmz6[42] = Bgrh07;
assign Gnzmz6[41] = Airh07;
assign Gnzmz6[40] = Zjrh07;
assign Gnzmz6[38] = Ylrh07;
assign Gnzmz6[37] = Xnrh07;
assign Gnzmz6[36] = Wprh07;
assign Gnzmz6[35] = Vrrh07;
assign Gnzmz6[34] = Gxps07;
assign Gnzmz6[33] = Fzps07;
assign Gnzmz6[32] = E1qs07;
assign Gnzmz6[30] = D3qs07;
assign Gnzmz6[29] = C5qs07;
assign Gnzmz6[28] = B7qs07;
assign Gnzmz6[27] = A9qs07;
assign Gnzmz6[26] = Zaqs07;
assign Gnzmz6[25] = Ycqs07;
assign Gnzmz6[24] = Xeqs07;
assign Gnzmz6[22] = Wgqs07;
assign Gnzmz6[21] = Viqs07;
assign Gnzmz6[20] = Ukqs07;
assign Gnzmz6[19] = Tmqs07;
assign Gnzmz6[18] = Soqs07;
assign Gnzmz6[17] = Rqqs07;
assign Gnzmz6[16] = Qsqs07;
assign Gnzmz6[14] = Puqs07;
assign Gnzmz6[13] = Owqs07;
assign Gnzmz6[12] = Nyqs07;
assign Gnzmz6[11] = M0rs07;
assign Gnzmz6[10] = L2rs07;
assign Gnzmz6[9] = K4rs07;
assign Gnzmz6[8] = I6rs07;
assign Gnzmz6[6] = G8rs07;
assign Gnzmz6[5] = Ears07;
assign Gnzmz6[4] = Ccrs07;
assign Gnzmz6[3] = Aers07;
assign Gnzmz6[2] = Yfrs07;
assign Gnzmz6[1] = Whrs07;
assign Sgymz6[9] = Ujrs07;
assign Sgymz6[4] = Dmrs07;
assign Sgymz6[6] = Mors07;
assign Sgymz6[7] = Vqrs07;
assign Sgymz6[0] = Etrs07;
assign Sgymz6[1] = Nvrs07;
assign Sgymz6[2] = Wxrs07;
assign Sgymz6[3] = F0ss07;
assign Sgymz6[8] = O2ss07;
assign Ok77v6 = X4ss07;
assign Jdymz6[3] = L7ss07;
assign Jdymz6[0] = G9ss07;
assign Jdymz6[1] = Bbss07;
assign J02nz6[2] = Wcss07;
assign Jw1nz6[3] = Tess07;
assign Jw1nz6[1] = Ngss07;
assign Jw1nz6[0] = Hiss07;
assign Hce7v6 = Bkss07;
assign Nl1nz6[0] = Cmss07;
assign Nl1nz6[1] = Aoss07;
assign Pk1nz6[1] = Ypss07;
assign Pk1nz6[3] = Vrss07;
assign Pk1nz6[6] = Stss07;
assign Pk1nz6[7] = Pvss07;
assign Pk1nz6[10] = Mxss07;
assign Pk1nz6[11] = Kzss07;
assign Pk1nz6[12] = I1ts07;
assign Nyd7v6 = G3ts07;
assign N6h7v6 = C5ts07;
assign M7e7v6 = P7ts07;
assign Fhh7v6 = (!P7ts07);
assign Drf7v6 = Cats07;
assign Td2nz6[1] = Fcts07;
assign Td2nz6[2] = Dets07;
assign Td2nz6[3] = Bgts07;
assign Td2nz6[4] = Zhts07;
assign Td2nz6[5] = Xjts07;
assign Td2nz6[6] = Vlts07;
assign Td2nz6[7] = Tnts07;
assign Td2nz6[8] = Rpts07;
assign Td2nz6[9] = Prts07;
assign Td2nz6[10] = Ntts07;
assign Td2nz6[11] = Mvts07;
assign Td2nz6[12] = Lxts07;
assign Pk1nz6[0] = Kzts07;
assign Pk1nz6[9] = H1us07;
assign Lge7v6 = E3us07;
assign Iy1nz6[1] = D5us07;
assign Gie7v6 = F7us07;
assign Iy1nz6[0] = C9us07;
assign Eee7v6 = Ebus07;
assign Hae7v6 = Fdus07;
assign Ja1nz6[0] = Gfus07;
assign Brg7v6 = Thus07;
assign Fg1nz6[0] = Mkus07;
assign Ti2nz6[0] = Fnus07;
assign Or27v6 = Lous07;
assign Q097z6 = (!Bqus07);
assign Ig27v6 = Prus07;
assign Ln6ft6 = Ntus07;
assign Pp1nz6[0] = Mvus07;
assign U81nz6[0] = Kxus07;
assign Uyg7v6 = Xzus07;
assign Af1nz6[0] = Q2vs07;
assign Oo1nz6[6] = J5vs07;
assign Oo1nz6[5] = H7vs07;
assign Oo1nz6[4] = F9vs07;
assign Oo1nz6[3] = Dbvs07;
assign Oo1nz6[2] = Bdvs07;
assign Oo1nz6[1] = Zevs07;
assign Nn1nz6[6] = Xgvs07;
assign Nn1nz6[5] = Vivs07;
assign Nn1nz6[4] = Tkvs07;
assign Nn1nz6[3] = Rmvs07;
assign Nn1nz6[2] = Povs07;
assign Nn1nz6[1] = Nqvs07;
assign Mm1nz6[1] = Lsvs07;
assign Mm1nz6[0] = Juvs07;
assign U81nz6[2] = Hwvs07;
assign Y3h7v6 = Uyvs07;
assign Af1nz6[2] = N1ws07;
assign Mqb7z6[1] = G4ws07;
assign Mqb7z6[2] = X5ws07;
assign Mqb7z6[3] = O7ws07;
assign Mqb7z6[4] = F9ws07;
assign Mqb7z6[5] = Waws07;
assign Mqb7z6[6] = Ncws07;
assign Rj27v6 = Eews07;
assign Ci6ft6 = Wfws07;
assign D86ft6 = Yhws07;
assign Og6ft6 = Qjws07;
assign Zm37v6 = Ilws07;
assign R8s7z6[0] = Lnws07;
assign R8s7z6[1] = Hpws07;
assign Scs7z6[1] = Drws07;
assign Scs7z6[3] = Atws07;
assign Scs7z6[0] = Xuws07;
assign Ies7z6[24] = Uwws07;
assign Ies7z6[31] = Tyws07;
assign Ies7z6[30] = S0xs07;
assign Ies7z6[29] = R2xs07;
assign Ies7z6[28] = Q4xs07;
assign Ies7z6[27] = P6xs07;
assign Ies7z6[26] = O8xs07;
assign Ies7z6[25] = Naxs07;
assign Ies7z6[15] = Mcxs07;
assign Ies7z6[14] = Lexs07;
assign Ies7z6[13] = Kgxs07;
assign Ies7z6[12] = Jixs07;
assign Ies7z6[11] = Ikxs07;
assign Ies7z6[10] = Hmxs07;
assign Ies7z6[9] = Goxs07;
assign Ies7z6[0] = Fqxs07;
assign Ies7z6[7] = Esxs07;
assign Ies7z6[6] = Duxs07;
assign Ies7z6[5] = Cwxs07;
assign Ies7z6[4] = Byxs07;
assign Ies7z6[3] = A0ys07;
assign Ies7z6[1] = Z1ys07;
assign Ex7et6 = Y3ys07;
assign K1i7z6[1] = V6ys07;
assign K1i7z6[2] = Y9ys07;
assign K1i7z6[5] = Bdys07;
assign K1i7z6[11] = Egys07;
assign K1i7z6[13] = Ijys07;
assign K1i7z6[14] = Mmys07;
assign K1i7z6[15] = Qpys07;
assign K1i7z6[19] = Usys07;
assign K1i7z6[23] = Yvys07;
assign K1i7z6[24] = Czys07;
assign E8h7z6[1] = G2zs07;
assign E3c7z6[0] = D5zs07;
assign Fhc7z6[20] = M7zs07;
assign Fhc7z6[23] = W9zs07;
assign Fhc7z6[14] = Gczs07;
assign Fhc7z6[22] = Qezs07;
assign Fhc7z6[13] = Ahzs07;
assign Fhc7z6[21] = Kjzs07;
assign Fhc7z6[12] = Ulzs07;
assign Fhc7z6[19] = Eozs07;
assign Fhc7z6[17] = Oqzs07;
assign Fhc7z6[9] = Yszs07;
assign Fhc7z6[16] = Hvzs07;
assign Fhc7z6[24] = Rxzs07;
assign Fhc7z6[25] = B00t07;
assign Fhc7z6[10] = L20t07;
assign Fhc7z6[18] = V40t07;
assign E3c7z6[2] = F70t07;
assign Fth7z6[2] = O90t07;
assign Fhc7z6[15] = Lc0t07;
assign Pxg7z6[2] = Ve0t07;
assign Z8c7z6[2] = Sh0t07;
assign Oyfdt6 = Dk0t07;
assign X0cdt6 = Gm0t07;
assign Qdcdt6 = Lo0t07;
assign Osd7z6[1] = Kr0t07;
assign Osd7z6[2] = Ju0t07;
assign Oac7z6[2] = Ix0t07;
assign Xwe7z6[2] = L01t07;
assign Ntg7z6[2] = M31t07;
assign O5h7z6[2] = J61t07;
assign V1c7z6[4] = G91t07;
assign V1c7z6[2] = Lb1t07;
assign Byc7z6[2] = Qd1t07;
assign Y7q7z6[1] = Tg1t07;
assign Bqp7z6[2] = Qi1t07;
assign Gop7z6[2] = Sk1t07;
assign Rip7z6[2] = Um1t07;
assign Hmp7z6[2] = Wo1t07;
assign B82ft6 = Cr1t07;
assign Sgp7z6[2] = Jt1t07;
assign E6p7z6[2] = Pv1t07;
assign Q8p7z6[2] = Nx1t07;
assign B2q7z6[2] = Lz1t07;
assign G0q7z6[2] = N12t07;
assign I7p7z6[2] = P32t07;
assign Zdp7z6[0] = R52t07;
assign Iwymz6[0] = Z72t07;
assign Um4ft6 = Ba2t07;
assign Hyp7z6[2] = Ac2t07;
assign Fy4ft6 = Ge2t07;
assign Dw4ft6 = Fg2t07;
assign Zdp7z6[1] = Li2t07;
assign Iwymz6[1] = Tk2t07;
assign Mkp7z6[2] = Vm2t07;
assign Y52ft6 = Xo2t07;
assign Ayeet6 = Er2t07;
assign Qij7z6[2] = It2t07;
assign Nmadt6 = Pv2t07;
assign U3cet6 = Ox2t07;
assign Hcget6 = Qz2t07;
assign Fjb7z6[0] = J23t07;
assign WICENACK = K33t07;
assign Dpadt6 = J43t07;
assign Me77z6 = (!K63t07);
assign Qg67z6 = (!Q83t07);
assign As67z6 = (!Pa3t07);
assign Cndet6 = Pc3t07;
assign H1j7z6[2] = Qe3t07;
assign X66ft6 = Ug3t07;
assign Scs7z6[2] = Ni3t07;
assign Ies7z6[23] = Kk3t07;
assign Ies7z6[22] = Jm3t07;
assign Ies7z6[21] = Io3t07;
assign Ies7z6[20] = Hq3t07;
assign Ies7z6[19] = Gs3t07;
assign Ies7z6[18] = Fu3t07;
assign Ies7z6[17] = Ew3t07;
assign Ies7z6[2] = Dy3t07;
assign Ee77z6 = C04t07;
assign Kmymz6[2] = H24t07;
assign Biymz6[2] = Q44t07;
assign Hyj7z6[1] = Y64t07;
assign Hyj7z6[3] = V94t07;
assign Hyj7z6[0] = Sc4t07;
assign Hyj7z6[2] = Pf4t07;
assign Bwi7z6[2] = Mi4t07;
assign P6l7z6[20] = Ik4t07;
assign P6l7z6[21] = Zn4t07;
assign P6l7z6[22] = Qr4t07;
assign P6l7z6[23] = Hv4t07;
assign P6l7z6[18] = Vy4t07;
assign P6l7z6[17] = N25t07;
assign P6l7z6[16] = F65t07;
assign P6l7z6[15] = X95t07;
assign P6l7z6[19] = Pd5t07;
assign P6l7z6[10] = Hh5t07;
assign P6l7z6[9] = Tk5t07;
assign P6l7z6[8] = Fo5t07;
assign P6l7z6[7] = Rr5t07;
assign P6l7z6[11] = Dv5t07;
assign P6l7z6[12] = Py5t07;
assign P6l7z6[13] = B26t07;
assign I097z6 = (!N56t07);
assign A097z6 = (!Z86t07);
assign Sz87z6 = (!Lc6t07);
assign Kz87z6 = (!Xf6t07);
assign Cz87z6 = (!Jj6t07);
assign Uy87z6 = (!Vm6t07);
assign Bal7z6[24] = Hq6t07;
assign My87z6 = (!Tt6t07);
assign Ey87z6 = (!Fx6t07);
assign Wx87z6 = (!R07t07);
assign Ox87z6 = (!D47t07);
assign Gx87z6 = (!P77t07);
assign Yw87z6 = (!Bb7t07);
assign Qw87z6 = (!Ne7t07);
assign Iw87z6 = (!Zh7t07);
assign Aw87z6 = (!Ll7t07);
assign Sv87z6 = (!Xo7t07);
assign Kv87z6 = (!Js7t07);
assign Cv87z6 = (!Uv7t07);
assign Uu87z6 = (!Gz7t07);
assign Mu87z6 = (!S28t07);
assign Bal7z6[5] = E68t07;
assign Eu87z6 = (!P98t07);
assign Wt87z6 = (!Ad8t07);
assign P6l7z6[0] = Lg8t07;
assign P6l7z6[1] = Tj8t07;
assign P6l7z6[3] = Gn8t07;
assign P6l7z6[4] = Tq8t07;
assign P6l7z6[5] = Gu8t07;
assign Hwk7z6[20] = Tx8t07;
assign Hwk7z6[21] = K19t07;
assign Hwk7z6[22] = B59t07;
assign Hwk7z6[23] = S89t07;
assign Hwk7z6[18] = Gc9t07;
assign Hwk7z6[17] = Yf9t07;
assign Hwk7z6[16] = Qj9t07;
assign Hwk7z6[15] = In9t07;
assign Hwk7z6[19] = Ar9t07;
assign Hwk7z6[10] = Su9t07;
assign Hwk7z6[9] = Ey9t07;
assign Hwk7z6[8] = Q1at07;
assign Hwk7z6[7] = C5at07;
assign Hwk7z6[11] = O8at07;
assign Hwk7z6[12] = Acat07;
assign Hwk7z6[13] = Mfat07;
assign Ot87z6 = (!Yiat07);
assign Gt87z6 = (!Kmat07);
assign Ys87z6 = (!Wpat07);
assign Qs87z6 = (!Itat07);
assign Is87z6 = (!Uwat07);
assign As87z6 = (!G0bt07);
assign Tzk7z6[24] = S3bt07;
assign Sr87z6 = (!E7bt07);
assign Kr87z6 = (!Qabt07);
assign Cr87z6 = (!Cebt07);
assign Uq87z6 = (!Ohbt07);
assign Mq87z6 = (!Albt07);
assign Eq87z6 = (!Mobt07);
assign Wp87z6 = (!Yrbt07);
assign Op87z6 = (!Kvbt07);
assign Gp87z6 = (!Wybt07);
assign Yo87z6 = (!I2ct07);
assign Qo87z6 = (!U5ct07);
assign Io87z6 = (!F9ct07);
assign Ao87z6 = (!Rcct07);
assign Sn87z6 = (!Dgct07);
assign Tzk7z6[5] = Pjct07;
assign Kn87z6 = (!Anct07);
assign Cn87z6 = (!Lqct07);
assign Hwk7z6[0] = Wtct07;
assign Hwk7z6[1] = Exct07;
assign Hwk7z6[3] = R0dt07;
assign Hwk7z6[4] = E4dt07;
assign Hwk7z6[5] = R7dt07;
assign Zlk7z6[20] = Ebdt07;
assign Zlk7z6[21] = Vedt07;
assign Zlk7z6[22] = Midt07;
assign Zlk7z6[23] = Dmdt07;
assign Zlk7z6[18] = Rpdt07;
assign Zlk7z6[17] = Jtdt07;
assign Zlk7z6[16] = Bxdt07;
assign Zlk7z6[15] = T0et07;
assign Zlk7z6[19] = L4et07;
assign Zlk7z6[10] = D8et07;
assign Zlk7z6[9] = Pbet07;
assign Zlk7z6[8] = Bfet07;
assign Zlk7z6[7] = Niet07;
assign Zlk7z6[11] = Zlet07;
assign Zlk7z6[12] = Lpet07;
assign Zlk7z6[13] = Xset07;
assign Um87z6 = (!Jwet07);
assign Mm87z6 = (!Vzet07);
assign Em87z6 = (!H3ft07);
assign Wl87z6 = (!T6ft07);
assign Ol87z6 = (!Faft07);
assign Gl87z6 = (!Rdft07);
assign Lpk7z6[24] = Dhft07;
assign Yk87z6 = (!Pkft07);
assign Qk87z6 = (!Boft07);
assign Ik87z6 = (!Nrft07);
assign Ak87z6 = (!Zuft07);
assign Sj87z6 = (!Lyft07);
assign Kj87z6 = (!X1gt07);
assign Cj87z6 = (!J5gt07);
assign Ui87z6 = (!V8gt07);
assign Mi87z6 = (!Hcgt07);
assign Ei87z6 = (!Tfgt07);
assign Wh87z6 = (!Fjgt07);
assign Oh87z6 = (!Qmgt07);
assign Gh87z6 = (!Cqgt07);
assign Yg87z6 = (!Otgt07);
assign Lpk7z6[5] = Axgt07;
assign Qg87z6 = (!L0ht07);
assign Ig87z6 = (!W3ht07);
assign Zlk7z6[0] = H7ht07;
assign Zlk7z6[1] = Paht07;
assign Zlk7z6[3] = Ceht07;
assign Zlk7z6[4] = Phht07;
assign Zlk7z6[5] = Clht07;
assign Rbk7z6[20] = Poht07;
assign Rbk7z6[21] = Gsht07;
assign Rbk7z6[22] = Xvht07;
assign Rbk7z6[23] = Ozht07;
assign Rbk7z6[18] = C3it07;
assign Rbk7z6[17] = U6it07;
assign Rbk7z6[16] = Mait07;
assign Rbk7z6[15] = Eeit07;
assign Rbk7z6[19] = Whit07;
assign Rbk7z6[10] = Olit07;
assign Rbk7z6[9] = Apit07;
assign Rbk7z6[8] = Msit07;
assign Rbk7z6[7] = Yvit07;
assign Rbk7z6[11] = Kzit07;
assign Rbk7z6[12] = W2jt07;
assign Rbk7z6[13] = I6jt07;
assign Dfk7z6[30] = U9jt07;
assign Dfk7z6[29] = Gdjt07;
assign Dfk7z6[28] = Sgjt07;
assign Dfk7z6[27] = Ekjt07;
assign Dfk7z6[26] = Qnjt07;
assign Dfk7z6[25] = Crjt07;
assign Dfk7z6[24] = Oujt07;
assign Dfk7z6[31] = Ayjt07;
assign Dfk7z6[22] = M1kt07;
assign Dfk7z6[21] = Y4kt07;
assign Dfk7z6[17] = K8kt07;
assign Dfk7z6[18] = Wbkt07;
assign Dfk7z6[19] = Ifkt07;
assign Dfk7z6[20] = Uikt07;
assign Dfk7z6[15] = Gmkt07;
assign Dfk7z6[14] = Spkt07;
assign Dfk7z6[13] = Etkt07;
assign Dfk7z6[9] = Qwkt07;
assign Dfk7z6[10] = B0lt07;
assign Dfk7z6[11] = N3lt07;
assign Dfk7z6[12] = Z6lt07;
assign Dfk7z6[5] = Lalt07;
assign Dfk7z6[6] = Wdlt07;
assign Dfk7z6[7] = Hhlt07;
assign Rbk7z6[0] = Sklt07;
assign Rbk7z6[1] = Aolt07;
assign Rbk7z6[3] = Nrlt07;
assign Rbk7z6[4] = Avlt07;
assign Rbk7z6[5] = Nylt07;
assign Jw1nz6[2] = A2mt07;
assign Wui7z6[2] = U3mt07;
assign Jdymz6[2] = V5mt07;
assign Apget6 = Q7mt07;
assign Ohj7z6[34] = Pamt07;
assign Ohj7z6[2] = Scmt07;
assign Hyj7z6[5] = Uemt07;
assign Frl7z6[20] = Rhmt07;
assign Frl7z6[21] = Ilmt07;
assign Frl7z6[22] = Zomt07;
assign Frl7z6[23] = Qsmt07;
assign Frl7z6[18] = Ewmt07;
assign Frl7z6[17] = Wzmt07;
assign Frl7z6[16] = O3nt07;
assign Frl7z6[15] = G7nt07;
assign Frl7z6[19] = Yant07;
assign Frl7z6[10] = Qent07;
assign Frl7z6[9] = Cint07;
assign Frl7z6[8] = Olnt07;
assign Frl7z6[7] = Apnt07;
assign Frl7z6[11] = Msnt07;
assign Frl7z6[12] = Yvnt07;
assign Frl7z6[13] = Kznt07;
assign Ag87z6 = (!W2ot07);
assign Sf87z6 = (!I6ot07);
assign Kf87z6 = (!U9ot07);
assign Cf87z6 = (!Gdot07);
assign Ue87z6 = (!Sgot07);
assign Me87z6 = (!Ekot07);
assign Rul7z6[24] = Qnot07;
assign Ee87z6 = (!Crot07);
assign Wd87z6 = (!Ouot07);
assign Od87z6 = (!Ayot07);
assign Gd87z6 = (!M1pt07);
assign Yc87z6 = (!Y4pt07);
assign Qc87z6 = (!K8pt07);
assign Ic87z6 = (!Wbpt07);
assign Ac87z6 = (!Ifpt07);
assign Sb87z6 = (!Uipt07);
assign Kb87z6 = (!Gmpt07);
assign Cb87z6 = (!Sppt07);
assign Ua87z6 = (!Dtpt07);
assign Ma87z6 = (!Pwpt07);
assign Ea87z6 = (!B0qt07);
assign Rul7z6[5] = N3qt07;
assign W987z6 = (!Y6qt07);
assign O987z6 = (!Jaqt07);
assign Frl7z6[0] = Udqt07;
assign Frl7z6[1] = Chqt07;
assign Frl7z6[3] = Pkqt07;
assign Frl7z6[4] = Coqt07;
assign Frl7z6[5] = Prqt07;
assign Hyj7z6[4] = Cvqt07;
assign Xgl7z6[20] = Zxqt07;
assign Xgl7z6[21] = Q1rt07;
assign Xgl7z6[22] = H5rt07;
assign Xgl7z6[23] = Y8rt07;
assign Xgl7z6[18] = Mcrt07;
assign Xgl7z6[17] = Egrt07;
assign Xgl7z6[16] = Wjrt07;
assign Xgl7z6[15] = Onrt07;
assign Xgl7z6[19] = Grrt07;
assign Xgl7z6[10] = Yurt07;
assign Xgl7z6[9] = Kyrt07;
assign Xgl7z6[8] = W1st07;
assign Xgl7z6[7] = I5st07;
assign Xgl7z6[11] = U8st07;
assign Xgl7z6[12] = Gcst07;
assign Xgl7z6[13] = Sfst07;
assign Jkl7z6[30] = Ejst07;
assign Jkl7z6[29] = Qmst07;
assign Jkl7z6[28] = Cqst07;
assign Jkl7z6[27] = Otst07;
assign Jkl7z6[26] = Axst07;
assign Jkl7z6[25] = M0tt07;
assign Jkl7z6[24] = Y3tt07;
assign Jkl7z6[31] = K7tt07;
assign Jkl7z6[22] = Watt07;
assign Jkl7z6[21] = Iett07;
assign Jkl7z6[17] = Uhtt07;
assign Jkl7z6[18] = Gltt07;
assign Jkl7z6[19] = Sott07;
assign Jkl7z6[20] = Estt07;
assign Jkl7z6[15] = Qvtt07;
assign Jkl7z6[14] = Cztt07;
assign Jkl7z6[13] = O2ut07;
assign Jkl7z6[9] = A6ut07;
assign Jkl7z6[10] = L9ut07;
assign Jkl7z6[11] = Xcut07;
assign Jkl7z6[12] = Jgut07;
assign Jkl7z6[5] = Vjut07;
assign Jkl7z6[6] = Gnut07;
assign Jkl7z6[7] = Rqut07;
assign Xgl7z6[0] = Cuut07;
assign Xgl7z6[1] = Kxut07;
assign Xgl7z6[3] = X0vt07;
assign Xgl7z6[4] = K4vt07;
assign Xgl7z6[5] = X7vt07;
assign Hyj7z6[6] = Kbvt07;
assign N1m7z6[20] = Hevt07;
assign N1m7z6[21] = Yhvt07;
assign N1m7z6[22] = Plvt07;
assign N1m7z6[23] = Gpvt07;
assign N1m7z6[18] = Usvt07;
assign N1m7z6[17] = Mwvt07;
assign N1m7z6[16] = E0wt07;
assign N1m7z6[15] = W3wt07;
assign N1m7z6[19] = O7wt07;
assign N1m7z6[10] = Gbwt07;
assign N1m7z6[9] = Sewt07;
assign N1m7z6[8] = Eiwt07;
assign N1m7z6[7] = Qlwt07;
assign N1m7z6[11] = Cpwt07;
assign N1m7z6[12] = Oswt07;
assign N1m7z6[13] = Awwt07;
assign G987z6 = (!Mzwt07);
assign Y887z6 = (!Y2xt07);
assign Q887z6 = (!K6xt07);
assign I887z6 = (!W9xt07);
assign A887z6 = (!Idxt07);
assign S787z6 = (!Ugxt07);
assign Z4m7z6[24] = Gkxt07;
assign K787z6 = (!Snxt07);
assign C787z6 = (!Erxt07);
assign U687z6 = (!Quxt07);
assign M687z6 = (!Cyxt07);
assign E687z6 = (!O1yt07);
assign W587z6 = (!A5yt07);
assign O587z6 = (!M8yt07);
assign G587z6 = (!Ybyt07);
assign Y487z6 = (!Kfyt07);
assign Q487z6 = (!Wiyt07);
assign I487z6 = (!Imyt07);
assign A487z6 = (!Tpyt07);
assign S387z6 = (!Ftyt07);
assign K387z6 = (!Rwyt07);
assign Z4m7z6[5] = D0zt07;
assign C387z6 = (!O3zt07);
assign U287z6 = (!Z6zt07);
assign N1m7z6[0] = Kazt07;
assign N1m7z6[1] = Sdzt07;
assign N1m7z6[3] = Fhzt07;
assign N1m7z6[5] = Skzt07;
assign Hyj7z6[7] = Fozt07;
assign Vbm7z6[20] = Crzt07;
assign Vbm7z6[21] = Tuzt07;
assign Vbm7z6[22] = Kyzt07;
assign Vbm7z6[23] = B20u07;
assign Vbm7z6[15] = P50u07;
assign Vbm7z6[16] = H90u07;
assign Vbm7z6[17] = Zc0u07;
assign Vbm7z6[18] = Rg0u07;
assign Vbm7z6[19] = Jk0u07;
assign Vbm7z6[10] = Bo0u07;
assign Vbm7z6[9] = Nr0u07;
assign Vbm7z6[8] = Zu0u07;
assign Vbm7z6[7] = Ly0u07;
assign Vbm7z6[11] = X11u07;
assign Vbm7z6[12] = J51u07;
assign Vbm7z6[13] = V81u07;
assign Vbm7z6[0] = Hc1u07;
assign Vbm7z6[1] = Pf1u07;
assign Vbm7z6[3] = Cj1u07;
assign Vbm7z6[5] = Pm1u07;
assign M287z6 = (!Cq1u07);
assign E287z6 = (!Ot1u07);
assign W187z6 = (!Ax1u07);
assign O187z6 = (!M02u07);
assign G187z6 = (!Y32u07);
assign Y087z6 = (!K72u07);
assign Q087z6 = (!Wa2u07);
assign I087z6 = (!Ie2u07);
assign A087z6 = (!Uh2u07);
assign Sz77z6 = (!Fl2u07);
assign Kz77z6 = (!Ro2u07);
assign Cz77z6 = (!Ds2u07);
assign Hfm7z6[5] = Pv2u07;
assign Uy77z6 = (!Az2u07);
assign My77z6 = (!L23u07);
assign Ey77z6 = (!W53u07);
assign Wx77z6 = (!I93u07);
assign Ox77z6 = (!Uc3u07);
assign Gx77z6 = (!Gg3u07);
assign Yw77z6 = (!Sj3u07);
assign Qw77z6 = (!En3u07);
assign Hfm7z6[25] = Qq3u07;
assign Iw77z6 = (!Cu3u07);
assign Dri7z6[2] = Ox3u07;
assign Rbk7z6[2] = Oz3u07;
assign Zlk7z6[2] = B34u07;
assign Hwk7z6[2] = O64u07;
assign P6l7z6[2] = Ba4u07;
assign Xgl7z6[2] = Od4u07;
assign Frl7z6[2] = Bh4u07;
assign N1m7z6[2] = Ok4u07;
assign Vbm7z6[2] = Bo4u07;
assign Pk1nz6[2] = Or4u07;
assign W3p7z6[2] = Lt4u07;
assign T2p7z6[2] = Av4u07;
assign A0p7z6[0] = Pw4u07;
assign Hxo7z6[0] = Ey4u07;
assign Ouo7z6[0] = Tz4u07;
assign Vro7z6[0] = I15u07;
assign Nqo7z6[0] = X25u07;
assign Fpo7z6[0] = M45u07;
assign Pdq7z6[2] = B65u07;
assign Cjq7z6[2] = H85u07;
assign vis_pc_o[27] = Na5u07;
assign Fhc7z6[27] = Uc5u07;
assign K1i7z6[27] = Ef5u07;
assign vis_pc_o[28] = Ii5u07;
assign Fhc7z6[28] = Pk5u07;
assign Fth7z6[28] = Zm5u07;
assign K1i7z6[28] = Xp5u07;
assign vis_pc_o[29] = Bt5u07;
assign Fhc7z6[29] = Iv5u07;
assign K1i7z6[29] = Sx5u07;
assign vis_pc_o[30] = W06u07;
assign Dvc7z6[2] = D36u07;
assign Dvc7z6[9] = I66u07;
assign Dvc7z6[12] = N96u07;
assign Dvc7z6[13] = Tc6u07;
assign Dvc7z6[14] = Zf6u07;
assign Dvc7z6[15] = Fj6u07;
assign Dvc7z6[17] = Lm6u07;
assign Dvc7z6[21] = Rp6u07;
assign Dvc7z6[25] = Xs6u07;
assign Dvc7z6[26] = Dw6u07;
assign Dvc7z6[27] = Jz6u07;
assign Dvc7z6[28] = P27u07;
assign Dvc7z6[29] = V57u07;
assign K1i7z6[30] = B97u07;
assign Aw77z6 = Fc7u07;
assign Rzr7z6[1] = Fe7u07;
assign Sv77z6 = Qg7u07;
assign Rzr7z6[2] = Qi7u07;
assign Kv77z6 = Bl7u07;
assign Rzr7z6[3] = Bn7u07;
assign Cv77z6 = Mp7u07;
assign Rzr7z6[4] = Mr7u07;
assign Uu77z6 = Xt7u07;
assign Rzr7z6[5] = Xv7u07;
assign Mu77z6 = Iy7u07;
assign Rzr7z6[6] = I08u07;
assign Eu77z6 = T28u07;
assign Rzr7z6[7] = T48u07;
assign Wt77z6 = E78u07;
assign Rzr7z6[8] = E98u07;
assign Ot77z6 = Pb8u07;
assign Rzr7z6[9] = Pd8u07;
assign Gt77z6 = Ag8u07;
assign Rzr7z6[10] = Bi8u07;
assign Ys77z6 = Nk8u07;
assign Rzr7z6[11] = Om8u07;
assign Qs77z6 = Ap8u07;
assign Rzr7z6[12] = Br8u07;
assign Is77z6 = Nt8u07;
assign Rzr7z6[13] = Ov8u07;
assign As77z6 = Ay8u07;
assign Rzr7z6[14] = B09u07;
assign Sr77z6 = N29u07;
assign Rzr7z6[15] = O49u07;
assign Kr77z6 = A79u07;
assign Rzr7z6[16] = B99u07;
assign Cr77z6 = Nb9u07;
assign Rzr7z6[17] = Od9u07;
assign Uq77z6 = Ag9u07;
assign Rzr7z6[18] = Bi9u07;
assign Mq77z6 = Nk9u07;
assign Rzr7z6[19] = Om9u07;
assign Eq77z6 = Ap9u07;
assign Rzr7z6[20] = Br9u07;
assign Wp77z6 = Nt9u07;
assign Rzr7z6[21] = Ov9u07;
assign Op77z6 = Ay9u07;
assign Rzr7z6[22] = B0au07;
assign Gp77z6 = N2au07;
assign Rzr7z6[23] = O4au07;
assign Yo77z6 = A7au07;
assign Rzr7z6[24] = B9au07;
assign Qo77z6 = Nbau07;
assign Rzr7z6[25] = Odau07;
assign Io77z6 = Agau07;
assign Rzr7z6[26] = Biau07;
assign Ao77z6 = Nkau07;
assign Rzr7z6[27] = Omau07;
assign Sn77z6 = Apau07;
assign Rzr7z6[28] = Brau07;
assign Kn77z6 = Ntau07;
assign Rzr7z6[29] = Ovau07;
assign Cn77z6 = Ayau07;
assign Rzr7z6[30] = B0bu07;
assign Um77z6 = N2bu07;
assign Rzr7z6[31] = O4bu07;
assign Slzmz6[31] = A7bu07;
assign Qk67z6 = (!A7bu07);
assign Slzmz6[1] = A9bu07;
assign Rjzmz6[1] = Zabu07;
assign Jezmz6[1] = Ldbu07;
assign Slzmz6[2] = Sfbu07;
assign Rjzmz6[2] = Rhbu07;
assign Jezmz6[2] = Dkbu07;
assign Slzmz6[3] = Kmbu07;
assign Rjzmz6[3] = Jobu07;
assign Jezmz6[3] = Vqbu07;
assign Slzmz6[4] = Ctbu07;
assign Rjzmz6[4] = Bvbu07;
assign Jezmz6[4] = Nxbu07;
assign Slzmz6[5] = Uzbu07;
assign Rjzmz6[5] = T1cu07;
assign Jezmz6[5] = F4cu07;
assign Slzmz6[6] = M6cu07;
assign Rjzmz6[6] = L8cu07;
assign Jezmz6[6] = Xacu07;
assign Slzmz6[7] = Edcu07;
assign Ik67z6 = (!Edcu07);
assign Rjzmz6[7] = Dfcu07;
assign Slzmz6[8] = Phcu07;
assign Kr67z6 = (!Phcu07);
assign Rjzmz6[8] = Ojcu07;
assign Slzmz6[9] = Amcu07;
assign Cr67z6 = (!Amcu07);
assign Rjzmz6[9] = Zncu07;
assign Slzmz6[10] = Lqcu07;
assign Uq67z6 = (!Lqcu07);
assign Rjzmz6[10] = Lscu07;
assign Slzmz6[11] = Yucu07;
assign Mq67z6 = (!Yucu07);
assign Rjzmz6[11] = Ywcu07;
assign Slzmz6[12] = Lzcu07;
assign Eq67z6 = (!Lzcu07);
assign Rjzmz6[12] = L1du07;
assign Slzmz6[13] = Y3du07;
assign Wp67z6 = (!Y3du07);
assign Rjzmz6[13] = Y5du07;
assign Slzmz6[14] = L8du07;
assign Op67z6 = (!L8du07);
assign Rjzmz6[14] = Ladu07;
assign Slzmz6[15] = Ycdu07;
assign Gp67z6 = (!Ycdu07);
assign Rjzmz6[15] = Yedu07;
assign Slzmz6[16] = Lhdu07;
assign Yo67z6 = (!Lhdu07);
assign Rjzmz6[16] = Ljdu07;
assign Slzmz6[17] = Yldu07;
assign Qo67z6 = (!Yldu07);
assign Rjzmz6[17] = Yndu07;
assign Slzmz6[18] = Lqdu07;
assign Io67z6 = (!Lqdu07);
assign Rjzmz6[18] = Lsdu07;
assign Slzmz6[19] = Yudu07;
assign Ao67z6 = (!Yudu07);
assign Rjzmz6[19] = Ywdu07;
assign Slzmz6[20] = Lzdu07;
assign Rjzmz6[20] = L1eu07;
assign Slzmz6[21] = Y3eu07;
assign Sn67z6 = (!Y3eu07);
assign Rjzmz6[21] = Y5eu07;
assign Slzmz6[22] = L8eu07;
assign Kn67z6 = (!L8eu07);
assign Rjzmz6[22] = Laeu07;
assign Slzmz6[23] = Yceu07;
assign Cn67z6 = (!Yceu07);
assign Rjzmz6[23] = Yeeu07;
assign Slzmz6[24] = Lheu07;
assign Um67z6 = (!Lheu07);
assign Rjzmz6[24] = Ljeu07;
assign Slzmz6[25] = Yleu07;
assign Mm67z6 = (!Yleu07);
assign Rjzmz6[25] = Yneu07;
assign Slzmz6[26] = Lqeu07;
assign Em67z6 = (!Lqeu07);
assign Rjzmz6[26] = Lseu07;
assign Slzmz6[27] = Yueu07;
assign Wl67z6 = (!Yueu07);
assign Rjzmz6[27] = Yweu07;
assign Slzmz6[28] = Lzeu07;
assign Ol67z6 = (!Lzeu07);
assign Rjzmz6[28] = L1fu07;
assign Slzmz6[29] = Y3fu07;
assign Gl67z6 = (!Y3fu07);
assign Rjzmz6[29] = Y5fu07;
assign Slzmz6[30] = L8fu07;
assign Yk67z6 = (!L8fu07);
assign Rjzmz6[30] = Lafu07;
assign Rjzmz6[31] = Ycfu07;
assign Hk5ft6 = Lffu07;
assign Mi5ft6 = Mhfu07;
assign Kg5ft6 = Ljfu07;
assign Lfp7z6[3] = Rlfu07;
assign Zdp7z6[3] = Rnfu07;
assign Iwymz6[3] = Zpfu07;
assign A05ft6 = Bsfu07;
assign Po4ft6 = Cufu07;
assign J95ft6 = Dwfu07;
assign O75ft6 = Eyfu07;
assign Lfp7z6[2] = D0gu07;
assign Zdp7z6[2] = D2gu07;
assign Iwymz6[2] = L4gu07;
assign Jqj7z6[3] = N6gu07;
assign Cmbdt6 = O9gu07;
assign LOCKUP = Pbgu07;
assign Mhh7v6 = (!Pbgu07);
assign Ac77z6 = Ndgu07;
assign Qjh7v6 = (!Ofgu07);
assign W1a7v6 = Uhgu07;
assign Pqddt6 = Akgu07;
assign Loddt6 = Imgu07;
assign H1j7z6[8] = Qogu07;
assign H56ft6 = Uqgu07;
assign Ies7z6[8] = Xsgu07;
assign T077v6 = Wugu07;
assign Q4c7v6 = Vwgu07;
assign Ro87v6 = Azgu07;
assign Oob7v6 = D1hu07;
assign Qxb7v6 = E3hu07;
assign P3zmz6[8] = H5hu07;
assign P3zmz6[9] = K7hu07;
assign P3zmz6[10] = N9hu07;
assign P3zmz6[11] = Rbhu07;
assign P3zmz6[12] = Vdhu07;
assign P3zmz6[13] = Zfhu07;
assign P3zmz6[14] = Dihu07;
assign P3zmz6[15] = Hkhu07;
assign P3zmz6[16] = Lmhu07;
assign P3zmz6[17] = Pohu07;
assign P3zmz6[18] = Tqhu07;
assign P3zmz6[19] = Xshu07;
assign P3zmz6[20] = Bvhu07;
assign P3zmz6[21] = Fxhu07;
assign P3zmz6[22] = Jzhu07;
assign P3zmz6[23] = N1iu07;
assign P3zmz6[24] = R3iu07;
assign P3zmz6[25] = V5iu07;
assign P3zmz6[26] = Z7iu07;
assign P3zmz6[27] = Daiu07;
assign P3zmz6[28] = Hciu07;
assign P3zmz6[29] = Leiu07;
assign P3zmz6[30] = Pgiu07;
assign P3zmz6[31] = Tiiu07;
assign Jezmz6[15] = Xkiu07;
assign Jezmz6[23] = Fniu07;
assign Jezmz6[31] = Npiu07;
assign P3zmz6[7] = Vriu07;
assign Jezmz6[10] = Ytiu07;
assign Jezmz6[11] = Gwiu07;
assign Jezmz6[12] = Oyiu07;
assign Jezmz6[13] = W0ju07;
assign Jezmz6[16] = E3ju07;
assign Jezmz6[17] = M5ju07;
assign Jezmz6[18] = U7ju07;
assign Jezmz6[19] = Caju07;
assign Jezmz6[20] = Kcju07;
assign Jezmz6[21] = Seju07;
assign Jezmz6[24] = Ahju07;
assign Jezmz6[25] = Ijju07;
assign Jezmz6[26] = Qlju07;
assign Jezmz6[27] = Ynju07;
assign Jezmz6[28] = Gqju07;
assign Jezmz6[29] = Osju07;
assign Jezmz6[34] = Wuju07;
assign Jezmz6[35] = Exju07;
assign Jezmz6[8] = Mzju07;
assign Jezmz6[9] = T1ku07;
assign Sgymz6[5] = A4ku07;
assign Ojymz6[5] = J6ku07;
assign Biymz6[8] = A9ku07;
assign Ruymz6[8] = Ibku07;
assign Uh77v6 = Gdku07;
assign Ruymz6[15] = Afku07;
assign Ruymz6[0] = Zgku07;
assign Ruymz6[1] = Xiku07;
assign Ruymz6[2] = Vkku07;
assign Ruymz6[3] = Tmku07;
assign Ruymz6[4] = Roku07;
assign Ruymz6[5] = Pqku07;
assign Ruymz6[6] = Nsku07;
assign Ruymz6[7] = Luku07;
assign Ruymz6[9] = Jwku07;
assign Ruymz6[10] = Hyku07;
assign Ruymz6[11] = G0lu07;
assign Ruymz6[12] = F2lu07;
assign Ruymz6[13] = E4lu07;
assign Ruymz6[14] = D6lu07;
assign Unymz6[5] = C8lu07;
assign Bwi7z6[8] = Ualu07;
assign Bzi7z6[8] = Qclu07;
assign Wui7z6[8] = Pelu07;
assign Dri7z6[8] = Qglu07;
assign Ohj7z6[40] = Qilu07;
assign Ohj7z6[8] = Tklu07;
assign Rbk7z6[6] = Vmlu07;
assign Dfk7z6[8] = Hqlu07;
assign Zlk7z6[6] = Stlu07;
assign Lpk7z6[8] = Exlu07;
assign Hwk7z6[6] = P0mu07;
assign Tzk7z6[8] = B4mu07;
assign P6l7z6[6] = M7mu07;
assign Bal7z6[8] = Yamu07;
assign Xgl7z6[6] = Jemu07;
assign Jkl7z6[8] = Vhmu07;
assign Frl7z6[6] = Glmu07;
assign Rul7z6[8] = Somu07;
assign N1m7z6[6] = Dsmu07;
assign Z4m7z6[8] = Pvmu07;
assign Vbm7z6[6] = Azmu07;
assign Hfm7z6[8] = M2nu07;
assign Pk1nz6[8] = X5nu07;
assign Qti7z6[8] = U7nu07;
assign Sctet6 = W9nu07;
assign W3p7z6[8] = Mbnu07;
assign T2p7z6[8] = Bdnu07;
assign A0p7z6[6] = Qenu07;
assign Hxo7z6[6] = Fgnu07;
assign Ouo7z6[6] = Uhnu07;
assign Vro7z6[6] = Jjnu07;
assign Nqo7z6[6] = Yknu07;
assign Fpo7z6[6] = Nmnu07;
assign K1i7z6[8] = Conu07;
assign vis_psp_o[7] = Frnu07;
assign K1i7z6[7] = Wtnu07;
assign Fhc7z6[7] = Ee9917;
assign Dvc7z6[7] = Ng9917;
assign vis_psp_o[6] = Sj9917;
assign K1i7z6[6] = Jm9917;
assign Fhc7z6[6] = Mp9917;
assign Dvc7z6[6] = Vr9917;
assign Ppb7z6[6] = Av9917;
assign vis_psp_o[4] = Ix9917;
assign E3c7z6[4] = Zz9917;
assign vis_psp_o[3] = I2a917;
assign K1i7z6[3] = Z4a917;
assign E3c7z6[3] = C8a917;
assign Qmb7z6[1] = Laa917;
assign Qmb7z6[3] = Hda917;
assign Qmb7z6[5] = Dga917;
assign Qmb7z6[6] = Zia917;
assign Qmb7z6[7] = Vla917;
assign Qmb7z6[0] = Roa917;
assign Ykcet6 = Nra917;
assign E1cet6 = Mta917;
assign H1j7z6[16] = Mva917;
assign A0j7z6[16] = Rxa917;
assign A0j7z6[0] = Vza917;
assign M5bdt6 = Y1b917;
assign Jqj7z6[8] = W3b917;
assign Macet6 = X6b917;
assign A0j7z6[1] = A9b917;
assign A0j7z6[2] = Dbb917;
assign A0j7z6[3] = Gdb917;
assign A0j7z6[4] = Jfb917;
assign A0j7z6[5] = Mhb917;
assign A0j7z6[6] = Pjb917;
assign A0j7z6[7] = Slb917;
assign A0j7z6[8] = Vnb917;
assign A0j7z6[9] = Ypb917;
assign A0j7z6[10] = Bsb917;
assign A0j7z6[11] = Fub917;
assign A0j7z6[12] = Jwb917;
assign A0j7z6[13] = Nyb917;
assign A0j7z6[14] = R0c917;
assign A0j7z6[15] = V2c917;
assign A0j7z6[17] = Z4c917;
assign A0j7z6[18] = D7c917;
assign A0j7z6[19] = H9c917;
assign A0j7z6[20] = Lbc917;
assign A0j7z6[21] = Pdc917;
assign A0j7z6[22] = Tfc917;
assign A0j7z6[23] = Xhc917;
assign Mqb7z6[0] = Bkc917;
assign Ies7z6[16] = Slc917;
assign Bfymz6[0] = Rnc917;
assign Sgymz6[10] = Mpc917;
assign Ojymz6[10] = Vrc917;
assign Blymz6[0] = Muc917;
assign Tn77v6 = Uwc917;
assign Unymz6[10] = Vyc917;
assign Fjd7v6 = N1d917;
assign Hcymz6[1] = C4d917;
assign Hcymz6[2] = R6d917;
assign Hcymz6[3] = G9d917;
assign G7bdt6 = Vbd917;
assign Nob7z6[0] = Ydd917;
assign Tjr7z6[2] = Dgd917;
assign Yhzmz6[0] = Nid917;
assign Nob7z6[7] = Rkd917;
assign Tjr7z6[9] = Wmd917;
assign Zxymz6[7] = Gpd917;
assign Pazmz6[7] = Krd917;
assign Nob7z6[6] = Rtd917;
assign Tjr7z6[8] = Wvd917;
assign Zxymz6[6] = Gyd917;
assign Pazmz6[6] = K0e917;
assign Nob7z6[5] = R2e917;
assign G5j7z6[32] = W4e917;
assign M6j7z6[32] = V7e917;
assign G5j7z6[0] = Uae917;
assign M6j7z6[0] = Sde917;
assign G5j7z6[16] = Qge917;
assign M6j7z6[16] = Pje917;
assign Tjr7z6[7] = Ome917;
assign Zxymz6[5] = Yoe917;
assign Pazmz6[5] = Cre917;
assign Nob7z6[3] = Jte917;
assign Tjr7z6[5] = Ove917;
assign Yhzmz6[3] = Yxe917;
assign Nob7z6[1] = C0f917;
assign G5j7z6[44] = H2f917;
assign M6j7z6[44] = G5f917;
assign G5j7z6[28] = F8f917;
assign M6j7z6[28] = Ebf917;
assign G5j7z6[12] = Def917;
assign M6j7z6[12] = Chf917;
assign Z3j7z6[8] = Bkf917;
assign Bxi7z6[4] = Zmf917;
assign G5j7z6[35] = Wof917;
assign M6j7z6[35] = Vrf917;
assign G5j7z6[19] = Uuf917;
assign M6j7z6[19] = Txf917;
assign G5j7z6[3] = S0g917;
assign M6j7z6[3] = R3g917;
assign G5j7z6[43] = Q6g917;
assign M6j7z6[43] = P9g917;
assign G5j7z6[27] = Ocg917;
assign M6j7z6[27] = Nfg917;
assign G5j7z6[11] = Mig917;
assign M6j7z6[11] = Llg917;
assign G5j7z6[31] = Kog917;
assign M6j7z6[31] = Jrg917;
assign G5j7z6[15] = Iug917;
assign Z3j7z6[11] = Hxg917;
assign Zfcet6 = F0h917;
assign G5j7z6[46] = D3h917;
assign M6j7z6[46] = C6h917;
assign G5j7z6[14] = B9h917;
assign M6j7z6[14] = Ach917;
assign G5j7z6[30] = Zeh917;
assign M6j7z6[30] = Yhh917;
assign G5j7z6[33] = Xkh917;
assign M6j7z6[33] = Wnh917;
assign G5j7z6[17] = Vqh917;
assign M6j7z6[17] = Uth917;
assign G5j7z6[1] = Twh917;
assign M6j7z6[1] = Szh917;
assign G5j7z6[41] = R2i917;
assign M6j7z6[41] = Q5i917;
assign G5j7z6[25] = P8i917;
assign M6j7z6[25] = Obi917;
assign G5j7z6[9] = Nei917;
assign M6j7z6[9] = Mhi917;
assign G5j7z6[61] = Lki917;
assign M6j7z6[61] = Kni917;
assign G5j7z6[13] = Jqi917;
assign M6j7z6[13] = Iti917;
assign G5j7z6[29] = Hwi917;
assign M6j7z6[29] = Gzi917;
assign G5j7z6[45] = F2j917;
assign M6j7z6[45] = E5j917;
assign Tjr7z6[3] = D8j917;
assign Yhzmz6[1] = Naj917;
assign G5j7z6[47] = Rcj917;
assign M6j7z6[47] = Qfj917;
assign G5j7z6[62] = Pij917;
assign M6j7z6[62] = Olj917;
assign X3get6 = Noj917;
assign SYSRESETREQ = Lrj917;
assign Hsi7z6[2] = Qtj917;
assign Hsi7z6[1] = Vvj917;
assign Hsi7z6[0] = Ayj917;
assign Dri7z6[16] = F0k917;
assign Ohj7z6[16] = G2k917;
assign Ohj7z6[48] = J4k917;
assign Bwi7z6[16] = M6k917;
assign Rbk7z6[14] = J8k917;
assign Dfk7z6[16] = Bck917;
assign Zlk7z6[14] = Nfk917;
assign Lpk7z6[16] = Fjk917;
assign Hwk7z6[14] = Rmk917;
assign Tzk7z6[16] = Jqk917;
assign P6l7z6[14] = Vtk917;
assign Bal7z6[16] = Nxk917;
assign Xgl7z6[14] = Z0l917;
assign Jkl7z6[16] = R4l917;
assign Frl7z6[14] = D8l917;
assign Rul7z6[16] = Vbl917;
assign N1m7z6[14] = Hfl917;
assign Z4m7z6[16] = Zil917;
assign Vbm7z6[14] = Lml917;
assign Hfm7z6[16] = Dql917;
assign Pnb7z6[16] = Ptl917;
assign Dvc7z6[16] = Svl917;
assign Kwset6 = Yyl917;
assign W3p7z6[16] = P0m917;
assign T2p7z6[16] = F2m917;
assign A0p7z6[14] = V3m917;
assign Hxo7z6[14] = L5m917;
assign Ouo7z6[14] = B7m917;
assign Vro7z6[14] = R8m917;
assign Nqo7z6[14] = Ham917;
assign Fpo7z6[14] = Xbm917;
assign Bzi7z6[16] = Ndm917;
assign Wui7z6[16] = Nfm917;
assign Iynet6 = Phm917;
assign Bxi7z6[3] = Ikm917;
assign Lgj7z6[8] = Emm917;
assign Lgj7z6[20] = Hom917;
assign Lgj7z6[32] = Lqm917;
assign Lgj7z6[44] = Psm917;
assign Lgj7z6[56] = Tum917;
assign Lgj7z6[68] = Xwm917;
assign Lgj7z6[80] = Bzm917;
assign Lgj7z6[92] = F1n917;
assign Lgj7z6[104] = J3n917;
assign Lgj7z6[116] = O5n917;
assign Lgj7z6[128] = T7n917;
assign Lgj7z6[140] = Y9n917;
assign Lgj7z6[152] = Dcn917;
assign Lgj7z6[164] = Ien917;
assign Lgj7z6[176] = Ngn917;
assign Lgj7z6[188] = Sin917;
assign Ohj7z6[23] = Xkn917;
assign Ohj7z6[55] = Ann917;
assign Dri7z6[23] = Dpn917;
assign Bwi7z6[23] = Ern917;
assign Dfk7z6[23] = Btn917;
assign Mm77z6 = (!Nwn917);
assign Em77z6 = (!Zzn917);
assign Wl77z6 = (!L3o917);
assign Jkl7z6[23] = X6o917;
assign Ol77z6 = (!Jao917);
assign Gl77z6 = (!Vdo917);
assign Yk77z6 = (!Hho917);
assign U9p7z6[23] = Tko917;
assign U9p7z6[0] = Vmo917;
assign U9p7z6[1] = Woo917;
assign U9p7z6[2] = Xqo917;
assign U9p7z6[3] = Yso917;
assign U9p7z6[4] = Zuo917;
assign U9p7z6[5] = Axo917;
assign U9p7z6[6] = Bzo917;
assign U9p7z6[7] = C1p917;
assign U9p7z6[8] = D3p917;
assign U9p7z6[9] = E5p917;
assign U9p7z6[10] = F7p917;
assign Gy2ft6 = H9p917;
assign W3q7z6[0] = Nbp917;
assign W3q7z6[1] = Udp917;
assign W3q7z6[2] = Bgp917;
assign W3q7z6[3] = Iip917;
assign V1s7z6[5] = Pkp917;
assign Cu5ft6 = Dnp917;
assign Gqr7z6[31] = Spp917;
assign Gqr7z6[30] = Bsp917;
assign Gqr7z6[29] = Kup917;
assign Gqr7z6[28] = Twp917;
assign Gqr7z6[27] = Czp917;
assign Gqr7z6[26] = L1q917;
assign Gqr7z6[25] = U3q917;
assign Gqr7z6[24] = D6q917;
assign Gqr7z6[23] = M8q917;
assign Gqr7z6[22] = Vaq917;
assign Gqr7z6[21] = Edq917;
assign Gqr7z6[20] = Nfq917;
assign Gqr7z6[19] = Whq917;
assign Gqr7z6[18] = Fkq917;
assign Gqr7z6[17] = Omq917;
assign Gqr7z6[16] = Xoq917;
assign Gqr7z6[15] = Grq917;
assign Gqr7z6[14] = Ptq917;
assign Gqr7z6[13] = Yvq917;
assign Gqr7z6[12] = Hyq917;
assign Gqr7z6[11] = Q0r917;
assign Gqr7z6[10] = Z2r917;
assign Gqr7z6[9] = I5r917;
assign Gqr7z6[8] = Q7r917;
assign Gqr7z6[7] = Y9r917;
assign Gqr7z6[6] = Gcr917;
assign Gqr7z6[5] = Oer917;
assign Gqr7z6[4] = Wgr917;
assign Gqr7z6[3] = Ejr917;
assign Gqr7z6[2] = Mlr917;
assign Gqr7z6[1] = Unr917;
assign U9p7z6[11] = Cqr917;
assign U9p7z6[12] = Esr917;
assign U9p7z6[13] = Gur917;
assign U9p7z6[14] = Iwr917;
assign U9p7z6[15] = Kyr917;
assign U9p7z6[16] = M0s917;
assign U9p7z6[17] = O2s917;
assign U9p7z6[18] = Q4s917;
assign U9p7z6[19] = S6s917;
assign U9p7z6[20] = U8s917;
assign U9p7z6[21] = Was917;
assign U9p7z6[22] = Ycs917;
assign U9p7z6[25] = Afs917;
assign U9p7z6[26] = Chs917;
assign U9p7z6[27] = Ejs917;
assign U9p7z6[28] = Gls917;
assign Hu2ft6 = Ins917;
assign Txadt6 = Lps917;
assign Ur37v6 = Krs917;
assign I96ft6 = Ats917;
assign X9s7z6[16] = Tus917;
assign X9s7z6[11] = Qws917;
assign X9s7z6[10] = Nys917;
assign X9s7z6[8] = K0t917;
assign X9s7z6[7] = G2t917;
assign X9s7z6[6] = C4t917;
assign X9s7z6[5] = Y5t917;
assign X9s7z6[4] = U7t917;
assign X9s7z6[3] = Q9t917;
assign X9s7z6[1] = Mbt917;
assign X9s7z6[22] = Idt917;
assign X9s7z6[23] = Fft917;
assign X9s7z6[24] = Cht917;
assign X9s7z6[0] = Zit917;
assign G1e7v6 = Vkt917;
assign Cmg7v6 = Tmt917;
assign L9e7v6 = Ipt917;
assign I6e7v6 = Xrt917;
assign Iyf7v6 = Qtt917;
assign Ekh7v6 = (!Bwt917);
assign Xre7v6 = Myt917;
assign Md1nz6[2] = K0u917;
assign X7g7v6 = X2u917;
assign Lj1nz6[2] = N5u917;
assign Md1nz6[1] = D8u917;
assign L5g7v6 = Qau917;
assign Fah7v6 = (!Gdu917);
assign Md1nz6[0] = Wfu917;
assign Z2g7v6 = Jiu917;
assign Lj1nz6[0] = Zku917;
assign F2f7v6 = Pnu917;
assign J7f7v6 = Opu917;
assign B5e7v6 = Mru917;
assign P0g7v6 = Ktu917;
assign Lkh7v6 = (!Yvu917);
assign Xzd7v6 = Myu917;
assign Nog7v6 = N0v917;
assign M8e7v6 = F3v917;
assign T5f7v6 = X5v917;
assign Od77z6 = (!R7v917);
assign Qa2nz6[1] = J9v917;
assign Yb1nz6[2] = Ebv917;
assign Hfg7v6 = Rdv917;
assign Hi1nz6[2] = Hgv917;
assign Yb1nz6[1] = Xiv917;
assign Vcg7v6 = Klv917;
assign Y9h7v6 = (!Aov917);
assign Yb1nz6[0] = Qqv917;
assign Jag7v6 = Dtv917;
assign Hi1nz6[0] = Tvv917;
assign Mwf7v6 = Jyv917;
assign Ctf7v6 = J0w917;
assign Qk77z6 = (!G2w917);
assign Kf2nz6[0] = G4w917;
assign Kf2nz6[1] = D6w917;
assign Kf2nz6[2] = A8w917;
assign D92nz6[0] = X9w917;
assign Ec2nz6[0] = Rbw917;
assign Ec2nz6[1] = Ndw917;
assign Ec2nz6[2] = Jfw917;
assign Ec2nz6[3] = Fhw917;
assign Dxe7v6 = Bjw917;
assign D92nz6[1] = Ykw917;
assign Kve7v6 = Smw917;
assign T32nz6[0] = Pow917;
assign T32nz6[1] = Qqw917;
assign T32nz6[2] = Rsw917;
assign T32nz6[3] = Suw917;
assign Qa2nz6[0] = Tww917;
assign Ah2nz6[0] = Oyw917;
assign Ah2nz6[1] = O0x917;
assign Ah2nz6[2] = O2x917;
assign M2e7v6 = O4x917;
assign Vjg7v6 = T6x917;
assign Hbe7v6 = E9x917;
assign Ak6ft6 = Pbx917;
assign Id6ft6 = Mdx917;
assign Vis7z6[3] = Efx917;
assign Vis7z6[2] = Dhx917;
assign Vis7z6[1] = Cjx917;
assign Vis7z6[0] = Blx917;
assign Vis7z6[4] = Anx917;
assign A4f7v6 = Zox917;
assign R0f7v6 = Wqx917;
assign Ik77z6 = (!Osx917);
assign U9p7z6[29] = Jux917;
assign U9p7z6[30] = Lwx917;
assign U9p7z6[31] = Nyx917;
assign Pnb7z6[23] = P0y917;
assign Dvc7z6[23] = S2y917;
assign Diset6 = Y5y917;
assign W3p7z6[23] = P7y917;
assign T2p7z6[23] = F9y917;
assign A0p7z6[21] = Vay917;
assign Hxo7z6[21] = Lcy917;
assign Ouo7z6[21] = Bey917;
assign Vro7z6[21] = Rfy917;
assign Nqo7z6[21] = Hhy917;
assign Fpo7z6[21] = Xiy917;
assign Wui7z6[23] = Nky917;
assign X9s7z6[31] = Pmy917;
assign Coxmz6[31] = Moy917;
assign Krxmz6[31] = Hqy917;
assign TDO = Zry917;
assign Pmh7v6 = (!Lty917);
assign Sk4ft6 = Ovy917;
assign M55ft6 = Uxy917;
assign Wlr7z6[1] = A0z917;
assign Wlr7z6[2] = N2z917;
assign Wlr7z6[3] = A5z917;
assign Wlr7z6[5] = N7z917;
assign Wlr7z6[6] = Aaz917;
assign Wlr7z6[8] = Ncz917;
assign Wlr7z6[9] = Afz917;
assign Wlr7z6[10] = Nhz917;
assign Wlr7z6[11] = Bkz917;
assign Wlr7z6[13] = Pmz917;
assign Wlr7z6[14] = Dpz917;
assign Wlr7z6[16] = Rrz917;
assign Wlr7z6[17] = Fuz917;
assign Wlr7z6[18] = Twz917;
assign Wlr7z6[19] = Hzz917;
assign Wlr7z6[21] = V10a17;
assign Wlr7z6[22] = J40a17;
assign Wlr7z6[24] = X60a17;
assign Wlr7z6[25] = L90a17;
assign Wlr7z6[26] = Zb0a17;
assign Wlr7z6[27] = Ne0a17;
assign Wlr7z6[29] = Bh0a17;
assign Wlr7z6[30] = Pj0a17;
assign Dfr7z6[0] = Dm0a17;
assign Dfr7z6[1] = Qo0a17;
assign Vr5ft6 = Dr0a17;
assign Xcr7z6[0] = Ot0a17;
assign Xcr7z6[1] = Bw0a17;
assign Wlr7z6[0] = Oy0a17;
assign J5n7z6[1] = B11a17;
assign BRCHSTAT[3] = R31a17;
assign Byc7z6[28] = N61a17;
assign Jexmz6[28] = R91a17;
assign Wlr7z6[28] = Jb1a17;
assign Wlr7z6[20] = Xd1a17;
assign Wlr7z6[12] = Lg1a17;
assign Wlr7z6[4] = Zi1a17;
assign K1i7z6[4] = Ml1a17;
assign G5j7z6[49] = Po1a17;
assign M6j7z6[49] = Or1a17;
assign G5j7z6[51] = Nu1a17;
assign M6j7z6[51] = Mx1a17;
assign G5j7z6[57] = L02a17;
assign M6j7z6[57] = K32a17;
assign G5j7z6[59] = J62a17;
assign M6j7z6[59] = I92a17;
assign G5j7z6[63] = Hc2a17;
assign K1i7z6[16] = Gf2a17;
assign G5j7z6[56] = Ki2a17;
assign M6j7z6[56] = Jl2a17;
assign G5j7z6[40] = Io2a17;
assign M6j7z6[40] = Hr2a17;
assign G5j7z6[24] = Gu2a17;
assign M6j7z6[24] = Fx2a17;
assign G5j7z6[8] = E03a17;
assign M6j7z6[8] = D33a17;
assign G5j7z6[50] = C63a17;
assign M6j7z6[50] = B93a17;
assign G5j7z6[34] = Ac3a17;
assign M6j7z6[34] = Ze3a17;
assign G5j7z6[18] = Yh3a17;
assign M6j7z6[18] = Xk3a17;
assign G5j7z6[2] = Wn3a17;
assign M6j7z6[2] = Vq3a17;
assign G5j7z6[58] = Ut3a17;
assign M6j7z6[58] = Tw3a17;
assign G5j7z6[42] = Sz3a17;
assign M6j7z6[42] = R24a17;
assign G5j7z6[26] = Q54a17;
assign M6j7z6[26] = P84a17;
assign G5j7z6[10] = Ob4a17;
assign M6j7z6[10] = Ne4a17;
assign G5j7z6[52] = Mh4a17;
assign M6j7z6[52] = Lk4a17;
assign G5j7z6[36] = Kn4a17;
assign M6j7z6[36] = Jq4a17;
assign G5j7z6[20] = It4a17;
assign M6j7z6[20] = Hw4a17;
assign G5j7z6[4] = Gz4a17;
assign M6j7z6[4] = F25a17;
assign Z3j7z6[0] = E55a17;
assign G5j7z6[53] = C85a17;
assign M6j7z6[53] = Bb5a17;
assign G5j7z6[37] = Ae5a17;
assign M6j7z6[37] = Zg5a17;
assign G5j7z6[5] = Yj5a17;
assign G5j7z6[21] = Xm5a17;
assign M6j7z6[21] = Wp5a17;
assign G5j7z6[54] = Vs5a17;
assign M6j7z6[54] = Uv5a17;
assign G5j7z6[38] = Ty5a17;
assign M6j7z6[38] = S16a17;
assign G5j7z6[6] = R46a17;
assign M6j7z6[6] = Q76a17;
assign G5j7z6[22] = Pa6a17;
assign M6j7z6[22] = Od6a17;
assign Z3j7z6[3] = Ng6a17;
assign Z3j7z6[12] = Lj6a17;
assign G5j7z6[55] = Jm6a17;
assign G5j7z6[39] = Ip6a17;
assign M6j7z6[39] = Hs6a17;
assign G5j7z6[23] = Gv6a17;
assign M6j7z6[23] = Fy6a17;
assign Moj7z6[0] = E17a17;
assign G5j7z6[7] = I37a17;
assign M6j7z6[7] = H67a17;
assign Tjr7z6[4] = G97a17;
assign Yhzmz6[2] = Qb7a17;
assign Pazmz6[4] = Ud7a17;
assign Hbb7v6 = Bg7a17;
assign Fgzmz6[1] = Ei7a17;
assign L587v6 = Ik7a17;
assign Ka87v6 = Gm7a17;
assign Gnzmz6[39] = Fo7a17;
assign Gnzmz6[31] = Eq7a17;
assign Gnzmz6[23] = Ds7a17;
assign Gnzmz6[15] = Cu7a17;
assign B987v6 = Bw7a17;
assign De87v6 = Zx7a17;
assign Jezmz6[33] = Tz7a17;
assign Ztb7v6 = B28a17;
assign Cdb7v6 = A48a17;
assign Xfd7v6 = O68a17;
assign E11nz6[0] = O88a17;
assign E11nz6[1] = Ma8a17;
assign E11nz6[2] = Kc8a17;
assign E11nz6[3] = Ie8a17;
assign E11nz6[4] = Gg8a17;
assign Uu0nz6[3] = Ei8a17;
assign Uu0nz6[2] = Ck8a17;
assign Uu0nz6[0] = Am8a17;
assign Uu0nz6[1] = Yn8a17;
assign R21nz6[0] = Wp8a17;
assign T51nz6[0] = Nr8a17;
assign R21nz6[1] = Mt8a17;
assign T51nz6[1] = Dv8a17;
assign Jezmz6[32] = Cx8a17;
assign Zt67v6 = Kz8a17;
assign T51nz6[2] = M19a17;
assign Vm0nz6[3] = L39a17;
assign Vm0nz6[6] = I59a17;
assign Lo0nz6[3] = F79a17;
assign Lo0nz6[6] = C99a17;
assign R21nz6[2] = Za9a17;
assign Ttzmz6[0] = Qc9a17;
assign Jvzmz6[0] = Ne9a17;
assign Zwzmz6[0] = Kg9a17;
assign Dd0nz6[0] = Hi9a17;
assign Te0nz6[0] = Ek9a17;
assign Jg0nz6[0] = Bm9a17;
assign L30nz6[0] = Yn9a17;
assign B50nz6[0] = Vp9a17;
assign R60nz6[0] = Sr9a17;
assign Vm0nz6[0] = Pt9a17;
assign Lo0nz6[0] = Mv9a17;
assign Bq0nz6[0] = Jx9a17;
assign Pazmz6[3] = Gz9a17;
assign Pazmz6[0] = N1aa17;
assign Pazmz6[1] = U3aa17;
assign Xozmz6[2] = B6aa17;
assign Nqzmz6[2] = Y7aa17;
assign Dszmz6[2] = V9aa17;
assign H80nz6[2] = Sbaa17;
assign X90nz6[2] = Pdaa17;
assign Nb0nz6[2] = Mfaa17;
assign Ttzmz6[2] = Jhaa17;
assign Jvzmz6[2] = Gjaa17;
assign Zwzmz6[2] = Dlaa17;
assign Dd0nz6[2] = Anaa17;
assign Te0nz6[2] = Xoaa17;
assign Jg0nz6[2] = Uqaa17;
assign Pyzmz6[2] = Rsaa17;
assign F00nz6[2] = Ouaa17;
assign V10nz6[2] = Lwaa17;
assign Zh0nz6[2] = Iyaa17;
assign Pj0nz6[2] = F0ba17;
assign Fl0nz6[2] = C2ba17;
assign L30nz6[2] = Z3ba17;
assign B50nz6[2] = W5ba17;
assign R60nz6[2] = T7ba17;
assign Vm0nz6[2] = Q9ba17;
assign Lo0nz6[2] = Nbba17;
assign Bq0nz6[2] = Kdba17;
assign Pazmz6[2] = Hfba17;
assign K1i7z6[10] = Ohba17;
assign X9s7z6[34] = Skba17;
assign K1i7z6[18] = Pmba17;
assign Yr1nz6[2] = Tpba17;
assign Xq1nz6[2] = Rrba17;
assign Ft0nz6[2] = Ptba17;
assign Ft0nz6[3] = Pvba17;
assign Jezmz6[30] = Pxba17;
assign Jezmz6[22] = Xzba17;
assign Jezmz6[14] = F2ca17;
assign Xozmz6[3] = N4ca17;
assign Nqzmz6[3] = K6ca17;
assign Dszmz6[3] = H8ca17;
assign H80nz6[3] = Eaca17;
assign X90nz6[3] = Bcca17;
assign Nb0nz6[3] = Ydca17;
assign Ttzmz6[3] = Vfca17;
assign Jvzmz6[3] = Shca17;
assign Zwzmz6[3] = Pjca17;
assign Dd0nz6[3] = Mlca17;
assign Te0nz6[3] = Jnca17;
assign Jg0nz6[3] = Gpca17;
assign Pyzmz6[3] = Drca17;
assign F00nz6[3] = Atca17;
assign V10nz6[3] = Xuca17;
assign Zh0nz6[3] = Uwca17;
assign Pj0nz6[3] = Ryca17;
assign Fl0nz6[3] = O0da17;
assign L30nz6[3] = L2da17;
assign B50nz6[3] = I4da17;
assign R60nz6[3] = F6da17;
assign Xozmz6[1] = C8da17;
assign Nqzmz6[1] = Z9da17;
assign Dszmz6[1] = Wbda17;
assign H80nz6[1] = Tdda17;
assign X90nz6[1] = Qfda17;
assign Nb0nz6[1] = Nhda17;
assign Ttzmz6[1] = Kjda17;
assign Jvzmz6[1] = Hlda17;
assign Zwzmz6[1] = Enda17;
assign Dd0nz6[1] = Bpda17;
assign Te0nz6[1] = Yqda17;
assign Jg0nz6[1] = Vsda17;
assign Pyzmz6[1] = Suda17;
assign F00nz6[1] = Pwda17;
assign V10nz6[1] = Myda17;
assign Zh0nz6[1] = J0ea17;
assign Pj0nz6[1] = G2ea17;
assign Fl0nz6[1] = D4ea17;
assign L30nz6[1] = A6ea17;
assign B50nz6[1] = X7ea17;
assign R60nz6[1] = U9ea17;
assign Vm0nz6[1] = Rbea17;
assign Lo0nz6[1] = Odea17;
assign Bq0nz6[1] = Lfea17;
assign Wh67z6 = Ihea17;
assign Bv1nz6[1] = Djea17;
assign Au1nz6[1] = Blea17;
assign Zs1nz6[1] = Zmea17;
assign S677v6 = Xoea17;
assign Qch7v6 = (!Xqea17);
assign Byc7z6[9] = Tsea17;
assign Tim7z6[8] = Wvea17;
assign Svn7z6[0] = Kyea17;
assign Svn7z6[2] = J1fa17;
assign Svn7z6[1] = I4fa17;
assign Vbm7z6[4] = H7fa17;
assign Tbq7z6[4] = Uafa17;
assign Tbq7z6[0] = Bdfa17;
assign Tbq7z6[1] = Iffa17;
assign Tbq7z6[2] = Phfa17;
assign Tbq7z6[3] = Wjfa17;
assign Tbq7z6[5] = Dmfa17;
assign Tbq7z6[6] = Kofa17;
assign Tbq7z6[7] = Rqfa17;
assign V1s7z6[4] = Ysfa17;
assign Kfq7z6[4] = Mvfa17;
assign Kfq7z6[1] = Uxfa17;
assign Kfq7z6[2] = C0ga17;
assign Kfq7z6[3] = K2ga17;
assign Kfq7z6[5] = S4ga17;
assign Kfq7z6[6] = A7ga17;
assign Kfq7z6[7] = I9ga17;
assign Pk1nz6[4] = Qbga17;
assign W3p7z6[4] = Ndga17;
assign T2p7z6[4] = Cfga17;
assign A0p7z6[2] = Rgga17;
assign Hxo7z6[2] = Giga17;
assign Ouo7z6[2] = Vjga17;
assign Vro7z6[2] = Klga17;
assign Nqo7z6[2] = Zmga17;
assign Fpo7z6[2] = Ooga17;
assign Pdq7z6[4] = Dqga17;
assign Cjq7z6[4] = Jsga17;
assign X9s7z6[12] = Puga17;
assign Hcymz6[4] = Mwga17;
assign Mi77z6 = Bzga17;
assign L9cdt6 = V0ha17;
assign D6c7z6[4] = V2ha17;
assign D6c7z6[1] = X5ha17;
assign D7hdt6 = Z8ha17;
assign Mpe7z6[5] = Qbha17;
assign Xpgdt6 = Ieha17;
assign Bsgdt6 = Ahha17;
assign Pne7z6[0] = Sjha17;
assign Mpe7z6[2] = Omha17;
assign Mpe7z6[3] = Gpha17;
assign Mpe7z6[4] = Yrha17;
assign Pne7z6[1] = Quha17;
assign Ple7z6[1] = Mxha17;
assign Ple7z6[2] = L0ia17;
assign Ple7z6[3] = K3ia17;
assign Ple7z6[4] = J6ia17;
assign Ple7z6[5] = I9ia17;
assign Ple7z6[6] = Hcia17;
assign Ple7z6[0] = Gfia17;
assign Ple7z6[7] = Fiia17;
assign Yxf7z6[2] = Elia17;
assign Yxf7z6[6] = Ynia17;
assign Yxf7z6[10] = Sqia17;
assign Yxf7z6[14] = Ntia17;
assign Yxf7z6[18] = Iwia17;
assign Yxf7z6[22] = Dzia17;
assign Yxf7z6[26] = Y1ja17;
assign Yxf7z6[30] = T4ja17;
assign Yxf7z6[34] = O7ja17;
assign Alf7z6[24] = Jaja17;
assign Alf7z6[21] = Hdja17;
assign Cngdt6 = Fgja17;
assign Ppb7z6[5] = Ejja17;
assign Kxb7z6[5] = Mlja17;
assign Alf7z6[0] = Vnja17;
assign Alf7z6[1] = Sqja17;
assign Alf7z6[2] = Ptja17;
assign Alf7z6[3] = Mwja17;
assign Alf7z6[4] = Jzja17;
assign Alf7z6[5] = G2ka17;
assign Alf7z6[6] = D5ka17;
assign Alf7z6[7] = A8ka17;
assign Alf7z6[15] = Xaka17;
assign Alf7z6[16] = Vdka17;
assign Alf7z6[8] = Tgka17;
assign Alf7z6[9] = Qjka17;
assign Alf7z6[10] = Nmka17;
assign Alf7z6[11] = Lpka17;
assign Alf7z6[12] = Jska17;
assign Alf7z6[13] = Hvka17;
assign Alf7z6[14] = Fyka17;
assign Alf7z6[17] = D1la17;
assign Alf7z6[18] = B4la17;
assign Alf7z6[19] = Z6la17;
assign Alf7z6[20] = X9la17;
assign Alf7z6[22] = Vcla17;
assign Alf7z6[23] = Tfla17;
assign Alf7z6[25] = Rila17;
assign Alf7z6[26] = Plla17;
assign Alf7z6[27] = Nola17;
assign Alf7z6[30] = Lrla17;
assign Alf7z6[28] = Jula17;
assign Alf7z6[29] = Hxla17;
assign Yxf7z6[1] = F0ma17;
assign Yxf7z6[5] = Z2ma17;
assign Yxf7z6[9] = T5ma17;
assign Yxf7z6[13] = N8ma17;
assign Yxf7z6[17] = Ibma17;
assign Yxf7z6[21] = Dema17;
assign Yxf7z6[25] = Ygma17;
assign Yxf7z6[29] = Tjma17;
assign Yxf7z6[33] = Omma17;
assign Onf7z6[0] = Jpma17;
assign Onf7z6[1] = Gsma17;
assign Onf7z6[2] = Dvma17;
assign Onf7z6[3] = Ayma17;
assign Onf7z6[4] = X0na17;
assign Onf7z6[5] = U3na17;
assign Onf7z6[6] = R6na17;
assign Onf7z6[7] = O9na17;
assign Onf7z6[8] = Lcna17;
assign Onf7z6[9] = Ifna17;
assign Onf7z6[10] = Fina17;
assign Onf7z6[11] = Dlna17;
assign Onf7z6[12] = Bona17;
assign Onf7z6[13] = Zqna17;
assign Onf7z6[14] = Xtna17;
assign Onf7z6[15] = Vwna17;
assign Onf7z6[16] = Tzna17;
assign Onf7z6[17] = R2oa17;
assign Onf7z6[18] = P5oa17;
assign Onf7z6[19] = N8oa17;
assign Onf7z6[20] = Lboa17;
assign Onf7z6[21] = Jeoa17;
assign Onf7z6[22] = Hhoa17;
assign Onf7z6[23] = Fkoa17;
assign Onf7z6[24] = Dnoa17;
assign Onf7z6[25] = Bqoa17;
assign Onf7z6[26] = Zsoa17;
assign Onf7z6[27] = Xvoa17;
assign Onf7z6[28] = Vyoa17;
assign Onf7z6[29] = T1pa17;
assign Fth7z6[5] = R4pa17;
assign Pdc7z6[5] = O7pa17;
assign Dvc7z6[5] = Oapa17;
assign Iufdt6 = Tdpa17;
assign Uyb7z6[1] = Agpa17;
assign Uyb7z6[4] = Kipa17;
assign Uyb7z6[3] = Ukpa17;
assign Uyb7z6[0] = Enpa17;
assign Z3j7z6[1] = Oppa17;
assign Z3j7z6[14] = Mspa17;
assign Wbcet6 = Kvpa17;
assign Efcdt6 = Pxpa17;
assign Fk2ft6 = M0qa17;
assign HTMDHTRANS[0] = O2qa17;
assign Gg2ft6 = G4qa17;
assign Xy5ft6 = I6qa17;
assign Jhr7z6[0] = S8qa17;
assign Jhr7z6[1] = Jbqa17;
assign Cor7z6[0] = Aeqa17;
assign Cor7z6[1] = Lgqa17;
assign Cor7z6[2] = Wiqa17;
assign Cor7z6[3] = Hlqa17;
assign Cor7z6[4] = Snqa17;
assign Cor7z6[5] = Dqqa17;
assign Cor7z6[6] = Osqa17;
assign Cor7z6[7] = Zuqa17;
assign Cor7z6[8] = Kxqa17;
assign Cor7z6[9] = Vzqa17;
assign Cor7z6[10] = G2ra17;
assign Cor7z6[11] = S4ra17;
assign Cor7z6[12] = E7ra17;
assign Cor7z6[13] = Q9ra17;
assign Cor7z6[14] = Ccra17;
assign Cor7z6[15] = Oera17;
assign Cor7z6[16] = Ahra17;
assign Cor7z6[17] = Mjra17;
assign Cor7z6[18] = Ylra17;
assign Cor7z6[19] = Kora17;
assign Cor7z6[20] = Wqra17;
assign Cor7z6[21] = Itra17;
assign Cor7z6[22] = Uvra17;
assign Cor7z6[23] = Gyra17;
assign Cor7z6[24] = S0sa17;
assign Cor7z6[25] = E3sa17;
assign Cor7z6[26] = Q5sa17;
assign Cor7z6[27] = C8sa17;
assign Cor7z6[28] = Oasa17;
assign Cor7z6[29] = Adsa17;
assign Cor7z6[30] = Mfsa17;
assign Cor7z6[31] = Yhsa17;
assign Xwadt6 = Kksa17;
assign Hsr7z6[1] = Rnsa17;
assign P7s7z6[8] = Arsa17;
assign P7s7z6[9] = Tssa17;
assign P7s7z6[10] = Musa17;
assign P7s7z6[11] = Fwsa17;
assign P7s7z6[12] = Yxsa17;
assign P7s7z6[13] = Rzsa17;
assign P7s7z6[14] = K1ta17;
assign P7s7z6[16] = D3ta17;
assign P7s7z6[17] = W4ta17;
assign P7s7z6[18] = P6ta17;
assign P7s7z6[19] = I8ta17;
assign P7s7z6[20] = Cata17;
assign P7s7z6[21] = Wbta17;
assign P7s7z6[22] = Qdta17;
assign P7s7z6[24] = Kfta17;
assign P7s7z6[25] = Ehta17;
assign P7s7z6[26] = Yita17;
assign P7s7z6[27] = Skta17;
assign P7s7z6[28] = Mmta17;
assign P7s7z6[30] = Gota17;
assign Y26ft6 = Aqta17;
assign Jch7v6 = (!Trta17);
assign Gq37v6 = Qtta17;
assign I347v6 = Ivta17;
assign Fbxmz6[3] = Bxta17;
assign Ak77z6 = (!Yyta17);
assign Vcxmz6[0] = Q0ua17;
assign Vcxmz6[47] = L2ua17;
assign Vcxmz6[46] = H4ua17;
assign Vcxmz6[45] = D6ua17;
assign Vcxmz6[44] = Z7ua17;
assign Vcxmz6[43] = V9ua17;
assign Vcxmz6[42] = Rbua17;
assign Vcxmz6[41] = Ndua17;
assign Vcxmz6[40] = Jfua17;
assign Vcxmz6[39] = Fhua17;
assign Vcxmz6[38] = Bjua17;
assign Vcxmz6[37] = Xkua17;
assign Vcxmz6[36] = Tmua17;
assign Vcxmz6[35] = Poua17;
assign Vcxmz6[34] = Lqua17;
assign Vcxmz6[33] = Hsua17;
assign Vcxmz6[32] = Duua17;
assign Vcxmz6[31] = Zvua17;
assign Vcxmz6[30] = Vxua17;
assign Vcxmz6[29] = Rzua17;
assign Vcxmz6[28] = N1va17;
assign Vcxmz6[27] = J3va17;
assign Vcxmz6[26] = F5va17;
assign Vcxmz6[25] = B7va17;
assign Vcxmz6[24] = X8va17;
assign Vcxmz6[23] = Tava17;
assign Vcxmz6[22] = Pcva17;
assign Vcxmz6[21] = Leva17;
assign Vcxmz6[20] = Hgva17;
assign Vcxmz6[19] = Diva17;
assign Vcxmz6[18] = Zjva17;
assign Vcxmz6[17] = Vlva17;
assign Vcxmz6[16] = Rnva17;
assign Vcxmz6[15] = Npva17;
assign Vcxmz6[14] = Jrva17;
assign Vcxmz6[13] = Ftva17;
assign Vcxmz6[12] = Bvva17;
assign Vcxmz6[11] = Xwva17;
assign Vcxmz6[10] = Tyva17;
assign Vcxmz6[9] = P0wa17;
assign Vcxmz6[8] = K2wa17;
assign Vcxmz6[7] = F4wa17;
assign Vcxmz6[6] = A6wa17;
assign Vcxmz6[5] = V7wa17;
assign Vcxmz6[4] = Q9wa17;
assign Vcxmz6[3] = Lbwa17;
assign Vcxmz6[2] = Gdwa17;
assign Vcxmz6[1] = Bfwa17;
assign P647v6 = Wgwa17;
assign O9xmz6[0] = Oiwa17;
assign O9xmz6[2] = Mkwa17;
assign O9xmz6[1] = Kmwa17;
assign Fbxmz6[2] = Iowa17;
assign V147v6 = Fqwa17;
assign Oo1nz6[7] = Wrwa17;
assign Nn1nz6[7] = Utwa17;
assign Mm1nz6[7] = Svwa17;
assign Kh1nz6[7] = Qxwa17;
assign Vs27v6 = Ozwa17;
assign Ixr7z6[1] = K1xa17;
assign Ixr7z6[0] = M4xa17;
assign Uur7z6[1] = O7xa17;
assign Uur7z6[0] = Vaxa17;
assign Nw5ft6 = Cexa17;
assign Hsr7z6[0] = Jhxa17;
assign Enwmz6[0] = Skxa17;
assign Enwmz6[1] = Knxa17;
assign Mgwmz6[8] = Cqxa17;
assign Qiwmz6[8] = Nsxa17;
assign K5xmz6[0] = Yuxa17;
assign K5xmz6[1] = Qxxa17;
assign Sywmz6[8] = I0ya17;
assign W0xmz6[3] = T2ya17;
assign W0xmz6[2] = E5ya17;
assign W0xmz6[0] = P7ya17;
assign W0xmz6[8] = Aaya17;
assign Hwwmz6[0] = Lcya17;
assign Hwwmz6[1] = Dfya17;
assign Ppwmz6[8] = Vhya17;
assign Trwmz6[8] = Gkya17;
assign C4s7z6[0] = Rmya17;
assign Yr1nz6[3] = Vpya17;
assign Xq1nz6[3] = Trya17;
assign Xozmz6[4] = Rtya17;
assign Nqzmz6[4] = Ovya17;
assign Dszmz6[4] = Lxya17;
assign H80nz6[4] = Izya17;
assign X90nz6[4] = F1za17;
assign Nb0nz6[4] = C3za17;
assign Pyzmz6[4] = Z4za17;
assign F00nz6[4] = W6za17;
assign V10nz6[4] = T8za17;
assign Zh0nz6[4] = Qaza17;
assign Pj0nz6[4] = Ncza17;
assign Fl0nz6[4] = Keza17;
assign Ttzmz6[4] = Hgza17;
assign Jvzmz6[4] = Eiza17;
assign Zwzmz6[4] = Bkza17;
assign Dd0nz6[4] = Ylza17;
assign Te0nz6[4] = Vnza17;
assign Jg0nz6[4] = Spza17;
assign L30nz6[4] = Prza17;
assign B50nz6[4] = Mtza17;
assign R60nz6[4] = Jvza17;
assign Vm0nz6[4] = Gxza17;
assign Lo0nz6[4] = Dzza17;
assign Bq0nz6[4] = A10b17;
assign Ui67z6 = X20b17;
assign Au1nz6[4] = S40b17;
assign Zs1nz6[4] = Q60b17;
assign Yr1nz6[4] = O80b17;
assign Xq1nz6[4] = Ma0b17;
assign Xozmz6[6] = Kc0b17;
assign Nqzmz6[6] = He0b17;
assign Dszmz6[6] = Eg0b17;
assign H80nz6[6] = Bi0b17;
assign X90nz6[6] = Yj0b17;
assign Nb0nz6[6] = Vl0b17;
assign Ttzmz6[6] = Sn0b17;
assign Jvzmz6[6] = Pp0b17;
assign Zwzmz6[6] = Mr0b17;
assign Dd0nz6[6] = Jt0b17;
assign Te0nz6[6] = Gv0b17;
assign Jg0nz6[6] = Dx0b17;
assign Pyzmz6[6] = Az0b17;
assign F00nz6[6] = X01b17;
assign V10nz6[6] = U21b17;
assign Zh0nz6[6] = R41b17;
assign Pj0nz6[6] = O61b17;
assign Fl0nz6[6] = L81b17;
assign L30nz6[6] = Ia1b17;
assign B50nz6[6] = Fc1b17;
assign R60nz6[6] = Ce1b17;
assign Xozmz6[7] = Zf1b17;
assign Nqzmz6[7] = Wh1b17;
assign Dszmz6[7] = Tj1b17;
assign H80nz6[7] = Ql1b17;
assign X90nz6[7] = Nn1b17;
assign Nb0nz6[7] = Kp1b17;
assign Ttzmz6[7] = Hr1b17;
assign Jvzmz6[7] = Et1b17;
assign Dd0nz6[7] = Bv1b17;
assign Te0nz6[7] = Yw1b17;
assign Jg0nz6[7] = Vy1b17;
assign Pyzmz6[7] = S02b17;
assign F00nz6[7] = P22b17;
assign V10nz6[7] = M42b17;
assign Zh0nz6[7] = J62b17;
assign Pj0nz6[7] = G82b17;
assign Fl0nz6[7] = Da2b17;
assign L30nz6[7] = Ac2b17;
assign B50nz6[7] = Xd2b17;
assign R60nz6[7] = Uf2b17;
assign Vm0nz6[7] = Rh2b17;
assign Lo0nz6[7] = Oj2b17;
assign Bq0nz6[7] = Ll2b17;
assign Xozmz6[0] = In2b17;
assign Nqzmz6[0] = Fp2b17;
assign Dszmz6[0] = Cr2b17;
assign H80nz6[0] = Zs2b17;
assign X90nz6[0] = Wu2b17;
assign Nb0nz6[0] = Tw2b17;
assign Pyzmz6[0] = Qy2b17;
assign F00nz6[0] = N03b17;
assign V10nz6[0] = K23b17;
assign Zh0nz6[0] = H43b17;
assign Pj0nz6[0] = E63b17;
assign Fl0nz6[0] = B83b17;
assign Xozmz6[5] = Y93b17;
assign Nqzmz6[5] = Vb3b17;
assign Dszmz6[5] = Sd3b17;
assign H80nz6[5] = Pf3b17;
assign X90nz6[5] = Mh3b17;
assign Nb0nz6[5] = Jj3b17;
assign Pyzmz6[5] = Gl3b17;
assign F00nz6[5] = Dn3b17;
assign V10nz6[5] = Ap3b17;
assign Zh0nz6[5] = Xq3b17;
assign Pj0nz6[5] = Us3b17;
assign Fl0nz6[5] = Ru3b17;
assign Ttzmz6[5] = Ow3b17;
assign Jvzmz6[5] = Ly3b17;
assign Zwzmz6[5] = I04b17;
assign Dd0nz6[5] = F24b17;
assign Te0nz6[5] = C44b17;
assign Jg0nz6[5] = Z54b17;
assign L30nz6[5] = W74b17;
assign B50nz6[5] = T94b17;
assign R60nz6[5] = Qb4b17;
assign Vm0nz6[5] = Nd4b17;
assign Lo0nz6[5] = Kf4b17;
assign Bq0nz6[5] = Hh4b17;
assign Cj67z6 = Ej4b17;
assign Au1nz6[5] = Zk4b17;
assign Zs1nz6[5] = Xm4b17;
assign Yr1nz6[5] = Vo4b17;
assign Xq1nz6[5] = Tq4b17;
assign W94ft6 = Rs4b17;
assign Bxi7z6[2] = Pu4b17;
assign Hc2ft6 = Nw4b17;
assign Pnb7z6[24] = Uy4b17;
assign Dvc7z6[24] = X05b17;
assign Cgset6 = D45b17;
assign W3p7z6[24] = U55b17;
assign T2p7z6[24] = K75b17;
assign A0p7z6[22] = A95b17;
assign Hxo7z6[22] = Qa5b17;
assign Ouo7z6[22] = Gc5b17;
assign Vro7z6[22] = Wd5b17;
assign Nqo7z6[22] = Mf5b17;
assign Fpo7z6[22] = Ch5b17;
assign Bzi7z6[24] = Si5b17;
assign Wui7z6[24] = Sk5b17;
assign X9s7z6[32] = Um5b17;
assign K0wmz6[0] = Ro5b17;
assign Gyvmz6[0] = Cr5b17;
assign J7wmz6[0] = Nt5b17;
assign Qiwmz6[0] = Yv5b17;
assign Mgwmz6[0] = Jy5b17;
assign Trwmz6[0] = U06b17;
assign Ppwmz6[0] = F36b17;
assign E277z6 = (!Q56b17);
assign O177z6 = (!T86b17);
assign J0n7z6[0] = Wb6b17;
assign Pnb7z6[18] = Qe6b17;
assign Dvc7z6[18] = Tg6b17;
assign Isset6 = Zj6b17;
assign W3p7z6[18] = Ql6b17;
assign T2p7z6[18] = Gn6b17;
assign A0p7z6[16] = Wo6b17;
assign Hxo7z6[16] = Mq6b17;
assign Ouo7z6[16] = Cs6b17;
assign Vro7z6[16] = St6b17;
assign Nqo7z6[16] = Iv6b17;
assign Fpo7z6[16] = Yw6b17;
assign X9s7z6[26] = Oy6b17;
assign Pdc7z6[10] = L07b17;
assign Moj7z6[1] = M37b17;
assign Fjb7z6[2] = Q57b17;
assign Fjb7z6[66] = R67b17;
assign Fjb7z6[65] = T77b17;
assign Fjb7z6[4] = V87b17;
assign Fjb7z6[5] = W97b17;
assign Fjb7z6[6] = Xa7b17;
assign Fjb7z6[7] = Yb7b17;
assign Fjb7z6[9] = Zc7b17;
assign Fjb7z6[10] = Yg5m17;
assign Fjb7z6[11] = Ai5m17;
assign Fjb7z6[12] = Cj5m17;
assign Fjb7z6[13] = Ek5m17;
assign Fjb7z6[14] = Gl5m17;
assign Fjb7z6[15] = Im5m17;
assign Fjb7z6[16] = Kn5m17;
assign Fjb7z6[17] = Mo5m17;
assign Fjb7z6[19] = Op5m17;
assign Fjb7z6[20] = Qq5m17;
assign Fjb7z6[21] = Sr5m17;
assign Fjb7z6[22] = Us5m17;
assign Fjb7z6[23] = Wt5m17;
assign Fjb7z6[24] = Yu5m17;
assign Fjb7z6[25] = Aw5m17;
assign Fjb7z6[26] = Cx5m17;
assign Fjb7z6[27] = Ey5m17;
assign Fjb7z6[28] = Gz5m17;
assign Fjb7z6[29] = I06m17;
assign Fjb7z6[30] = K16m17;
assign Fjb7z6[31] = M26m17;
assign Fjb7z6[32] = O36m17;
assign Fjb7z6[33] = Q46m17;
assign Fjb7z6[34] = S56m17;
assign Fjb7z6[35] = U66m17;
assign Fjb7z6[36] = W76m17;
assign Fjb7z6[37] = Y86m17;
assign Fjb7z6[38] = Aa6m17;
assign Fjb7z6[39] = Cb6m17;
assign Fjb7z6[40] = Ec6m17;
assign Fjb7z6[41] = Gd6m17;
assign Fjb7z6[42] = Ie6m17;
assign Fjb7z6[43] = Kf6m17;
assign Fjb7z6[44] = Mg6m17;
assign Fjb7z6[45] = Oh6m17;
assign Fjb7z6[46] = Qi6m17;
assign Fjb7z6[47] = Sj6m17;
assign Fjb7z6[48] = Uk6m17;
assign Fjb7z6[49] = Wl6m17;
assign Fjb7z6[50] = Ym6m17;
assign Fjb7z6[51] = Ao6m17;
assign Fjb7z6[52] = Cp6m17;
assign Fjb7z6[53] = Eq6m17;
assign Fjb7z6[54] = Gr6m17;
assign Fjb7z6[55] = Is6m17;
assign Fjb7z6[56] = Kt6m17;
assign Fjb7z6[57] = Mu6m17;
assign Fjb7z6[59] = Ov6m17;
assign Fjb7z6[60] = Qw6m17;
assign Fjb7z6[61] = Sx6m17;
assign Fjb7z6[62] = Uy6m17;
assign Fjb7z6[63] = Wz6m17;
assign Fjb7z6[64] = Y07m17;
assign Fjb7z6[3] = A27m17;
assign Yr1nz6[7] = B37m17;
assign Xq1nz6[7] = Z47m17;
assign J72nz6[7] = X67m17;
assign Qc77z6 = (!Y87m17);
assign K1i7z6[12] = Fb7m17;
assign K1i7z6[20] = Je7m17;
assign Hhq7z6[3] = Nh7m17;
assign Hhq7z6[2] = Tj7m17;
assign Hhq7z6[1] = Zl7m17;
assign Hhq7z6[0] = Fo7m17;
assign Yr1nz6[6] = Lq7m17;
assign Xq1nz6[6] = Js7m17;
assign Bxi7z6[0] = Hu7m17;
assign Qubet6 = Fw7m17;
assign X9s7z6[15] = Jy7m17;
assign Bv37v6 = G08m17;
assign Xtwmz6[0] = N28m17;
assign Xtwmz6[1] = E58m17;
assign Cnvmz6[0] = V78m17;
assign Cnvmz6[8] = Ka8m17;
assign Kwvmz6[0] = Zc8m17;
assign A3xmz6[0] = Ye8m17;
assign A3xmz6[1] = Ph8m17;
assign Jt37v6 = Gk8m17;
assign Kms7z6[8] = Nm8m17;
assign Kwvmz6[1] = Cp8m17;
assign Kwvmz6[2] = Br8m17;
assign Kwvmz6[3] = At8m17;
assign Kwvmz6[4] = Zu8m17;
assign Tw37v6 = Yw8m17;
assign Ukwmz6[0] = Fz8m17;
assign Ukwmz6[1] = W19m17;
assign Xovmz6[0] = N49m17;
assign Xovmz6[8] = C79m17;
assign D047v6 = R99m17;
assign O2wmz6[0] = Yb9m17;
assign O2wmz6[1] = Pe9m17;
assign Nsvmz6[0] = Gh9m17;
assign Rbwmz6[0] = Vj9m17;
assign Rbwmz6[1] = Mm9m17;
assign N9wmz6[0] = Dp9m17;
assign Sqvmz6[0] = Or9m17;
assign N9wmz6[8] = Du9m17;
assign Sqvmz6[8] = Ow9m17;
assign Vitet6 = Dz9m17;
assign W3p7z6[5] = T0am17;
assign T2p7z6[5] = I2am17;
assign A0p7z6[3] = X3am17;
assign Hxo7z6[3] = M5am17;
assign Ouo7z6[3] = B7am17;
assign Vro7z6[3] = Q8am17;
assign Nqo7z6[3] = Faam17;
assign Fpo7z6[3] = Ubam17;
assign Pdq7z6[5] = Jdam17;
assign Cjq7z6[5] = Pfam17;
assign X9s7z6[13] = Vham17;
assign K1i7z6[21] = Sjam17;
assign X9s7z6[37] = Wmam17;
assign Hhq7z6[7] = Toam17;
assign V1s7z6[1] = Zqam17;
assign Cjq7z6[6] = Ntam17;
assign X9s7z6[14] = Tvam17;
assign K1i7z6[22] = Qxam17;
assign Pdq7z6[7] = U0bm17;
assign V1s7z6[3] = A3bm17;
assign X9s7z6[28] = O5bm17;
assign X9s7z6[20] = L7bm17;
assign W0xmz6[4] = I9bm17;
assign Sywmz6[4] = Tbbm17;
assign Kms7z6[4] = Eebm17;
assign Trwmz6[4] = Tgbm17;
assign Ppwmz6[4] = Ejbm17;
assign Cnvmz6[4] = Plbm17;
assign Qiwmz6[4] = Eobm17;
assign Mgwmz6[4] = Pqbm17;
assign Xovmz6[4] = Atbm17;
assign N9wmz6[4] = Pvbm17;
assign J7wmz6[4] = Aybm17;
assign Sqvmz6[4] = L0cm17;
assign Pdc7z6[20] = A3cm17;
assign Dvc7z6[20] = B6cm17;
assign Kxb7z6[11] = H9cm17;
assign Fth7z6[11] = Rbcm17;
assign X9s7z6[35] = Pecm17;
assign vis_r1_o[31] = Mgcm17;
assign vis_r2_o[31] = Djcm17;
assign vis_r3_o[31] = Ulcm17;
assign vis_r4_o[31] = Locm17;
assign vis_r5_o[31] = Crcm17;
assign vis_r6_o[31] = Ttcm17;
assign vis_r7_o[31] = Kwcm17;
assign vis_r8_o[31] = Bzcm17;
assign vis_r9_o[31] = S1dm17;
assign vis_r10_o[31] = J4dm17;
assign vis_r11_o[31] = B7dm17;
assign vis_r12_o[31] = T9dm17;
assign vis_msp_o[31] = Lcdm17;
assign Pic7z6[31] = Dfdm17;
assign vis_psp_o[31] = Vhdm17;
assign vis_r0_o[31] = Nkdm17;
assign Fjb7z6[1] = Endm17;
assign K1i7z6[9] = Fodm17;
assign X9s7z6[33] = Irdm17;
assign K1i7z6[17] = Ftdm17;
assign Pnb7z6[22] = Jwdm17;
assign Ekset6 = Mydm17;
assign W3p7z6[22] = D0em17;
assign T2p7z6[22] = T1em17;
assign A0p7z6[20] = J3em17;
assign Hxo7z6[20] = Z4em17;
assign Ouo7z6[20] = P6em17;
assign Vro7z6[20] = F8em17;
assign Nqo7z6[20] = V9em17;
assign Fpo7z6[20] = Lbem17;
assign Wui7z6[22] = Bdem17;
assign X9s7z6[30] = Dfem17;
assign W0xmz6[6] = Ahem17;
assign Sywmz6[6] = Ljem17;
assign Kms7z6[6] = Wlem17;
assign Trwmz6[6] = Loem17;
assign Ppwmz6[6] = Wqem17;
assign Cnvmz6[6] = Htem17;
assign Qiwmz6[6] = Wvem17;
assign Mgwmz6[6] = Hyem17;
assign Xovmz6[6] = S0fm17;
assign N9wmz6[6] = H3fm17;
assign J7wmz6[6] = S5fm17;
assign Sqvmz6[6] = D8fm17;
assign Pdc7z6[22] = Safm17;
assign Dvc7z6[22] = Tdfm17;
assign Byc7z6[29] = Zgfm17;
assign Wlr7z6[23] = Dkfm17;
assign Wlr7z6[15] = Rmfm17;
assign Wlr7z6[7] = Fpfm17;
assign W0xmz6[7] = Srfm17;
assign Sywmz6[7] = Dufm17;
assign Kms7z6[7] = Owfm17;
assign Trwmz6[7] = Dzfm17;
assign Ppwmz6[7] = O1gm17;
assign Cnvmz6[7] = Z3gm17;
assign Qiwmz6[7] = O6gm17;
assign Mgwmz6[7] = Z8gm17;
assign Xovmz6[7] = Kbgm17;
assign N9wmz6[7] = Zdgm17;
assign J7wmz6[7] = Kggm17;
assign Sqvmz6[7] = Vigm17;
assign K1i7z6[31] = Klgm17;
assign X9s7z6[9] = Oogm17;
assign K1i7z6[25] = Kqgm17;
assign X9s7z6[17] = Otgm17;
assign Pdc7z6[0] = Lvgm17;
assign Pdc7z6[31] = Lygm17;
assign Fjb7z6[58] = M1hm17;
assign Fjb7z6[18] = O2hm17;
assign Fjb7z6[8] = Q3hm17;
assign X9s7z6[18] = R4hm17;
assign K0wmz6[2] = O6hm17;
assign Gyvmz6[2] = Z8hm17;
assign Nsvmz6[2] = Kbhm17;
assign N9wmz6[2] = Zdhm17;
assign J7wmz6[2] = Kghm17;
assign Sqvmz6[2] = Vihm17;
assign Qiwmz6[2] = Klhm17;
assign Mgwmz6[2] = Vnhm17;
assign Xovmz6[2] = Gqhm17;
assign Trwmz6[2] = Vshm17;
assign Ppwmz6[2] = Gvhm17;
assign Cnvmz6[2] = Rxhm17;
assign Oyh7z6[1] = G0im17;
assign K1i7z6[26] = J3im17;
assign Kh1nz6[2] = N6im17;
assign J72nz6[2] = L8im17;
assign Pnb7z6[19] = Maim17;
assign Dvc7z6[19] = Pcim17;
assign Hqset6 = Vfim17;
assign W3p7z6[19] = Mhim17;
assign T2p7z6[19] = Cjim17;
assign A0p7z6[17] = Skim17;
assign Hxo7z6[17] = Imim17;
assign Ouo7z6[17] = Ynim17;
assign Vro7z6[17] = Opim17;
assign Nqo7z6[17] = Erim17;
assign Fpo7z6[17] = Usim17;
assign X9s7z6[27] = Kuim17;
assign K0wmz6[3] = Hwim17;
assign Gyvmz6[3] = Syim17;
assign Nsvmz6[3] = D1jm17;
assign N9wmz6[3] = S3jm17;
assign J7wmz6[3] = D6jm17;
assign Sqvmz6[3] = O8jm17;
assign Qiwmz6[3] = Dbjm17;
assign Mgwmz6[3] = Odjm17;
assign Xovmz6[3] = Zfjm17;
assign Trwmz6[3] = Oijm17;
assign Ppwmz6[3] = Zkjm17;
assign Cnvmz6[3] = Knjm17;
assign Kh1nz6[3] = Zpjm17;
assign J72nz6[3] = Xrjm17;
assign Pdc7z6[3] = Ytjm17;
assign Dvc7z6[3] = Ywjm17;
assign Byc7z6[24] = D0km17;
assign Xmtet6 = H3km17;
assign Yotet6 = A5km17;
assign Gsb7z6[0] = T6km17;
assign Gsb7z6[1] = M8km17;
assign Ozadt6 = Fakm17;
assign Y9pet6 = Wbkm17;
assign X7pet6 = Pdkm17;
assign V3pet6 = Ifkm17;
assign Wktet6 = Fhkm17;
assign Wui7z6[21] = Yikm17;
assign X9s7z6[29] = Alkm17;
assign X9s7z6[21] = Xmkm17;
assign W0xmz6[5] = Uokm17;
assign Sywmz6[5] = Frkm17;
assign Kms7z6[5] = Qtkm17;
assign Trwmz6[5] = Fwkm17;
assign Ppwmz6[5] = Qykm17;
assign Cnvmz6[5] = B1lm17;
assign Qiwmz6[5] = Q3lm17;
assign Mgwmz6[5] = B6lm17;
assign Xovmz6[5] = M8lm17;
assign N9wmz6[5] = Bblm17;
assign J7wmz6[5] = Mdlm17;
assign Sqvmz6[5] = Xflm17;
assign K0wmz6[5] = Milm17;
assign Gyvmz6[5] = Xklm17;
assign Nsvmz6[5] = Inlm17;
assign V7xmz6[5] = Xplm17;
assign Kh1nz6[5] = Xrlm17;
assign J72nz6[5] = Vtlm17;
assign Eqn7z6[0] = Wvlm17;
assign Eqn7z6[2] = Xylm17;
assign Eqn7z6[1] = Y1mm17;
assign Dvc7z6[4] = Z4mm17;
assign D5f7z6[2] = E8mm17;
assign D5f7z6[0] = Abmm17;
assign D5f7z6[1] = Wdmm17;
assign W2n7z6[0] = Sgmm17;
assign J5n7z6[2] = Mjmm17;
assign G4i7z6[0] = Cmmm17;
assign Oyh7z6[2] = Xomm17;
assign G4i7z6[1] = Asmm17;
assign Oyh7z6[3] = Vumm17;
assign G4i7z6[2] = Yxmm17;
assign Oyh7z6[4] = T0nm17;
assign G4i7z6[3] = W3nm17;
assign G4i7z6[4] = R6nm17;
assign Oyh7z6[6] = M9nm17;
assign G4i7z6[5] = Pcnm17;
assign Oyh7z6[7] = Kfnm17;
assign G4i7z6[6] = Ninm17;
assign Oyh7z6[8] = Ilnm17;
assign G4i7z6[7] = Lonm17;
assign Oyh7z6[9] = Grnm17;
assign G4i7z6[8] = Junm17;
assign Oyh7z6[10] = Exnm17;
assign G4i7z6[9] = I0om17;
assign Oyh7z6[11] = D3om17;
assign Oyh7z6[12] = H6om17;
assign Oyh7z6[13] = L9om17;
assign Oyh7z6[14] = Pcom17;
assign Oyh7z6[15] = Tfom17;
assign Oyh7z6[16] = Xiom17;
assign Oyh7z6[17] = Bmom17;
assign Oyh7z6[18] = Fpom17;
assign Oyh7z6[19] = Jsom17;
assign Oyh7z6[20] = Nvom17;
assign Oyh7z6[21] = Ryom17;
assign Oyh7z6[22] = V1pm17;
assign Oyh7z6[23] = Z4pm17;
assign Oyh7z6[24] = D8pm17;
assign Oyh7z6[25] = Hbpm17;
assign Oyh7z6[26] = Lepm17;
assign Oyh7z6[27] = Phpm17;
assign Oyh7z6[28] = Tkpm17;
assign Oyh7z6[29] = Xnpm17;
assign Oyh7z6[30] = Brpm17;
assign Oyh7z6[31] = Fupm17;
assign Oyh7z6[0] = Jxpm17;
assign Byc7z6[0] = M0qm17;
assign Ryadt6 = P3qm17;
assign Oo1nz6[0] = A5qm17;
assign J72nz6[0] = Y6qm17;
assign N52nz6[6] = Z8qm17;
assign N52nz6[5] = Xaqm17;
assign N52nz6[4] = Wcqm17;
assign N52nz6[3] = Veqm17;
assign N52nz6[2] = Ugqm17;
assign N52nz6[1] = Tiqm17;
assign N52nz6[0] = Skqm17;
assign Wye7v6 = Rmqm17;
assign Z12nz6[2] = Qoqm17;
assign Z12nz6[3] = Rqqm17;
assign Z12nz6[5] = Ssqm17;
assign Z12nz6[7] = Tuqm17;
assign TRACEDATA[3] = Uwqm17;
assign Oih7v6 = (!Uwqm17);
assign Z12nz6[0] = Syqm17;
assign X9s7z6[25] = T0rm17;
assign K0wmz6[1] = Q2rm17;
assign Gyvmz6[1] = B5rm17;
assign Nsvmz6[1] = M7rm17;
assign N9wmz6[1] = Barm17;
assign J7wmz6[1] = Mcrm17;
assign Sqvmz6[1] = Xerm17;
assign Qiwmz6[1] = Mhrm17;
assign Mgwmz6[1] = Xjrm17;
assign Xovmz6[1] = Imrm17;
assign Trwmz6[1] = Xorm17;
assign Ppwmz6[1] = Irrm17;
assign Cnvmz6[1] = Ttrm17;
assign W0xmz6[1] = Iwrm17;
assign Sywmz6[1] = Tyrm17;
assign Kms7z6[1] = E1sm17;
assign T5fet6 = T3sm17;
assign HTMDHTRANS[1] = V5sm17;
assign Dgh7v6 = (!V5sm17);
assign Fb47v6 = N7sm17;
assign V947v6 = A9sm17;
assign Oyh7z6[5] = Oasm17;
assign Byc7z6[7] = Rdsm17;
assign R7fet6 = Ugsm17;
assign W5pet6 = Ajsm17;
assign J5n7z6[3] = Tksm17;
assign J0n7z6[1] = Jnsm17;
assign U1pet6 = Dqsm17;
assign W2n7z6[1] = Assm17;
assign S7f7z6[0] = Uusm17;
assign S7f7z6[2] = Sxsm17;
assign S7f7z6[5] = Q0tm17;
assign S7f7z6[1] = O3tm17;
assign S7f7z6[3] = M6tm17;
assign S7f7z6[4] = K9tm17;
assign Fre7z6[1] = Ictm17;
assign Kh1nz6[4] = Fftm17;
assign J72nz6[4] = Dhtm17;
assign Z12nz6[4] = Ejtm17;
assign Hjn7z6[7] = Fltm17;
assign Hjn7z6[8] = Vntm17;
assign Hjn7z6[9] = Lqtm17;
assign Hjn7z6[10] = Bttm17;
assign Hjn7z6[11] = Svtm17;
assign Hjn7z6[12] = Jytm17;
assign Hjn7z6[13] = A1um17;
assign Hjn7z6[14] = R3um17;
assign Hjn7z6[15] = I6um17;
assign Hjn7z6[16] = Z8um17;
assign Hjn7z6[17] = Qbum17;
assign Hjn7z6[18] = Heum17;
assign Hjn7z6[19] = Ygum17;
assign Hjn7z6[20] = Pjum17;
assign Hjn7z6[21] = Gmum17;
assign Hjn7z6[22] = Xoum17;
assign Hjn7z6[23] = Orum17;
assign Hjn7z6[24] = Fuum17;
assign Hjn7z6[25] = Wwum17;
assign Hjn7z6[26] = Nzum17;
assign Hjn7z6[27] = E2vm17;
assign Hjn7z6[28] = V4vm17;
assign Hjn7z6[29] = M7vm17;
assign Hjn7z6[30] = Davm17;
assign Hjn7z6[31] = Ucvm17;
assign X9s7z6[39] = Lfvm17;
assign Kh1nz6[6] = Ihvm17;
assign J72nz6[6] = Gjvm17;
assign Z12nz6[6] = Hlvm17;
assign TRACEDATA[2] = Invm17;
assign Hih7v6 = (!Invm17);
assign Byc7z6[31] = Gpvm17;
assign Cxtet6 = Ksvm17;
assign Bvtet6 = Duvm17;
assign Attet6 = Wvvm17;
assign Zqtet6 = Pxvm17;
assign Dztet6 = Izvm17;
assign Fopet6 = B1wm17;
assign Empet6 = U2wm17;
assign Dkpet6 = N4wm17;
assign Cipet6 = G6wm17;
assign Bgpet6 = Z7wm17;
assign Aepet6 = W9wm17;
assign J72nz6[1] = Tbwm17;
assign Z12nz6[1] = Udwm17;
assign TRACEDATA[1] = Vfwm17;
assign Vih7v6 = (!Vfwm17);
assign TRACEDATA[0] = Thwm17;
assign Aih7v6 = (!Thwm17);
assign SWV = Rjwm17;
assign H1m8v6 = (Hsi7z6[2] ? X5m8v6 : 1'b1);
assign Zyl8v6 = (Hsi7z6[2] ? Kja7z6 : 1'b1);
assign Rwl8v6 = (Hsi7z6[2] ? P3m8v6 : 1'b1);
assign X5m8v6 = (Hsi7z6[1] ? Sja7z6 : 1'b1);
assign Dpo8v6 = (O7c7z6[8] ? B9r8v6 : Ffr8v6);
assign Bmo8v6 = (O7c7z6[8] ? Z5r8v6 : Dcr8v6);
assign Zio8v6 = (O7c7z6[8] ? X2r8v6 : B9r8v6);
assign Xfo8v6 = (O7c7z6[8] ? Vzq8v6 : Z5r8v6);
assign Vco8v6 = (O7c7z6[8] ? Twq8v6 : X2r8v6);
assign T9o8v6 = (O7c7z6[8] ? Rtq8v6 : Vzq8v6);
assign R6o8v6 = (O7c7z6[8] ? Pqq8v6 : Twq8v6);
assign P3o8v6 = (O7c7z6[8] ? Nnq8v6 : Rtq8v6);
assign N0o8v6 = (O7c7z6[8] ? Lkq8v6 : Pqq8v6);
assign Lxn8v6 = (O7c7z6[8] ? Jhq8v6 : Nnq8v6);
assign Jun8v6 = (O7c7z6[8] ? Heq8v6 : Lkq8v6);
assign Hrn8v6 = (O7c7z6[8] ? Fbq8v6 : Jhq8v6);
assign Fon8v6 = (O7c7z6[8] ? D8q8v6 : Heq8v6);
assign Dln8v6 = (O7c7z6[8] ? B5q8v6 : Fbq8v6);
assign Bin8v6 = (O7c7z6[8] ? Z1q8v6 : D8q8v6);
assign Zen8v6 = (O7c7z6[8] ? Xyp8v6 : B5q8v6);
assign Xbn8v6 = (O7c7z6[8] ? Vvp8v6 : Z1q8v6);
assign V8n8v6 = (O7c7z6[8] ? Tsp8v6 : Xyp8v6);
assign T5n8v6 = (O7c7z6[8] ? Rpp8v6 : Vvp8v6);
assign R2n8v6 = (O7c7z6[8] ? Pmp8v6 : Tsp8v6);
assign Pzm8v6 = (O7c7z6[8] ? Ojp8v6 : Rpp8v6);
assign Nwm8v6 = (O7c7z6[8] ? Ngp8v6 : Pmp8v6);
assign Mtm8v6 = (O7c7z6[8] ? Mdp8v6 : Ojp8v6);
assign Lqm8v6 = (O7c7z6[8] ? Lap8v6 : Ngp8v6);
assign Knm8v6 = (O7c7z6[8] ? K7p8v6 : Mdp8v6);
assign Jkm8v6 = (O7c7z6[8] ? J4p8v6 : Lap8v6);
assign Ihm8v6 = (O7c7z6[8] ? I1p8v6 : K7p8v6);
assign Hem8v6 = (O7c7z6[8] ? Hyo8v6 : J4p8v6);
assign Gbm8v6 = (O7c7z6[8] ? Gvo8v6 : I1p8v6);
assign F8m8v6 = (O7c7z6[8] ? Fso8v6 : Hyo8v6);
assign Ffr8v6 = (O7c7z6[7] ? Zkh7z6[30] : Zkh7z6[31]);
assign Dcr8v6 = (O7c7z6[7] ? Zkh7z6[29] : Zkh7z6[30]);
assign B9r8v6 = (O7c7z6[7] ? Zkh7z6[28] : Zkh7z6[29]);
assign Z5r8v6 = (O7c7z6[7] ? Zkh7z6[27] : Zkh7z6[28]);
assign X2r8v6 = (O7c7z6[7] ? Zkh7z6[26] : Zkh7z6[27]);
assign Vzq8v6 = (O7c7z6[7] ? Zkh7z6[25] : Zkh7z6[26]);
assign Twq8v6 = (O7c7z6[7] ? Zkh7z6[24] : Zkh7z6[25]);
assign Rtq8v6 = (O7c7z6[7] ? Zkh7z6[23] : Zkh7z6[24]);
assign Pqq8v6 = (O7c7z6[7] ? Zkh7z6[22] : Zkh7z6[23]);
assign Nnq8v6 = (O7c7z6[7] ? Zkh7z6[21] : Zkh7z6[22]);
assign Lkq8v6 = (O7c7z6[7] ? Zkh7z6[20] : Zkh7z6[21]);
assign Jhq8v6 = (O7c7z6[7] ? Zkh7z6[19] : Zkh7z6[20]);
assign Heq8v6 = (O7c7z6[7] ? Zkh7z6[18] : Zkh7z6[19]);
assign Fbq8v6 = (O7c7z6[7] ? Zkh7z6[17] : Zkh7z6[18]);
assign D8q8v6 = (O7c7z6[7] ? Zkh7z6[16] : Zkh7z6[17]);
assign B5q8v6 = (O7c7z6[7] ? Zkh7z6[15] : Zkh7z6[16]);
assign Z1q8v6 = (O7c7z6[7] ? Zkh7z6[14] : Zkh7z6[15]);
assign Xyp8v6 = (O7c7z6[7] ? Zkh7z6[13] : Zkh7z6[14]);
assign Vvp8v6 = (O7c7z6[7] ? Zkh7z6[12] : Zkh7z6[13]);
assign Tsp8v6 = (O7c7z6[7] ? Zkh7z6[11] : Zkh7z6[12]);
assign Rpp8v6 = (O7c7z6[7] ? Zkh7z6[10] : Zkh7z6[11]);
assign Pmp8v6 = (O7c7z6[7] ? Zkh7z6[9] : Zkh7z6[10]);
assign Ojp8v6 = (O7c7z6[7] ? Zkh7z6[8] : Zkh7z6[9]);
assign Ngp8v6 = (O7c7z6[7] ? Zkh7z6[7] : Zkh7z6[8]);
assign Mdp8v6 = (O7c7z6[7] ? Zkh7z6[6] : Zkh7z6[7]);
assign Lap8v6 = (O7c7z6[7] ? Zkh7z6[5] : Zkh7z6[6]);
assign K7p8v6 = (O7c7z6[7] ? Zkh7z6[4] : Zkh7z6[5]);
assign J4p8v6 = (O7c7z6[7] ? Zkh7z6[3] : Zkh7z6[4]);
assign I1p8v6 = (O7c7z6[7] ? Zkh7z6[2] : Zkh7z6[3]);
assign Hyo8v6 = (O7c7z6[7] ? Zkh7z6[1] : Zkh7z6[2]);
assign Gvo8v6 = (O7c7z6[7] ? Zkh7z6[0] : Zkh7z6[1]);
assign Q1s8v6 = (Bat8v6 ? Nas8v6 : Jms8v6);
assign Ryr8v6 = (Bat8v6 ? O7s8v6 : Kjs8v6);
assign Svr8v6 = (Bat8v6 ? P4s8v6 : Lgs8v6);
assign Tsr8v6 = (Bat8v6 ? 1'b0 : Mds8v6);
assign Jms8v6 = (Kfa7z6 ? Fys8v6 : D4t8v6);
assign Kjs8v6 = (Kfa7z6 ? Gvs8v6 : E1t8v6);
assign Lgs8v6 = (Kfa7z6 ? Hss8v6 : Fys8v6);
assign Mds8v6 = (Kfa7z6 ? Ips8v6 : Gvs8v6);
assign Nas8v6 = (Kfa7z6 ? C7t8v6 : Hss8v6);
assign O7s8v6 = (Kfa7z6 ? 1'b0 : Ips8v6);
assign D4t8v6 = (Sfa7z6 ? Uqd7z6[21] : Uqd7z6[22]);
assign E1t8v6 = (Sfa7z6 ? Uqd7z6[20] : Uqd7z6[21]);
assign Fys8v6 = (Sfa7z6 ? Uqd7z6[19] : Uqd7z6[20]);
assign Gvs8v6 = (Sfa7z6 ? Uqd7z6[18] : Uqd7z6[19]);
assign Hss8v6 = (Sfa7z6 ? Uqd7z6[17] : Uqd7z6[18]);
assign Ips8v6 = (Sfa7z6 ? Ovbdt6 : Uqd7z6[17]);
assign {D9f7v6, Naf7v6, Xbf7v6, Hdf7v6, Ref7v6, Bgf7v6, Lhf7v6, Vif7v6,
 Fkf7v6, Plf7v6, Zmf7v6, Jof7v6, Tpf7v6} = (Td2nz6 + 1'b1);
assign {Bmd7v6, Lnd7v6, Vod7v6, Fqd7v6, Prd7v6, Zsd7v6, Jud7v6, Tvd7v6,
 Dxd7v6} = (H71nz6 - 1'b1);
assign Llwm17 = ({E11nz6, 1'b0} + {{1'b0, Rht8v6, Bgt8v6, Let8v6,
 Wsc7v6}, 1'b1});
assign {Mz0nz6, Ux0nz6} = Llwm17[33:1];
assign Cnwm17 = ({{G0d7v6, M1d7v6, S2d7v6, Y3d7v6, E5d7v6}, 1'b0} +
 {E11nz6, 1'b1});
assign {Cuc7v6, Ivc7v6, Owc7v6, Uxc7v6, Azc7v6} = Cnwm17[33:1];
assign Towm17 = ((E11nz6 - {Rr0nz6, Hw0nz6, E5d7v6}) - 1'b0);
assign {K6d7v6, Q7d7v6, W8d7v6, Cad7v6, Ibd7v6} = Towm17[4:0];
assign Jqwm17 = ({Slzmz6, 1'b0} + {{1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, W9c7v6}, 1'b1});
assign {Uq87v6, Ds87v6, Mt87v6, Vu87v6, Ew87v6, Nx87v6, Wy87v6, F097v6,
 O197v6, X297v6, G497v6, P597v6, Y697v6, H897v6, Q997v6, Za97v6,
 Ic97v6, Rd97v6, Af97v6, Jg97v6, Sh97v6, Bj97v6, Kk97v6, Tl97v6,
 Cn97v6, Lo97v6, Up97v6, Dr97v6, Ms97v6, Vt97v6, Ev97v6} =
 Jqwm17[33:1];
assign Ctymz6 = (Ruymz6 - 1'b1);
assign {Ub67v6, Uc67v6, Ud67v6, Ue67v6, Uf67v6, Ug67v6, Uh67v6, Ui67v6,
 Uj67v6, Uk67v6, Ul67v6, Um67v6} = (Hnxmz6 - 1'b1);
assign {Iw27v6, Px27v6, Wy27v6, D037v6, K137v6, R237v6, Y337v6, F537v6,
 M637v6, T737v6, A937v6, Ha37v6, Ob37v6, Vc37v6, Ce37v6, Jf37v6,
 Qg37v6, Xh37v6, Ej37v6, Lk37v6, Sl37v6} = ({P7s7z6[30:24],
 P7s7z6[22:16], P7s7z6[14:8]} + 1'b1);
assign Em5ft6 = (({Mkp7z6[31:15], S8r7z6} == {T6r7z6[31:16], Ve5ft6,
 T6r7z6[14:1], 1'b0}) ? 1'b1 : 1'b0);
assign Gb5ft6 = (({Bqp7z6[31:15], O2r7z6} == {T6r7z6[31:16], Ve5ft6,
 P0r7z6, 1'b0}) ? 1'b1 : 1'b0);
assign X15ft6 = (({B2q7z6[31:15], Kwq7z6} == {T6r7z6[31:16], Ve5ft6,
 Luq7z6, 1'b0}) ? 1'b1 : 1'b0);
assign Mq4ft6 = (({E6p7z6[31:15], Gqq7z6} == {T6r7z6[31:16], Ve5ft6,
 Hoq7z6, 1'b0}) ? 1'b1 : 1'b0);
assign {I03ft6, T13ft6, E33ft6, P43ft6, A63ft6, L73ft6, W83ft6, Ha3ft6,
 Sb3ft6, Dd3ft6, Oe3ft6, Zf3ft6, Kh3ft6, Vi3ft6, Gk3ft6, Rl3ft6,
 Cn3ft6, No3ft6, Yp3ft6, Jr3ft6, Us3ft6, Fu3ft6, Qv3ft6, Bx3ft6,
 My3ft6, Xz3ft6, I14ft6, T24ft6, E44ft6, P54ft6, A74ft6, L84ft6}
 = (U9p7z6 + 1'b1);
assign Zb1ft6 = (({1'b0, 1'b0, 1'b0, Fpo7z6} == Zmo7z6) ? 1'b1 : 1'b0);
assign Xc1ft6 = (({1'b0, 1'b0, 1'b0, Nqo7z6} == Zmo7z6) ? 1'b1 : 1'b0);
assign Vd1ft6 = (({1'b0, 1'b0, 1'b0, Vro7z6} == Coo7z6) ? 1'b1 : 1'b0);
assign Te1ft6 = (({1'b0, 1'b0, 1'b0, Ouo7z6} == Coo7z6) ? 1'b1 : 1'b0);
assign Rf1ft6 = (({1'b0, 1'b0, 1'b0, Hxo7z6} == Coo7z6) ? 1'b1 : 1'b0);
assign Pg1ft6 = (({1'b0, 1'b0, 1'b0, A0p7z6} == Coo7z6) ? 1'b1 : 1'b0);
assign Nh1ft6 = (({1'b0, 1'b0, 1'b0, T2p7z6} == Coo7z6) ? 1'b1 : 1'b0);
assign Li1ft6 = (({1'b0, 1'b0, 1'b0, W3p7z6} == Coo7z6) ? 1'b1 : 1'b0);
assign Dswm17 = ({{U3o7z6[11:4], Y9o7z6}, 1'b0} + {{1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, O7o7z6}, 1'b1});
assign {Pxzet6, Pzzet6, P10ft6, P30ft6, P50ft6, P70ft6, P90ft6, Pb0ft6,
 Pd0ft6, Pf0ft6, Ph0ft6, Pj0ft6} = Dswm17[33:1];
assign Puwm17 = ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, Kvxet6} << {Ean7z6, Ryyet6, S0zet6, T2zet6});
assign {Y8uet6, Zauet6, Aduet6, Bfuet6, Chuet6, Djuet6, Eluet6, Fnuet6,
 Gpuet6, Hruet6, Ituet6, Jvuet6, Kxuet6, Lzuet6, M1vet6, N3vet6,
 O5vet6, P7vet6, Q9vet6, Rbvet6, Sdvet6, Tfvet6, Uhvet6, Vjvet6,
 Wlvet6, Xnvet6, Ypvet6, Zrvet6, Auvet6, Bwvet6, Cyvet6, D0wet6}
 = Puwm17[31:0];
assign Dxwm17 = ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b1} << {Ean7z6, Ryyet6, S0zet6, T2zet6});
assign {E2wet6, F4wet6, G6wet6, H8wet6, Iawet6, Jcwet6, Kewet6, Lgwet6,
 Miwet6, Nkwet6, Omwet6, Powet6, Qqwet6, Rswet6, Suwet6, Twwet6,
 Uywet6, V0xet6, W2xet6, X4xet6, Y6xet6, Z8xet6, Abxet6, Bdxet6,
 Cfxet6, Dhxet6, Ejxet6, Flxet6, Gnxet6, Hpxet6, Irxet6, Jtxet6}
 = Dxwm17[31:0];
assign Rzwm17 = ({Chn7z6, 1'b0} + {{1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, M7yet6, 1'b0, 1'b0}, 1'b1});
assign Icn7z6 = Rzwm17[33:1];
assign H2xm17 = ({N3k7z6, 1'b0} + {{1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, Obo7v6}, 1'b1});
assign {X0k7z6, Aka7z6, Xka7z6, Ula7z6} = H2xm17[33:1];
assign P9get6 = (({Tib7z6, M5bdt6, Oqbet6, Zrbet6, Qmj7z6[5:4], E6a7z6,
 Pnfet6, Qmj7z6[1], S3a7z6} != Jqj7z6) ? 1'b1 : 1'b0);
assign Fs4ft6 = (({E6p7z6[31:15], Gqq7z6} == {Gsq7z6[31:16], Bu4ft6,
 Gsq7z6[14:0]}) ? 1'b1 : 1'b0);
assign Q35ft6 = (({B2q7z6[31:15], Kwq7z6} == {Sar7z6[31:16], Tp5ft6,
 Kyq7z6}) ? 1'b1 : 1'b0);
assign Zc5ft6 = (({Bqp7z6[31:15], O2r7z6} == {Sar7z6[31:16], Tp5ft6,
 O4r7z6}) ? 1'b1 : 1'b0);
assign Xn5ft6 = (({Mkp7z6[31:15], S8r7z6} == {Sar7z6[31:16], Tp5ft6,
 Sar7z6[14:0]}) ? 1'b1 : 1'b0);
assign {Emcet6, Sncet6, Gpcet6, Uqcet6, Iscet6, Wtcet6, Kvcet6, Ywcet6,
 Mycet6, A0det6, O1det6, C3det6, Q4det6, E6det6, S7det6, G9det6,
 Uadet6, Icdet6, Wddet6, Kfdet6, Ygdet6, Midet6, Akdet6, Oldet6}
 = (A0j7z6 - 1'b1);
assign W4xm17 = ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, T9fet6} << {Bmfet6, Nkfet6, Zifet6,
 Lhfet6, Xffet6, Jefet6, Vcfet6, Hbfet6});
assign Qkj7z6 = W4xm17[63:0];
assign Y6xm17 = ((vis_pc_o - {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b1, 1'b0}) - 1'b0);
assign Bni7z6 = Y6xm17[30:0];
assign A9xm17 = ((vis_pc_o - {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, Zei7z6}) - 1'b0);
assign Gli7z6 = A9xm17[30:0];
assign Cbxm17 = ({vis_pc_o, 1'b0} + {{1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, A4a7z6, Tao7v6}, 1'b1});
assign Bhi7z6 = Cbxm17[33:1];
assign Edxm17 = ({{Wt97z6, Eu97z6, Cv97z6, Uu97z6, Sv97z6, Qw97z6,
 Ox97z6, Wx97z6, Ey97z6, My97z6, Uy97z6, Cz97z6, Kz97z6, Yw97z6,
 Sz97z6, A0a7z6, Kv97z6, I0a7z6, Q0a7z6, Y0a7z6, G1a7z6, Gx97z6,
 O1a7z6, Aw97z6, W1a7z6, E2a7z6, M2a7z6, Iw97z6, U2a7z6, As97z6,
 Mu97z6}, 1'b0} + {{1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b1, 1'b0}, 1'b1});
assign Eji7z6 = Edxm17[33:1];
assign Gfxm17 = ({{Ca3et6, Lc3et6, Ue3et6, Dh3et6, Mj3et6, Vl3et6,
 Eo3et6, Nq3et6, Ws3et6, Fv3et6, Ox3et6, Xz3et6, G24et6, P44et6,
 Y64et6, H94et6, Qb4et6, Zd4et6, Ig4et6, Ri4et6, Al4et6, Jn4et6,
 Sp4et6, Bs4et6, Ku4et6, Tw4et6, Cz4et6, L15et6, U35et6, D65et6,
 M85et6, Va5et6}, 1'b0} + {{1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, Ueo7v6}, 1'b1});
assign Nqh7z6 = Gfxm17[33:1];
assign Cixm17 = ({Vvh7z6, 1'b0} + {{Xd7et6, Ob7et6, F97et6, W67et6,
 N47et6, E27et6, Vz6et6, Mx6et6, Dv6et6, Us6et6, Lq6et6, Co6et6,
 Tl6et6, Kj6et6, Bh6et6, Se6et6, Jc6et6, Aa6et6, R76et6, I56et6,
 Z26et6, Q06et6, Hy5et6, Yv5et6, Pt5et6, Gr5et6, Xo5et6, Om5et6,
 Fk5et6, Wh5et6, Nf5et6, Ed5et6}, 1'b1});
assign {Ca3et6, Lc3et6, Ue3et6, Dh3et6, Mj3et6, Vl3et6, Eo3et6, Nq3et6,
 Ws3et6, Fv3et6, Ox3et6, Xz3et6, G24et6, P44et6, Y64et6, H94et6,
 Qb4et6, Zd4et6, Ig4et6, Ri4et6, Al4et6, Jn4et6, Sp4et6, Bs4et6,
 Ku4et6, Tw4et6, Cz4et6, L15et6, U35et6, D65et6, M85et6, Va5et6}
 = Cixm17[33:1];
assign Wkxm17 = ({{Nbaet6, Wdaet6, Fgaet6, Oiaet6, Xkaet6, Gnaet6,
 Ppaet6, Yraet6, Huaet6, Qwaet6}, 1'b0} + {{1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, Cfa7z6}, 1'b1});
assign P9i7z6 = Wkxm17[33:1];
assign Snxm17 = ({{1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 Fci7z6}, 1'b0} + {{Cfa7z6, Cfa7z6, Kfbet6, Bdbet6, Sabet6,
 J8bet6, A6bet6, R3bet6, I1bet6, Zyaet6}, 1'b1});
assign {Nbaet6, Wdaet6, Fgaet6, Oiaet6, Xkaet6, Gnaet6, Ppaet6, Yraet6,
 Huaet6, Qwaet6} = Snxm17[33:1];
assign Mqxm17 = ((Pcg7z6 - {A4xdt6, A4xdt6, A4xdt6, Alf7z6[31:3]}) -
 1'b0);
assign {Epmdt6, Dsmdt6, Cvmdt6, Bymdt6, A1ndt6, Z3ndt6, Y6ndt6, X9ndt6,
 Wcndt6, Vfndt6, Uindt6, Tlndt6, Sondt6, Rrndt6, Qundt6, Pxndt6,
 O0odt6, N3odt6, M6odt6, L9odt6, Kcodt6, Jfodt6, Iiodt6, Hlodt6,
 Goodt6, Frodt6, Euodt6, Dxodt6, C0pdt6, A3pdt6, Y5pdt6, W8pdt6}
 = Mqxm17[31:0];
assign Wtxm17 = ({Pcg7z6, 1'b0} + {{A4xdt6, A4xdt6, A4xdt6,
 Alf7z6[31:3]}, 1'b1});
assign {Ubpdt6, Sepdt6, Qhpdt6, Okpdt6, Mnpdt6, Kqpdt6, Itpdt6, Gwpdt6,
 Ezpdt6, C2qdt6, A5qdt6, Y7qdt6, Waqdt6, Udqdt6, Sgqdt6, Qjqdt6,
 Omqdt6, Mpqdt6, Ksqdt6, Ivqdt6, Gyqdt6, E1rdt6, C4rdt6, A7rdt6,
 Y9rdt6, Wcrdt6, Ufrdt6, Sirdt6, Qlrdt6, Oordt6, Mrrdt6, Kurdt6}
 = Wtxm17[33:1];
assign Gxxm17 = ((Zfg7z6 - {A4xdt6, A4xdt6, Alf7z6[31:2]}) - 1'b0);
assign {Ixrdt6, G0sdt6, E3sdt6, C6sdt6, A9sdt6, Ybsdt6, Wesdt6, Uhsdt6,
 Sksdt6, Qnsdt6, Oqsdt6, Mtsdt6, Kwsdt6, Izsdt6, G2tdt6, E5tdt6,
 C8tdt6, Abtdt6, Ydtdt6, Wgtdt6, Ujtdt6, Smtdt6, Qptdt6, Ostdt6,
 Mvtdt6, Kytdt6, I1udt6, G4udt6, E7udt6, Caudt6, Adudt6, Yfudt6}
 = Gxxm17[31:0];
assign Q0ym17 = ({Zfg7z6, 1'b0} + {{A4xdt6, A4xdt6, Alf7z6[31:2]}, 1'b1}
 );
assign {Wiudt6, Uludt6, Soudt6, Qrudt6, Ouudt6, Mxudt6, K0vdt6, I3vdt6,
 G6vdt6, E9vdt6, Ccvdt6, Afvdt6, Yhvdt6, Wkvdt6, Unvdt6, Sqvdt6,
 Qtvdt6, Owvdt6, Mzvdt6, K2wdt6, I5wdt6, G8wdt6, Ebwdt6, Bewdt6,
 Ygwdt6, Vjwdt6, Smwdt6, Ppwdt6, Mswdt6, Jvwdt6, Gywdt6, D1xdt6}
 = Q0ym17[33:1];
assign A4ym17 = ({{Tmg7z6, 1'b1}, 1'b0} + {{Jjg7z6, Wvl8v6}, 1'b1});
assign {Zfg7z6, Rma7z6} = A4ym17[33:1];
assign K7ym17 = ({{Onf7z6, 1'b1}, 1'b0} + {{Dqg7z6, Geo7v6}, 1'b1});
assign {Tmg7z6, Ona7z6} = K7ym17[33:1];
assign Iphdt6 = ((Kif7z6 == {Uff7z6, Arkdt6}) ? 1'b1 : 1'b0);
assign Uaym17 = ({{Vrhdt6, Zthdt6, Dwhdt6, Hyhdt6, L0idt6, P2idt6,
 T4idt6, X6idt6, B9idt6, Fbidt6, Jdidt6, Nfidt6, Rhidt6, Vjidt6,
 Zlidt6, Doidt6}, 1'b0} + {{1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, Hqidt6},
 1'b1});
assign Cqf7z6 = Uaym17[33:1];
assign Ldym17 = ({Ivf7z6, 1'b0} + {Ssf7z6, 1'b1});
assign {Vrhdt6, Zthdt6, Dwhdt6, Hyhdt6, L0idt6, P2idt6, T4idt6, X6idt6,
 B9idt6, Fbidt6, Jdidt6, Nfidt6, Rhidt6, Vjidt6, Zlidt6, Doidt6}
 = Ldym17[33:1];
assign Agym17 = ({{Xsidt6, Bvidt6, Fxidt6, Jzidt6, N1jdt6, R3jdt6,
 V5jdt6, Z7jdt6, Dajdt6, Gcjdt6, Jejdt6, Mgjdt6, Pijdt6, Skjdt6,
 Vmjdt6, Yojdt6, Brjdt6, Etjdt6, Hvjdt6, Kxjdt6, Nzjdt6, Q1kdt6,
 T3kdt6, W5kdt6, Z7kdt6, Cakdt6, Fckdt6, Iekdt6, Lgkdt6, Oikdt6,
 Rkkdt6, Umkdt6, Xokdt6}, 1'b0} + {{1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, Arkdt6}, 1'b1});
assign L0g7z6 = Agym17[33:1];
assign Riym17 = ({{1'b0, J5g7z6}, 1'b0} + {{1'b0, X2g7z6}, 1'b1});
assign {Xsidt6, Bvidt6, Fxidt6, Jzidt6, N1jdt6, R3jdt6, V5jdt6, Z7jdt6,
 Dajdt6, Gcjdt6, Jejdt6, Mgjdt6, Pijdt6, Skjdt6, Vmjdt6, Yojdt6,
 Brjdt6, Etjdt6, Hvjdt6, Kxjdt6, Nzjdt6, Q1kdt6, T3kdt6, W5kdt6,
 Z7kdt6, Cakdt6, Fckdt6, Iekdt6, Lgkdt6, Oikdt6, Rkkdt6, Umkdt6,
 Xokdt6} = Riym17[33:1];
assign Glym17 = (Fag7z6 * V7g7z6);
assign {Loa7z6, Ipa7z6, Fqa7z6, Cra7z6, Zra7z6, Xsa7z6, Vta7z6, Tua7z6,
 Rva7z6, Pwa7z6, Nxa7z6, Lya7z6, Jza7z6, H0b7z6, F1b7z6, D2b7z6,
 B3b7z6, Z3b7z6, X4b7z6, V5b7z6, T6b7z6, R7b7z6, P8b7z6, N9b7z6,
 Lab7z6, Jbb7z6, Hcb7z6, Fdb7z6, Deb7z6, Bfb7z6, Zfb7z6, Xgb7z6,
 Mtkdt6, Pvkdt6, Sxkdt6, Vzkdt6, Y1ldt6, B4ldt6, E6ldt6, H8ldt6,
 Kaldt6, Ncldt6, Qeldt6, Tgldt6, Wildt6, Zkldt6, Cnldt6, Fpldt6,
 Irldt6, Ltldt6, Ovldt6, Rxldt6, Uzldt6, X1mdt6, A4mdt6, D6mdt6,
 G8mdt6, Jamdt6, Mcmdt6, Pemdt6, Sgmdt6, Vimdt6, Ykmdt6, Bnmdt6}
 = Glym17[63:0];
assign Xnym17 = ((K2f7z6 - Rze7z6) - 1'b0);
assign {Fugdt6, Jwgdt6, Nygdt6, R0hdt6, V2hdt6, Z4hdt6} = Xnym17[5:0];
assign Mqym17 = ({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
 1'b1, 1'b1, 1'b1} << Jaf7z6);
assign Rje7z6 = Mqym17[31:0];
assign Etym17 = ({V1c7z6[31:27], 1'b0} + {V1c7z6[4:0], 1'b1});
assign {Oehdt6, Sghdt6, Wihdt6, Alhdt6, Enhdt6} = Etym17[33:1];
assign Uvym17 = (({1'b0, S0e7z6} - {1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 Yxd7z6}) - 1'b0);
assign Gvd7z6 = Uvym17[6:0];
assign Nlcdt6 = (({Dvc7z6[31:2], 1'b0, 1'b0} == {X0d7z6, 1'b0, 1'b0}) ?
 1'b1 : 1'b0);
assign Jyym17 = ({{Pdc7z6[31:2], 1'b0}, 1'b0} + {{1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0}, 1'b1});
assign {Xhd7z6, Vhb7z6} = Jyym17[33:1];
assign H1zm17 = ({vis_pc_o, 1'b0} + {{Vjc7z6[31], Vjc7z6[31],
 Vjc7z6[31], Vjc7z6[31], Vjc7z6[31], Vjc7z6[31], Vjc7z6[31],
 Vjc7z6[31], Vjc7z6[31], Vjc7z6[31], Vjc7z6[31], Vjc7z6[31],
 Vjc7z6[31], Vjc7z6[31], Vjc7z6[31], Vjc7z6[31], Vjc7z6[31],
 Vjc7z6[31], Vjc7z6[31], Vjc7z6[31], Vjc7z6[31], Vjc7z6[31],
 Vjc7z6[31], Vjc7z6[31], Vjc7z6[31], Vjc7z6[6:1]}, 1'b1});
assign Wkd7z6 = H1zm17[33:1];
assign F4zm17 = ({vis_pc_o, 1'b0} + {{Flc7z6[31], Flc7z6[31],
 Flc7z6[31], Flc7z6[31], Flc7z6[31], Flc7z6[31], Flc7z6[31],
 Flc7z6[31], Flc7z6[23:1]}, 1'b1});
assign Vnd7z6 = F4zm17[33:1];
assign D7zm17 = ({{L88et6, Ua8et6, Dd8et6, Mf8et6, Vh8et6, Ek8et6,
 Nm8et6, Wo8et6, Fr8et6, Ot8et6, Xv8et6, Gy8et6, P09et6, Y29et6,
 H59et6, Q79et6, Z99et6, Ic9et6, Re9et6, Ah9et6, Jj9et6, Sl9et6,
 Bo9et6, Kq9et6, Ts9et6, Cv9et6, Lx9et6, Uz9et6, D2aet6, M4aet6,
 V6aet6, E9aet6}, 1'b0} + {{1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, P58et6}, 1'b1});
assign {Cmm7z6[31:3], U28et6, Cmm7z6[1:0]} = D7zm17[33:1];
assign Z9zm17 = ({K1i7z6, 1'b0} + {Oyh7z6, 1'b1});
assign {L88et6, Ua8et6, Dd8et6, Mf8et6, Vh8et6, Ek8et6, Nm8et6, Wo8et6,
 Fr8et6, Ot8et6, Xv8et6, Gy8et6, P09et6, Y29et6, H59et6, Q79et6,
 Z99et6, Ic9et6, Re9et6, Ah9et6, Jj9et6, Sl9et6, Bo9et6, Kq9et6,
 Ts9et6, Cv9et6, Lx9et6, Uz9et6, D2aet6, M4aet6, V6aet6, E9aet6}
 = Z9zm17[33:1];
assign Tpt8v6 = (S7gdt6 & H9gdt6);
assign Ojt8v6 = (~(Q1fdt6 & Tpt8v6));
assign Aqt8v6 = (S7gdt6 & But8v6);
assign Hjt8v6 = (~(B0fdt6 & Aqt8v6));
assign Qkt8v6 = (Ojt8v6 & Hjt8v6);
assign Vqt8v6 = (~(But8v6 | S7gdt6));
assign Ckt8v6 = (~(Myedt6 & Vqt8v6));
assign Crt8v6 = (~(H9gdt6 | S7gdt6));
assign Vjt8v6 = (~(Xwedt6 & Crt8v6));
assign Jkt8v6 = (Ckt8v6 & Vjt8v6);
assign Xkt8v6 = (~(Qkt8v6 & Jkt8v6));
assign Int8v6 = (~(D6gdt6 & Xkt8v6));
assign Llt8v6 = (~(Ivedt6 & Tpt8v6));
assign Elt8v6 = (~(Ttedt6 & Aqt8v6));
assign Nmt8v6 = (Llt8v6 & Elt8v6);
assign Zlt8v6 = (~(Esedt6 & Vqt8v6));
assign Slt8v6 = (~(Pqedt6 & Crt8v6));
assign Gmt8v6 = (Zlt8v6 & Slt8v6);
assign Umt8v6 = (~(Nmt8v6 & Gmt8v6));
assign Bnt8v6 = (~(Umt8v6 & Iut8v6));
assign Pnt8v6 = (~(Int8v6 & Bnt8v6));
assign Utt8v6 = (~(O4gdt6 & Pnt8v6));
assign Dot8v6 = (~(Apedt6 & Tpt8v6));
assign Wnt8v6 = (~(Lnedt6 & Aqt8v6));
assign Fpt8v6 = (Dot8v6 & Wnt8v6);
assign Rot8v6 = (~(Wledt6 & Vqt8v6));
assign Kot8v6 = (~(Hkedt6 & Crt8v6));
assign Yot8v6 = (Rot8v6 & Kot8v6);
assign Mpt8v6 = (~(Fpt8v6 & Yot8v6));
assign Zst8v6 = (~(Mpt8v6 & D6gdt6));
assign Oqt8v6 = (~(Siedt6 & Tpt8v6));
assign Hqt8v6 = (~(Dhedt6 & Aqt8v6));
assign Est8v6 = (Oqt8v6 & Hqt8v6);
assign Qrt8v6 = (~(Ofedt6 & Vqt8v6));
assign Jrt8v6 = (~(Zdedt6 & Crt8v6));
assign Xrt8v6 = (Qrt8v6 & Jrt8v6);
assign Lst8v6 = (~(Est8v6 & Xrt8v6));
assign Sst8v6 = (~(Lst8v6 & Iut8v6));
assign Gtt8v6 = (Zst8v6 & Sst8v6);
assign Ntt8v6 = (Gtt8v6 | O4gdt6);
assign Acedt6 = (~(Utt8v6 & Ntt8v6));
assign But8v6 = (!H9gdt6);
assign Iut8v6 = (!D6gdt6);
assign B1u8v6 = (Aegdt6 & Pfgdt6);
assign Wut8v6 = (~(Wqfdt6 & B1u8v6));
assign I1u8v6 = (Aegdt6 & J5u8v6);
assign Put8v6 = (~(Hpfdt6 & I1u8v6));
assign Yvt8v6 = (Wut8v6 & Put8v6);
assign D2u8v6 = (~(J5u8v6 | Aegdt6));
assign Kvt8v6 = (~(Snfdt6 & D2u8v6));
assign K2u8v6 = (~(Pfgdt6 | Aegdt6));
assign Dvt8v6 = (~(Dmfdt6 & K2u8v6));
assign Rvt8v6 = (Kvt8v6 & Dvt8v6);
assign Fwt8v6 = (~(Yvt8v6 & Rvt8v6));
assign Qyt8v6 = (~(Lcgdt6 & Fwt8v6));
assign Twt8v6 = (~(Okfdt6 & B1u8v6));
assign Mwt8v6 = (~(Zifdt6 & I1u8v6));
assign Vxt8v6 = (Twt8v6 & Mwt8v6);
assign Hxt8v6 = (~(Khfdt6 & D2u8v6));
assign Axt8v6 = (~(Vffdt6 & K2u8v6));
assign Oxt8v6 = (Hxt8v6 & Axt8v6);
assign Cyt8v6 = (~(Vxt8v6 & Oxt8v6));
assign Jyt8v6 = (~(Cyt8v6 & Q5u8v6));
assign Xyt8v6 = (~(Qyt8v6 & Jyt8v6));
assign C5u8v6 = (~(Wagdt6 & Xyt8v6));
assign Lzt8v6 = (~(Gefdt6 & B1u8v6));
assign Ezt8v6 = (~(Rcfdt6 & I1u8v6));
assign N0u8v6 = (Lzt8v6 & Ezt8v6);
assign Zzt8v6 = (~(Cbfdt6 & D2u8v6));
assign Szt8v6 = (~(N9fdt6 & K2u8v6));
assign G0u8v6 = (Zzt8v6 & Szt8v6);
assign U0u8v6 = (~(N0u8v6 & G0u8v6));
assign H4u8v6 = (~(U0u8v6 & Lcgdt6));
assign W1u8v6 = (~(Y7fdt6 & B1u8v6));
assign P1u8v6 = (~(J6fdt6 & I1u8v6));
assign M3u8v6 = (W1u8v6 & P1u8v6);
assign Y2u8v6 = (~(U4fdt6 & D2u8v6));
assign R2u8v6 = (~(F3fdt6 & K2u8v6));
assign F3u8v6 = (Y2u8v6 & R2u8v6);
assign T3u8v6 = (~(M3u8v6 & F3u8v6));
assign A4u8v6 = (~(T3u8v6 & Q5u8v6));
assign O4u8v6 = (H4u8v6 & A4u8v6);
assign V4u8v6 = (O4u8v6 | Wagdt6);
assign B8cdt6 = (~(C5u8v6 & V4u8v6));
assign J5u8v6 = (!Pfgdt6);
assign Q5u8v6 = (!Lcgdt6);
assign Imu8v6 = (Alhdt6 & Enhdt6);
assign E6u8v6 = (~(Neo7v6 & Imu8v6));
assign Pmu8v6 = (Alhdt6 & Lru8v6);
assign X5u8v6 = (~(Cve7z6[30] & Pmu8v6));
assign G7u8v6 = (E6u8v6 & X5u8v6);
assign Knu8v6 = (~(Lru8v6 | Alhdt6));
assign S6u8v6 = (~(Cve7z6[29] & Knu8v6));
assign Rnu8v6 = (~(Enhdt6 | Alhdt6));
assign L6u8v6 = (~(Cve7z6[28] & Rnu8v6));
assign Z6u8v6 = (S6u8v6 & L6u8v6);
assign N7u8v6 = (~(G7u8v6 & Z6u8v6));
assign Y9u8v6 = (~(Wihdt6 & N7u8v6));
assign B8u8v6 = (~(Cve7z6[27] & Imu8v6));
assign U7u8v6 = (~(Cve7z6[26] & Pmu8v6));
assign D9u8v6 = (B8u8v6 & U7u8v6);
assign P8u8v6 = (~(Cve7z6[25] & Knu8v6));
assign I8u8v6 = (~(Cve7z6[24] & Rnu8v6));
assign W8u8v6 = (P8u8v6 & I8u8v6);
assign K9u8v6 = (~(D9u8v6 & W8u8v6));
assign R9u8v6 = (~(K9u8v6 & Sru8v6));
assign Fau8v6 = (~(Y9u8v6 & R9u8v6));
assign Ifu8v6 = (~(Sghdt6 & Fau8v6));
assign Tau8v6 = (~(Cve7z6[23] & Imu8v6));
assign Mau8v6 = (~(Cve7z6[22] & Pmu8v6));
assign Vbu8v6 = (Tau8v6 & Mau8v6);
assign Hbu8v6 = (~(Cve7z6[21] & Knu8v6));
assign Abu8v6 = (~(Cve7z6[20] & Rnu8v6));
assign Obu8v6 = (Hbu8v6 & Abu8v6);
assign Ccu8v6 = (~(Vbu8v6 & Obu8v6));
assign Neu8v6 = (~(Ccu8v6 & Wihdt6));
assign Qcu8v6 = (~(Cve7z6[19] & Imu8v6));
assign Jcu8v6 = (~(Cve7z6[18] & Pmu8v6));
assign Sdu8v6 = (Qcu8v6 & Jcu8v6);
assign Edu8v6 = (~(Cve7z6[17] & Knu8v6));
assign Xcu8v6 = (~(Cve7z6[16] & Rnu8v6));
assign Ldu8v6 = (Edu8v6 & Xcu8v6);
assign Zdu8v6 = (~(Sdu8v6 & Ldu8v6));
assign Geu8v6 = (~(Zdu8v6 & Sru8v6));
assign Ueu8v6 = (~(Neu8v6 & Geu8v6));
assign Bfu8v6 = (~(Ueu8v6 & Zru8v6));
assign Pfu8v6 = (~(Ifu8v6 & Bfu8v6));
assign Eru8v6 = (~(Oehdt6 & Pfu8v6));
assign Dgu8v6 = (~(Cve7z6[15] & Imu8v6));
assign Wfu8v6 = (~(Cve7z6[14] & Pmu8v6));
assign Fhu8v6 = (Dgu8v6 & Wfu8v6);
assign Rgu8v6 = (~(Cve7z6[13] & Knu8v6));
assign Kgu8v6 = (~(Cve7z6[12] & Rnu8v6));
assign Ygu8v6 = (Rgu8v6 & Kgu8v6);
assign Mhu8v6 = (~(Fhu8v6 & Ygu8v6));
assign Xju8v6 = (~(Mhu8v6 & Wihdt6));
assign Aiu8v6 = (~(Cve7z6[11] & Imu8v6));
assign Thu8v6 = (~(Cve7z6[10] & Pmu8v6));
assign Cju8v6 = (Aiu8v6 & Thu8v6);
assign Oiu8v6 = (~(Cve7z6[9] & Knu8v6));
assign Hiu8v6 = (~(Cve7z6[8] & Rnu8v6));
assign Viu8v6 = (Oiu8v6 & Hiu8v6);
assign Jju8v6 = (~(Cju8v6 & Viu8v6));
assign Qju8v6 = (~(Jju8v6 & Sru8v6));
assign Eku8v6 = (~(Xju8v6 & Qju8v6));
assign Jqu8v6 = (~(Eku8v6 & Sghdt6));
assign Sku8v6 = (~(Cve7z6[7] & Imu8v6));
assign Lku8v6 = (~(Cve7z6[6] & Pmu8v6));
assign Ulu8v6 = (Sku8v6 & Lku8v6);
assign Glu8v6 = (~(Cve7z6[5] & Knu8v6));
assign Zku8v6 = (~(Cve7z6[4] & Rnu8v6));
assign Nlu8v6 = (Glu8v6 & Zku8v6);
assign Bmu8v6 = (~(Ulu8v6 & Nlu8v6));
assign Opu8v6 = (~(Bmu8v6 & Wihdt6));
assign Dnu8v6 = (~(Cve7z6[3] & Imu8v6));
assign Wmu8v6 = (~(Cve7z6[2] & Pmu8v6));
assign Tou8v6 = (Dnu8v6 & Wmu8v6);
assign Fou8v6 = (~(Cve7z6[1] & Knu8v6));
assign Ynu8v6 = (~(Cve7z6[0] & Rnu8v6));
assign Mou8v6 = (Fou8v6 & Ynu8v6);
assign Apu8v6 = (~(Tou8v6 & Mou8v6));
assign Hpu8v6 = (~(Apu8v6 & Sru8v6));
assign Vpu8v6 = (~(Opu8v6 & Hpu8v6));
assign Cqu8v6 = (~(Vpu8v6 & Zru8v6));
assign Qqu8v6 = (Jqu8v6 & Cqu8v6);
assign Xqu8v6 = (Qqu8v6 | Oehdt6);
assign Q9hdt6 = (~(Eru8v6 & Xqu8v6));
assign Lru8v6 = (!Enhdt6);
assign Sru8v6 = (!Wihdt6);
assign Zru8v6 = (!Sghdt6);
assign Nsu8v6 = (~(H8k7z6[7] & Pehet6));
assign Gsu8v6 = (~(H8k7z6[6] & Qxu8v6));
assign Usu8v6 = (~(Nsu8v6 & Gsu8v6));
assign Duu8v6 = (~(Cbhet6 & Usu8v6));
assign Itu8v6 = (~(H8k7z6[5] & Pehet6));
assign Btu8v6 = (~(H8k7z6[4] & Qxu8v6));
assign Ptu8v6 = (~(Itu8v6 & Btu8v6));
assign Wtu8v6 = (~(Ptu8v6 & Xxu8v6));
assign Kuu8v6 = (~(Duu8v6 & Wtu8v6));
assign Jxu8v6 = (~(P7het6 & Kuu8v6));
assign Yuu8v6 = (~(H8k7z6[3] & Pehet6));
assign Ruu8v6 = (~(H8k7z6[2] & Qxu8v6));
assign Fvu8v6 = (~(Yuu8v6 & Ruu8v6));
assign Owu8v6 = (~(Fvu8v6 & Cbhet6));
assign Tvu8v6 = (~(H8k7z6[1] & Pehet6));
assign Mvu8v6 = (~(H8k7z6[0] & Qxu8v6));
assign Awu8v6 = (~(Tvu8v6 & Mvu8v6));
assign Hwu8v6 = (~(Awu8v6 & Xxu8v6));
assign Vwu8v6 = (~(Owu8v6 & Hwu8v6));
assign Cxu8v6 = (Eyu8v6 | P7het6);
assign C4het6 = (~(Jxu8v6 & Cxu8v6));
assign Qxu8v6 = (!Pehet6);
assign Xxu8v6 = (!Cbhet6);
assign Eyu8v6 = (!Vwu8v6);
assign Syu8v6 = (~(H8k7z6[7] & Pshet6));
assign Lyu8v6 = (~(H8k7z6[6] & C4v8v6));
assign Zyu8v6 = (~(Syu8v6 & Lyu8v6));
assign I0v8v6 = (~(Cphet6 & Zyu8v6));
assign Nzu8v6 = (~(H8k7z6[5] & Pshet6));
assign Gzu8v6 = (~(H8k7z6[4] & C4v8v6));
assign Uzu8v6 = (~(Nzu8v6 & Gzu8v6));
assign B0v8v6 = (~(Uzu8v6 & V3v8v6));
assign P0v8v6 = (~(I0v8v6 & B0v8v6));
assign O3v8v6 = (~(Plhet6 & P0v8v6));
assign D1v8v6 = (~(H8k7z6[3] & Pshet6));
assign W0v8v6 = (~(H8k7z6[2] & C4v8v6));
assign K1v8v6 = (~(D1v8v6 & W0v8v6));
assign T2v8v6 = (~(K1v8v6 & Cphet6));
assign Y1v8v6 = (~(H8k7z6[1] & Pshet6));
assign R1v8v6 = (~(H8k7z6[0] & C4v8v6));
assign F2v8v6 = (~(Y1v8v6 & R1v8v6));
assign M2v8v6 = (~(F2v8v6 & V3v8v6));
assign A3v8v6 = (~(T2v8v6 & M2v8v6));
assign H3v8v6 = (J4v8v6 | Plhet6);
assign Cihet6 = (~(O3v8v6 & H3v8v6));
assign V3v8v6 = (!Cphet6);
assign C4v8v6 = (!Pshet6);
assign J4v8v6 = (!A3v8v6);
assign X4v8v6 = (~(Pik7z6[7] & P6iet6));
assign Q4v8v6 = (~(Pik7z6[6] & Aav8v6));
assign E5v8v6 = (~(X4v8v6 & Q4v8v6));
assign N6v8v6 = (~(C3iet6 & E5v8v6));
assign S5v8v6 = (~(Pik7z6[5] & P6iet6));
assign L5v8v6 = (~(Pik7z6[4] & Aav8v6));
assign Z5v8v6 = (~(S5v8v6 & L5v8v6));
assign G6v8v6 = (~(Z5v8v6 & Hav8v6));
assign U6v8v6 = (~(N6v8v6 & G6v8v6));
assign T9v8v6 = (~(Pzhet6 & U6v8v6));
assign I7v8v6 = (~(Pik7z6[3] & P6iet6));
assign B7v8v6 = (~(Pik7z6[2] & Aav8v6));
assign P7v8v6 = (~(I7v8v6 & B7v8v6));
assign Y8v8v6 = (~(P7v8v6 & C3iet6));
assign D8v8v6 = (~(Pik7z6[1] & P6iet6));
assign W7v8v6 = (~(Pik7z6[0] & Aav8v6));
assign K8v8v6 = (~(D8v8v6 & W7v8v6));
assign R8v8v6 = (~(K8v8v6 & Hav8v6));
assign F9v8v6 = (~(Y8v8v6 & R8v8v6));
assign M9v8v6 = (Oav8v6 | Pzhet6);
assign Cwhet6 = (~(T9v8v6 & M9v8v6));
assign Aav8v6 = (!P6iet6);
assign Hav8v6 = (!C3iet6);
assign Oav8v6 = (!F9v8v6);
assign Cbv8v6 = (~(Pik7z6[7] & Pkiet6));
assign Vav8v6 = (~(Pik7z6[6] & Mgv8v6));
assign Jbv8v6 = (~(Cbv8v6 & Vav8v6));
assign Scv8v6 = (~(Chiet6 & Jbv8v6));
assign Xbv8v6 = (~(Pik7z6[5] & Pkiet6));
assign Qbv8v6 = (~(Pik7z6[4] & Mgv8v6));
assign Ecv8v6 = (~(Xbv8v6 & Qbv8v6));
assign Lcv8v6 = (~(Ecv8v6 & Fgv8v6));
assign Zcv8v6 = (~(Scv8v6 & Lcv8v6));
assign Yfv8v6 = (~(Pdiet6 & Zcv8v6));
assign Ndv8v6 = (~(Pik7z6[3] & Pkiet6));
assign Gdv8v6 = (~(Pik7z6[2] & Mgv8v6));
assign Udv8v6 = (~(Ndv8v6 & Gdv8v6));
assign Dfv8v6 = (~(Udv8v6 & Chiet6));
assign Iev8v6 = (~(Pik7z6[1] & Pkiet6));
assign Bev8v6 = (~(Pik7z6[0] & Mgv8v6));
assign Pev8v6 = (~(Iev8v6 & Bev8v6));
assign Wev8v6 = (~(Pev8v6 & Fgv8v6));
assign Kfv8v6 = (~(Dfv8v6 & Wev8v6));
assign Rfv8v6 = (Tgv8v6 | Pdiet6);
assign Caiet6 = (~(Yfv8v6 & Rfv8v6));
assign Fgv8v6 = (!Chiet6);
assign Mgv8v6 = (!Pkiet6);
assign Tgv8v6 = (!Kfv8v6);
assign Hhv8v6 = (~(Xsk7z6[7] & Pyiet6));
assign Ahv8v6 = (~(Xsk7z6[6] & Kmv8v6));
assign Ohv8v6 = (~(Hhv8v6 & Ahv8v6));
assign Xiv8v6 = (~(Cviet6 & Ohv8v6));
assign Civ8v6 = (~(Xsk7z6[5] & Pyiet6));
assign Vhv8v6 = (~(Xsk7z6[4] & Kmv8v6));
assign Jiv8v6 = (~(Civ8v6 & Vhv8v6));
assign Qiv8v6 = (~(Jiv8v6 & Rmv8v6));
assign Ejv8v6 = (~(Xiv8v6 & Qiv8v6));
assign Dmv8v6 = (~(Priet6 & Ejv8v6));
assign Sjv8v6 = (~(Xsk7z6[3] & Pyiet6));
assign Ljv8v6 = (~(Xsk7z6[2] & Kmv8v6));
assign Zjv8v6 = (~(Sjv8v6 & Ljv8v6));
assign Ilv8v6 = (~(Zjv8v6 & Cviet6));
assign Nkv8v6 = (~(Xsk7z6[1] & Pyiet6));
assign Gkv8v6 = (~(Xsk7z6[0] & Kmv8v6));
assign Ukv8v6 = (~(Nkv8v6 & Gkv8v6));
assign Blv8v6 = (~(Ukv8v6 & Rmv8v6));
assign Plv8v6 = (~(Ilv8v6 & Blv8v6));
assign Wlv8v6 = (Ymv8v6 | Priet6);
assign Coiet6 = (~(Dmv8v6 & Wlv8v6));
assign Kmv8v6 = (!Pyiet6);
assign Rmv8v6 = (!Cviet6);
assign Ymv8v6 = (!Plv8v6);
assign Mnv8v6 = (~(Xsk7z6[7] & Pcjet6));
assign Fnv8v6 = (~(Xsk7z6[6] & Wsv8v6));
assign Tnv8v6 = (~(Mnv8v6 & Fnv8v6));
assign Cpv8v6 = (~(C9jet6 & Tnv8v6));
assign Hov8v6 = (~(Xsk7z6[5] & Pcjet6));
assign Aov8v6 = (~(Xsk7z6[4] & Wsv8v6));
assign Oov8v6 = (~(Hov8v6 & Aov8v6));
assign Vov8v6 = (~(Oov8v6 & Psv8v6));
assign Jpv8v6 = (~(Cpv8v6 & Vov8v6));
assign Isv8v6 = (~(P5jet6 & Jpv8v6));
assign Xpv8v6 = (~(Xsk7z6[3] & Pcjet6));
assign Qpv8v6 = (~(Xsk7z6[2] & Wsv8v6));
assign Eqv8v6 = (~(Xpv8v6 & Qpv8v6));
assign Nrv8v6 = (~(Eqv8v6 & C9jet6));
assign Sqv8v6 = (~(Xsk7z6[1] & Pcjet6));
assign Lqv8v6 = (~(Xsk7z6[0] & Wsv8v6));
assign Zqv8v6 = (~(Sqv8v6 & Lqv8v6));
assign Grv8v6 = (~(Zqv8v6 & Psv8v6));
assign Urv8v6 = (~(Nrv8v6 & Grv8v6));
assign Bsv8v6 = (Dtv8v6 | P5jet6);
assign C2jet6 = (~(Isv8v6 & Bsv8v6));
assign Psv8v6 = (!C9jet6);
assign Wsv8v6 = (!Pcjet6);
assign Dtv8v6 = (!Urv8v6);
assign Rtv8v6 = (~(F3l7z6[7] & Pqjet6));
assign Ktv8v6 = (~(F3l7z6[6] & Uyv8v6));
assign Ytv8v6 = (~(Rtv8v6 & Ktv8v6));
assign Hvv8v6 = (~(Cnjet6 & Ytv8v6));
assign Muv8v6 = (~(F3l7z6[5] & Pqjet6));
assign Fuv8v6 = (~(F3l7z6[4] & Uyv8v6));
assign Tuv8v6 = (~(Muv8v6 & Fuv8v6));
assign Avv8v6 = (~(Tuv8v6 & Bzv8v6));
assign Ovv8v6 = (~(Hvv8v6 & Avv8v6));
assign Nyv8v6 = (~(Pjjet6 & Ovv8v6));
assign Cwv8v6 = (~(F3l7z6[3] & Pqjet6));
assign Vvv8v6 = (~(F3l7z6[2] & Uyv8v6));
assign Jwv8v6 = (~(Cwv8v6 & Vvv8v6));
assign Sxv8v6 = (~(Jwv8v6 & Cnjet6));
assign Xwv8v6 = (~(F3l7z6[1] & Pqjet6));
assign Qwv8v6 = (~(F3l7z6[0] & Uyv8v6));
assign Exv8v6 = (~(Xwv8v6 & Qwv8v6));
assign Lxv8v6 = (~(Exv8v6 & Bzv8v6));
assign Zxv8v6 = (~(Sxv8v6 & Lxv8v6));
assign Gyv8v6 = (Izv8v6 | Pjjet6);
assign Cgjet6 = (~(Nyv8v6 & Gyv8v6));
assign Uyv8v6 = (!Pqjet6);
assign Bzv8v6 = (!Cnjet6);
assign Izv8v6 = (!Zxv8v6);
assign Wzv8v6 = (~(F3l7z6[7] & P4ket6));
assign Pzv8v6 = (~(F3l7z6[6] & G5w8v6));
assign D0w8v6 = (~(Wzv8v6 & Pzv8v6));
assign M1w8v6 = (~(C1ket6 & D0w8v6));
assign R0w8v6 = (~(F3l7z6[5] & P4ket6));
assign K0w8v6 = (~(F3l7z6[4] & G5w8v6));
assign Y0w8v6 = (~(R0w8v6 & K0w8v6));
assign F1w8v6 = (~(Y0w8v6 & Z4w8v6));
assign T1w8v6 = (~(M1w8v6 & F1w8v6));
assign S4w8v6 = (~(Pxjet6 & T1w8v6));
assign H2w8v6 = (~(F3l7z6[3] & P4ket6));
assign A2w8v6 = (~(F3l7z6[2] & G5w8v6));
assign O2w8v6 = (~(H2w8v6 & A2w8v6));
assign X3w8v6 = (~(O2w8v6 & C1ket6));
assign C3w8v6 = (~(F3l7z6[1] & P4ket6));
assign V2w8v6 = (~(F3l7z6[0] & G5w8v6));
assign J3w8v6 = (~(C3w8v6 & V2w8v6));
assign Q3w8v6 = (~(J3w8v6 & Z4w8v6));
assign E4w8v6 = (~(X3w8v6 & Q3w8v6));
assign L4w8v6 = (N5w8v6 | Pxjet6);
assign Cujet6 = (~(S4w8v6 & L4w8v6));
assign Z4w8v6 = (!C1ket6);
assign G5w8v6 = (!P4ket6);
assign N5w8v6 = (!E4w8v6);
assign B6w8v6 = (~(Ndl7z6[7] & Piket6));
assign U5w8v6 = (~(Ndl7z6[6] & Ebw8v6));
assign I6w8v6 = (~(B6w8v6 & U5w8v6));
assign R7w8v6 = (~(Cfket6 & I6w8v6));
assign W6w8v6 = (~(Ndl7z6[5] & Piket6));
assign P6w8v6 = (~(Ndl7z6[4] & Ebw8v6));
assign D7w8v6 = (~(W6w8v6 & P6w8v6));
assign K7w8v6 = (~(D7w8v6 & Lbw8v6));
assign Y7w8v6 = (~(R7w8v6 & K7w8v6));
assign Xaw8v6 = (~(Pbket6 & Y7w8v6));
assign M8w8v6 = (~(Ndl7z6[3] & Piket6));
assign F8w8v6 = (~(Ndl7z6[2] & Ebw8v6));
assign T8w8v6 = (~(M8w8v6 & F8w8v6));
assign Caw8v6 = (~(T8w8v6 & Cfket6));
assign H9w8v6 = (~(Ndl7z6[1] & Piket6));
assign A9w8v6 = (~(Ndl7z6[0] & Ebw8v6));
assign O9w8v6 = (~(H9w8v6 & A9w8v6));
assign V9w8v6 = (~(O9w8v6 & Lbw8v6));
assign Jaw8v6 = (~(Caw8v6 & V9w8v6));
assign Qaw8v6 = (Sbw8v6 | Pbket6);
assign C8ket6 = (~(Xaw8v6 & Qaw8v6));
assign Ebw8v6 = (!Piket6);
assign Lbw8v6 = (!Cfket6);
assign Sbw8v6 = (!Jaw8v6);
assign Gcw8v6 = (~(Ndl7z6[7] & Pwket6));
assign Zbw8v6 = (~(Ndl7z6[6] & Qhw8v6));
assign Ncw8v6 = (~(Gcw8v6 & Zbw8v6));
assign Wdw8v6 = (~(Ctket6 & Ncw8v6));
assign Bdw8v6 = (~(Ndl7z6[5] & Pwket6));
assign Ucw8v6 = (~(Ndl7z6[4] & Qhw8v6));
assign Idw8v6 = (~(Bdw8v6 & Ucw8v6));
assign Pdw8v6 = (~(Idw8v6 & Jhw8v6));
assign Dew8v6 = (~(Wdw8v6 & Pdw8v6));
assign Chw8v6 = (~(Ppket6 & Dew8v6));
assign Rew8v6 = (~(Ndl7z6[3] & Pwket6));
assign Kew8v6 = (~(Ndl7z6[2] & Qhw8v6));
assign Yew8v6 = (~(Rew8v6 & Kew8v6));
assign Hgw8v6 = (~(Yew8v6 & Ctket6));
assign Mfw8v6 = (~(Ndl7z6[1] & Pwket6));
assign Ffw8v6 = (~(Ndl7z6[0] & Qhw8v6));
assign Tfw8v6 = (~(Mfw8v6 & Ffw8v6));
assign Agw8v6 = (~(Tfw8v6 & Jhw8v6));
assign Ogw8v6 = (~(Hgw8v6 & Agw8v6));
assign Vgw8v6 = (Xhw8v6 | Ppket6);
assign Cmket6 = (~(Chw8v6 & Vgw8v6));
assign Jhw8v6 = (!Ctket6);
assign Qhw8v6 = (!Pwket6);
assign Xhw8v6 = (!Ogw8v6);
assign Liw8v6 = (~(Vnl7z6[7] & Palet6));
assign Eiw8v6 = (~(Vnl7z6[6] & Onw8v6));
assign Siw8v6 = (~(Liw8v6 & Eiw8v6));
assign Bkw8v6 = (~(C7let6 & Siw8v6));
assign Gjw8v6 = (~(Vnl7z6[5] & Palet6));
assign Ziw8v6 = (~(Vnl7z6[4] & Onw8v6));
assign Njw8v6 = (~(Gjw8v6 & Ziw8v6));
assign Ujw8v6 = (~(Njw8v6 & Vnw8v6));
assign Ikw8v6 = (~(Bkw8v6 & Ujw8v6));
assign Hnw8v6 = (~(P3let6 & Ikw8v6));
assign Wkw8v6 = (~(Vnl7z6[3] & Palet6));
assign Pkw8v6 = (~(Vnl7z6[2] & Onw8v6));
assign Dlw8v6 = (~(Wkw8v6 & Pkw8v6));
assign Mmw8v6 = (~(Dlw8v6 & C7let6));
assign Rlw8v6 = (~(Vnl7z6[1] & Palet6));
assign Klw8v6 = (~(Vnl7z6[0] & Onw8v6));
assign Ylw8v6 = (~(Rlw8v6 & Klw8v6));
assign Fmw8v6 = (~(Ylw8v6 & Vnw8v6));
assign Tmw8v6 = (~(Mmw8v6 & Fmw8v6));
assign Anw8v6 = (Cow8v6 | P3let6);
assign C0let6 = (~(Hnw8v6 & Anw8v6));
assign Onw8v6 = (!Palet6);
assign Vnw8v6 = (!C7let6);
assign Cow8v6 = (!Tmw8v6);
assign Qow8v6 = (~(Vnl7z6[7] & Polet6));
assign Jow8v6 = (~(Vnl7z6[6] & Auw8v6));
assign Xow8v6 = (~(Qow8v6 & Jow8v6));
assign Gqw8v6 = (~(Cllet6 & Xow8v6));
assign Lpw8v6 = (~(Vnl7z6[5] & Polet6));
assign Epw8v6 = (~(Vnl7z6[4] & Auw8v6));
assign Spw8v6 = (~(Lpw8v6 & Epw8v6));
assign Zpw8v6 = (~(Spw8v6 & Ttw8v6));
assign Nqw8v6 = (~(Gqw8v6 & Zpw8v6));
assign Mtw8v6 = (~(Phlet6 & Nqw8v6));
assign Brw8v6 = (~(Vnl7z6[3] & Polet6));
assign Uqw8v6 = (~(Vnl7z6[2] & Auw8v6));
assign Irw8v6 = (~(Brw8v6 & Uqw8v6));
assign Rsw8v6 = (~(Irw8v6 & Cllet6));
assign Wrw8v6 = (~(Vnl7z6[1] & Polet6));
assign Prw8v6 = (~(Vnl7z6[0] & Auw8v6));
assign Dsw8v6 = (~(Wrw8v6 & Prw8v6));
assign Ksw8v6 = (~(Dsw8v6 & Ttw8v6));
assign Ysw8v6 = (~(Rsw8v6 & Ksw8v6));
assign Ftw8v6 = (Huw8v6 | Phlet6);
assign Celet6 = (~(Mtw8v6 & Ftw8v6));
assign Ttw8v6 = (!Cllet6);
assign Auw8v6 = (!Polet6);
assign Huw8v6 = (!Ysw8v6);
assign Vuw8v6 = (~(Dyl7z6[7] & P2met6));
assign Ouw8v6 = (~(Dyl7z6[6] & Yzw8v6));
assign Cvw8v6 = (~(Vuw8v6 & Ouw8v6));
assign Lww8v6 = (~(Czlet6 & Cvw8v6));
assign Qvw8v6 = (~(Dyl7z6[5] & P2met6));
assign Jvw8v6 = (~(Dyl7z6[4] & Yzw8v6));
assign Xvw8v6 = (~(Qvw8v6 & Jvw8v6));
assign Eww8v6 = (~(Xvw8v6 & F0x8v6));
assign Sww8v6 = (~(Lww8v6 & Eww8v6));
assign Rzw8v6 = (~(Pvlet6 & Sww8v6));
assign Gxw8v6 = (~(Dyl7z6[3] & P2met6));
assign Zww8v6 = (~(Dyl7z6[2] & Yzw8v6));
assign Nxw8v6 = (~(Gxw8v6 & Zww8v6));
assign Wyw8v6 = (~(Nxw8v6 & Czlet6));
assign Byw8v6 = (~(Dyl7z6[1] & P2met6));
assign Uxw8v6 = (~(Dyl7z6[0] & Yzw8v6));
assign Iyw8v6 = (~(Byw8v6 & Uxw8v6));
assign Pyw8v6 = (~(Iyw8v6 & F0x8v6));
assign Dzw8v6 = (~(Wyw8v6 & Pyw8v6));
assign Kzw8v6 = (M0x8v6 | Pvlet6);
assign Cslet6 = (~(Rzw8v6 & Kzw8v6));
assign Yzw8v6 = (!P2met6);
assign F0x8v6 = (!Czlet6);
assign M0x8v6 = (!Dzw8v6);
assign A1x8v6 = (~(Dyl7z6[7] & Pgmet6));
assign T0x8v6 = (~(Dyl7z6[6] & K6x8v6));
assign H1x8v6 = (~(A1x8v6 & T0x8v6));
assign Q2x8v6 = (~(Cdmet6 & H1x8v6));
assign V1x8v6 = (~(Dyl7z6[5] & Pgmet6));
assign O1x8v6 = (~(Dyl7z6[4] & K6x8v6));
assign C2x8v6 = (~(V1x8v6 & O1x8v6));
assign J2x8v6 = (~(C2x8v6 & D6x8v6));
assign X2x8v6 = (~(Q2x8v6 & J2x8v6));
assign W5x8v6 = (~(P9met6 & X2x8v6));
assign L3x8v6 = (~(Dyl7z6[3] & Pgmet6));
assign E3x8v6 = (~(Dyl7z6[2] & K6x8v6));
assign S3x8v6 = (~(L3x8v6 & E3x8v6));
assign B5x8v6 = (~(S3x8v6 & Cdmet6));
assign G4x8v6 = (~(Dyl7z6[1] & Pgmet6));
assign Z3x8v6 = (~(Dyl7z6[0] & K6x8v6));
assign N4x8v6 = (~(G4x8v6 & Z3x8v6));
assign U4x8v6 = (~(N4x8v6 & D6x8v6));
assign I5x8v6 = (~(B5x8v6 & U4x8v6));
assign P5x8v6 = (R6x8v6 | P9met6);
assign C6met6 = (~(W5x8v6 & P5x8v6));
assign D6x8v6 = (!Cdmet6);
assign K6x8v6 = (!Pgmet6);
assign R6x8v6 = (!I5x8v6);
assign F7x8v6 = (~(L8m7z6[7] & Pumet6));
assign Y6x8v6 = (~(L8m7z6[6] & Icx8v6));
assign M7x8v6 = (~(F7x8v6 & Y6x8v6));
assign V8x8v6 = (~(Crmet6 & M7x8v6));
assign A8x8v6 = (~(L8m7z6[5] & Pumet6));
assign T7x8v6 = (~(L8m7z6[4] & Icx8v6));
assign H8x8v6 = (~(A8x8v6 & T7x8v6));
assign O8x8v6 = (~(H8x8v6 & Pcx8v6));
assign C9x8v6 = (~(V8x8v6 & O8x8v6));
assign Bcx8v6 = (~(Pnmet6 & C9x8v6));
assign Q9x8v6 = (~(L8m7z6[3] & Pumet6));
assign J9x8v6 = (~(L8m7z6[2] & Icx8v6));
assign X9x8v6 = (~(Q9x8v6 & J9x8v6));
assign Gbx8v6 = (~(X9x8v6 & Crmet6));
assign Lax8v6 = (~(L8m7z6[1] & Pumet6));
assign Eax8v6 = (~(L8m7z6[0] & Icx8v6));
assign Sax8v6 = (~(Lax8v6 & Eax8v6));
assign Zax8v6 = (~(Sax8v6 & Pcx8v6));
assign Nbx8v6 = (~(Gbx8v6 & Zax8v6));
assign Ubx8v6 = (Wcx8v6 | Pnmet6);
assign Ckmet6 = (~(Bcx8v6 & Ubx8v6));
assign Icx8v6 = (!Pumet6);
assign Pcx8v6 = (!Crmet6);
assign Wcx8v6 = (!Nbx8v6);
assign Kdx8v6 = (~(L8m7z6[7] & P8net6));
assign Ddx8v6 = (~(L8m7z6[6] & Uix8v6));
assign Rdx8v6 = (~(Kdx8v6 & Ddx8v6));
assign Afx8v6 = (~(C5net6 & Rdx8v6));
assign Fex8v6 = (~(L8m7z6[5] & P8net6));
assign Ydx8v6 = (~(L8m7z6[4] & Uix8v6));
assign Mex8v6 = (~(Fex8v6 & Ydx8v6));
assign Tex8v6 = (~(Mex8v6 & Nix8v6));
assign Hfx8v6 = (~(Afx8v6 & Tex8v6));
assign Gix8v6 = (~(P1net6 & Hfx8v6));
assign Vfx8v6 = (~(L8m7z6[3] & P8net6));
assign Ofx8v6 = (~(L8m7z6[2] & Uix8v6));
assign Cgx8v6 = (~(Vfx8v6 & Ofx8v6));
assign Lhx8v6 = (~(Cgx8v6 & C5net6));
assign Qgx8v6 = (~(L8m7z6[1] & P8net6));
assign Jgx8v6 = (~(L8m7z6[0] & Uix8v6));
assign Xgx8v6 = (~(Qgx8v6 & Jgx8v6));
assign Ehx8v6 = (~(Xgx8v6 & Nix8v6));
assign Shx8v6 = (~(Lhx8v6 & Ehx8v6));
assign Zhx8v6 = (Bjx8v6 | P1net6);
assign Cymet6 = (~(Gix8v6 & Zhx8v6));
assign Nix8v6 = (!C5net6);
assign Uix8v6 = (!P8net6);
assign Bjx8v6 = (!Shx8v6);
assign Tzx8v6 = (S0zet6 & T2zet6);
assign Pjx8v6 = (~(Vbo7v6 & Tzx8v6));
assign A0y8v6 = (S0zet6 & D5y8v6);
assign Ijx8v6 = (~(M6a7z6 & A0y8v6));
assign Rkx8v6 = (Pjx8v6 & Ijx8v6);
assign V0y8v6 = (~(D5y8v6 | S0zet6));
assign Dkx8v6 = (~(U6a7z6 & V0y8v6));
assign C1y8v6 = (~(T2zet6 | S0zet6));
assign Wjx8v6 = (~(C7a7z6 & C1y8v6));
assign Kkx8v6 = (Dkx8v6 & Wjx8v6);
assign Ykx8v6 = (~(Rkx8v6 & Kkx8v6));
assign Jnx8v6 = (~(Ryyet6 & Ykx8v6));
assign Mlx8v6 = (~(K7a7z6 & Tzx8v6));
assign Flx8v6 = (~(S7a7z6 & A0y8v6));
assign Omx8v6 = (Mlx8v6 & Flx8v6);
assign Amx8v6 = (~(A8a7z6 & V0y8v6));
assign Tlx8v6 = (~(I8a7z6 & C1y8v6));
assign Hmx8v6 = (Amx8v6 & Tlx8v6);
assign Vmx8v6 = (~(Omx8v6 & Hmx8v6));
assign Cnx8v6 = (~(Vmx8v6 & W4y8v6));
assign Qnx8v6 = (~(Jnx8v6 & Cnx8v6));
assign Tsx8v6 = (~(Ean7z6[3] & Qnx8v6));
assign Eox8v6 = (~(Q8a7z6 & Tzx8v6));
assign Xnx8v6 = (~(Y8a7z6 & A0y8v6));
assign Gpx8v6 = (Eox8v6 & Xnx8v6);
assign Sox8v6 = (~(G9a7z6 & V0y8v6));
assign Lox8v6 = (~(Cco7v6 & C1y8v6));
assign Zox8v6 = (Sox8v6 & Lox8v6);
assign Npx8v6 = (~(Gpx8v6 & Zox8v6));
assign Yrx8v6 = (~(Npx8v6 & Ryyet6));
assign Bqx8v6 = (~(O9a7z6 & Tzx8v6));
assign Upx8v6 = (~(W9a7z6 & A0y8v6));
assign Drx8v6 = (Bqx8v6 & Upx8v6);
assign Pqx8v6 = (~(Eaa7z6 & V0y8v6));
assign Iqx8v6 = (~(Maa7z6 & C1y8v6));
assign Wqx8v6 = (Pqx8v6 & Iqx8v6);
assign Krx8v6 = (~(Drx8v6 & Wqx8v6));
assign Rrx8v6 = (~(Krx8v6 & W4y8v6));
assign Fsx8v6 = (~(Yrx8v6 & Rrx8v6));
assign Msx8v6 = (~(Fsx8v6 & K5y8v6));
assign Atx8v6 = (~(Tsx8v6 & Msx8v6));
assign P4y8v6 = (~(Ean7z6[4] & Atx8v6));
assign Otx8v6 = (~(Uaa7z6 & Tzx8v6));
assign Htx8v6 = (~(Cba7z6 & A0y8v6));
assign Qux8v6 = (Otx8v6 & Htx8v6);
assign Cux8v6 = (~(Kba7z6 & V0y8v6));
assign Vtx8v6 = (~(Jco7v6 & C1y8v6));
assign Jux8v6 = (Cux8v6 & Vtx8v6);
assign Xux8v6 = (~(Qux8v6 & Jux8v6));
assign Ixx8v6 = (~(Xux8v6 & Ryyet6));
assign Lvx8v6 = (~(Sba7z6 & Tzx8v6));
assign Evx8v6 = (~(Aca7z6 & A0y8v6));
assign Nwx8v6 = (Lvx8v6 & Evx8v6);
assign Zvx8v6 = (~(Ica7z6 & V0y8v6));
assign Svx8v6 = (~(Qca7z6 & C1y8v6));
assign Gwx8v6 = (Zvx8v6 & Svx8v6);
assign Uwx8v6 = (~(Nwx8v6 & Gwx8v6));
assign Bxx8v6 = (~(Uwx8v6 & W4y8v6));
assign Pxx8v6 = (~(Ixx8v6 & Bxx8v6));
assign U3y8v6 = (~(Pxx8v6 & Ean7z6[3]));
assign Dyx8v6 = (~(Yca7z6 & Tzx8v6));
assign Wxx8v6 = (~(Gda7z6 & A0y8v6));
assign Fzx8v6 = (Dyx8v6 & Wxx8v6);
assign Ryx8v6 = (~(Oda7z6 & V0y8v6));
assign Kyx8v6 = (~(Qco7v6 & C1y8v6));
assign Yyx8v6 = (Ryx8v6 & Kyx8v6);
assign Mzx8v6 = (~(Fzx8v6 & Yyx8v6));
assign Z2y8v6 = (~(Mzx8v6 & Ryyet6));
assign O0y8v6 = (~(Wda7z6 & Tzx8v6));
assign H0y8v6 = (~(Eea7z6 & A0y8v6));
assign E2y8v6 = (O0y8v6 & H0y8v6);
assign Q1y8v6 = (~(Mea7z6 & V0y8v6));
assign J1y8v6 = (~(Uea7z6 & C1y8v6));
assign X1y8v6 = (Q1y8v6 & J1y8v6);
assign L2y8v6 = (~(E2y8v6 & X1y8v6));
assign S2y8v6 = (~(L2y8v6 & W4y8v6));
assign G3y8v6 = (~(Z2y8v6 & S2y8v6));
assign N3y8v6 = (~(G3y8v6 & K5y8v6));
assign B4y8v6 = (U3y8v6 & N3y8v6);
assign I4y8v6 = (B4y8v6 | Ean7z6[4]);
assign Qxxet6 = (~(P4y8v6 & I4y8v6));
assign W4y8v6 = (!Ryyet6);
assign D5y8v6 = (!T2zet6);
assign K5y8v6 = (!Ean7z6[3]);
assign Cmy8v6 = (Hq27v6 & Or27v6);
assign Y5y8v6 = (~(Ies7z6[31] & Cmy8v6));
assign Jmy8v6 = (Hq27v6 & Fry8v6);
assign R5y8v6 = (~(Ies7z6[30] & Jmy8v6));
assign A7y8v6 = (Y5y8v6 & R5y8v6);
assign Eny8v6 = (~(Fry8v6 | Hq27v6));
assign M6y8v6 = (~(Ies7z6[29] & Eny8v6));
assign Lny8v6 = (~(Or27v6 | Hq27v6));
assign F6y8v6 = (~(Ies7z6[28] & Lny8v6));
assign T6y8v6 = (M6y8v6 & F6y8v6);
assign H7y8v6 = (~(A7y8v6 & T6y8v6));
assign S9y8v6 = (~(Ap27v6 & H7y8v6));
assign V7y8v6 = (~(Ies7z6[27] & Cmy8v6));
assign O7y8v6 = (~(Ies7z6[26] & Jmy8v6));
assign X8y8v6 = (V7y8v6 & O7y8v6);
assign J8y8v6 = (~(Ies7z6[25] & Eny8v6));
assign C8y8v6 = (~(Ies7z6[24] & Lny8v6));
assign Q8y8v6 = (J8y8v6 & C8y8v6);
assign E9y8v6 = (~(X8y8v6 & Q8y8v6));
assign L9y8v6 = (~(E9y8v6 & Mry8v6));
assign Z9y8v6 = (~(S9y8v6 & L9y8v6));
assign Cfy8v6 = (~(Tn27v6 & Z9y8v6));
assign Nay8v6 = (~(Ies7z6[23] & Cmy8v6));
assign Gay8v6 = (~(Ies7z6[22] & Jmy8v6));
assign Pby8v6 = (Nay8v6 & Gay8v6);
assign Bby8v6 = (~(Ies7z6[21] & Eny8v6));
assign Uay8v6 = (~(Ies7z6[20] & Lny8v6));
assign Iby8v6 = (Bby8v6 & Uay8v6);
assign Wby8v6 = (~(Pby8v6 & Iby8v6));
assign Hey8v6 = (~(Wby8v6 & Ap27v6));
assign Kcy8v6 = (~(Ies7z6[19] & Cmy8v6));
assign Dcy8v6 = (~(Ies7z6[18] & Jmy8v6));
assign Mdy8v6 = (Kcy8v6 & Dcy8v6);
assign Ycy8v6 = (~(Ies7z6[17] & Eny8v6));
assign Rcy8v6 = (~(Ies7z6[16] & Lny8v6));
assign Fdy8v6 = (Ycy8v6 & Rcy8v6);
assign Tdy8v6 = (~(Mdy8v6 & Fdy8v6));
assign Aey8v6 = (~(Tdy8v6 & Mry8v6));
assign Oey8v6 = (~(Hey8v6 & Aey8v6));
assign Vey8v6 = (~(Oey8v6 & Try8v6));
assign Jfy8v6 = (~(Cfy8v6 & Vey8v6));
assign Yqy8v6 = (~(Mm27v6 & Jfy8v6));
assign Xfy8v6 = (~(Ies7z6[15] & Cmy8v6));
assign Qfy8v6 = (~(Ies7z6[14] & Jmy8v6));
assign Zgy8v6 = (Xfy8v6 & Qfy8v6);
assign Lgy8v6 = (~(Ies7z6[13] & Eny8v6));
assign Egy8v6 = (~(Ies7z6[12] & Lny8v6));
assign Sgy8v6 = (Lgy8v6 & Egy8v6);
assign Ghy8v6 = (~(Zgy8v6 & Sgy8v6));
assign Rjy8v6 = (~(Ghy8v6 & Ap27v6));
assign Uhy8v6 = (~(Ies7z6[11] & Cmy8v6));
assign Nhy8v6 = (~(Ies7z6[10] & Jmy8v6));
assign Wiy8v6 = (Uhy8v6 & Nhy8v6);
assign Iiy8v6 = (~(Ies7z6[9] & Eny8v6));
assign Biy8v6 = (~(Ies7z6[8] & Lny8v6));
assign Piy8v6 = (Iiy8v6 & Biy8v6);
assign Djy8v6 = (~(Wiy8v6 & Piy8v6));
assign Kjy8v6 = (~(Djy8v6 & Mry8v6));
assign Yjy8v6 = (~(Rjy8v6 & Kjy8v6));
assign Dqy8v6 = (~(Yjy8v6 & Tn27v6));
assign Mky8v6 = (~(Ies7z6[7] & Cmy8v6));
assign Fky8v6 = (~(Ies7z6[6] & Jmy8v6));
assign Oly8v6 = (Mky8v6 & Fky8v6);
assign Aly8v6 = (~(Ies7z6[5] & Eny8v6));
assign Tky8v6 = (~(Ies7z6[4] & Lny8v6));
assign Hly8v6 = (Aly8v6 & Tky8v6);
assign Vly8v6 = (~(Oly8v6 & Hly8v6));
assign Ipy8v6 = (~(Vly8v6 & Ap27v6));
assign Xmy8v6 = (~(Ies7z6[3] & Cmy8v6));
assign Qmy8v6 = (~(Ies7z6[2] & Jmy8v6));
assign Noy8v6 = (Xmy8v6 & Qmy8v6);
assign Zny8v6 = (~(Ies7z6[1] & Eny8v6));
assign Sny8v6 = (~(Ies7z6[0] & Lny8v6));
assign Goy8v6 = (Zny8v6 & Sny8v6);
assign Uoy8v6 = (~(Noy8v6 & Goy8v6));
assign Bpy8v6 = (~(Uoy8v6 & Mry8v6));
assign Ppy8v6 = (~(Ipy8v6 & Bpy8v6));
assign Wpy8v6 = (~(Ppy8v6 & Try8v6));
assign Kqy8v6 = (Dqy8v6 & Wpy8v6);
assign Rqy8v6 = (Kqy8v6 | Mm27v6);
assign Fl27v6 = (~(Yqy8v6 & Rqy8v6));
assign Fry8v6 = (!Or27v6);
assign Mry8v6 = (!Ap27v6);
assign Try8v6 = (!Tn27v6);
assign P209v6 = (~(Znn7z6[3] | Znn7z6[2]));
assign Hsy8v6 = (~(V3pet6 & P209v6));
assign I209v6 = (~(Znn7z6[1] | Znn7z6[3]));
assign Lfz8v6 = (Znn7z6[2] & I209v6);
assign Asy8v6 = (~(Bgpet6 & Lfz8v6));
assign Euy8v6 = (Hsy8v6 & Asy8v6);
assign Z009v6 = (~(Znn7z6[2] | D309v6));
assign Z8z8v6 = (Z009v6 & F409v6);
assign Cty8v6 = (~(Hspet6 & Z8z8v6));
assign Ivz8v6 = (~(R309v6 | D309v6));
assign Osy8v6 = (~(F409v6 | R309v6));
assign G109v6 = (Ivz8v6 | Osy8v6);
assign Vsy8v6 = (~(W2n7z6[0] & G109v6));
assign Qty8v6 = (Cty8v6 & Vsy8v6);
assign C7z8v6 = (Znn7z6[1] & Z009v6);
assign Jty8v6 = (~(N4qet6 & C7z8v6));
assign Xty8v6 = (Qty8v6 & Jty8v6);
assign Proet6 = (~(Euy8v6 & Xty8v6));
assign Suy8v6 = (~(U1pet6 & P209v6));
assign Luy8v6 = (~(Aepet6 & Lfz8v6));
assign Iwy8v6 = (Suy8v6 & Luy8v6);
assign Gvy8v6 = (~(Gqpet6 & Z8z8v6));
assign Zuy8v6 = (~(W2n7z6[1] & G109v6));
assign Uvy8v6 = (Gvy8v6 & Zuy8v6);
assign Nvy8v6 = (~(M2qet6 & C7z8v6));
assign Bwy8v6 = (Uvy8v6 & Nvy8v6);
assign Opoet6 = (~(Iwy8v6 & Bwy8v6));
assign Wwy8v6 = (~(Zbpet6 & P209v6));
assign Pwy8v6 = (~(Fopet6 & Lfz8v6));
assign Myy8v6 = (Wwy8v6 & Pwy8v6);
assign Kxy8v6 = (~(L0qet6 & Z8z8v6));
assign Dxy8v6 = (~(J5n7z6[0] & G109v6));
assign Yxy8v6 = (Kxy8v6 & Dxy8v6);
assign Rxy8v6 = (~(Rcqet6 & C7z8v6));
assign Fyy8v6 = (Yxy8v6 & Rxy8v6);
assign Tzoet6 = (~(Myy8v6 & Fyy8v6));
assign Azy8v6 = (~(Y9pet6 & P209v6));
assign Tyy8v6 = (~(Empet6 & Lfz8v6));
assign Q0z8v6 = (Azy8v6 & Tyy8v6);
assign Ozy8v6 = (~(Kypet6 & Z8z8v6));
assign Hzy8v6 = (~(J5n7z6[1] & G109v6));
assign C0z8v6 = (Ozy8v6 & Hzy8v6);
assign Vzy8v6 = (~(Qaqet6 & C7z8v6));
assign J0z8v6 = (C0z8v6 & Vzy8v6);
assign Sxoet6 = (~(Q0z8v6 & J0z8v6));
assign E1z8v6 = (~(X7pet6 & P209v6));
assign X0z8v6 = (~(Dkpet6 & Lfz8v6));
assign U2z8v6 = (E1z8v6 & X0z8v6);
assign S1z8v6 = (~(Jwpet6 & Z8z8v6));
assign L1z8v6 = (~(J5n7z6[2] & G109v6));
assign G2z8v6 = (S1z8v6 & L1z8v6);
assign Z1z8v6 = (~(P8qet6 & C7z8v6));
assign N2z8v6 = (G2z8v6 & Z1z8v6);
assign Rvoet6 = (~(U2z8v6 & N2z8v6));
assign I3z8v6 = (~(W5pet6 & P209v6));
assign B3z8v6 = (~(Cipet6 & Lfz8v6));
assign Y4z8v6 = (I3z8v6 & B3z8v6);
assign W3z8v6 = (~(Iupet6 & Z8z8v6));
assign P3z8v6 = (~(J5n7z6[3] & G109v6));
assign K4z8v6 = (W3z8v6 & P3z8v6);
assign D4z8v6 = (~(O6qet6 & C7z8v6));
assign R4z8v6 = (K4z8v6 & D4z8v6);
assign Qtoet6 = (~(Y4z8v6 & R4z8v6));
assign M5z8v6 = (~(Yotet6 & P209v6));
assign F5z8v6 = (~(Dztet6 & Lfz8v6));
assign V6z8v6 = (M5z8v6 & F5z8v6);
assign H6z8v6 = (~(Qvm7z6[0] & Ivz8v6));
assign T5z8v6 = (~(R309v6 | Znn7z6[3]));
assign Waz8v6 = (T5z8v6 & Znn7z6[1]);
assign A6z8v6 = (~(X9yet6 & Waz8v6));
assign O6z8v6 = (H6z8v6 & A6z8v6);
assign X5set6 = (~(V6z8v6 & O6z8v6));
assign Q7z8v6 = (~(Cxtet6 & Lfz8v6));
assign J7z8v6 = (~(Eia7z6 & C7z8v6));
assign E8z8v6 = (Q7z8v6 & J7z8v6);
assign X7z8v6 = (~(Xmtet6 & P209v6));
assign Baz8v6 = (E8z8v6 & X7z8v6);
assign S8z8v6 = (~(Qvm7z6[1] & Ivz8v6));
assign L8z8v6 = (~(Icyet6 & Waz8v6));
assign N9z8v6 = (S8z8v6 & L8z8v6);
assign G9z8v6 = (~(Mia7z6 & Z8z8v6));
assign U9z8v6 = (N9z8v6 & G9z8v6);
assign W3set6 = (~(Baz8v6 & U9z8v6));
assign Paz8v6 = (~(Wktet6 & P209v6));
assign Iaz8v6 = (~(Bvtet6 & Lfz8v6));
assign Ybz8v6 = (Paz8v6 & Iaz8v6);
assign Kbz8v6 = (~(Hjn7z6[7] & Ivz8v6));
assign Xzz8v6 = (Z009v6 | Waz8v6);
assign Dbz8v6 = (~(T2zet6 & Xzz8v6));
assign Rbz8v6 = (Kbz8v6 & Dbz8v6);
assign V1set6 = (~(Ybz8v6 & Rbz8v6));
assign Fcz8v6 = (~(Hjn7z6[8] & Ivz8v6));
assign Odz8v6 = (Fcz8v6 & K309v6);
assign Mcz8v6 = (F409v6 | Znn7z6[3]);
assign Cez8v6 = (~(Znn7z6[2] & Mcz8v6));
assign Adz8v6 = (~(S0zet6 & Cez8v6));
assign Tcz8v6 = (~(Attet6 & I209v6));
assign Hdz8v6 = (Adz8v6 & Tcz8v6);
assign Uzret6 = (~(Odz8v6 & Hdz8v6));
assign Vdz8v6 = (~(Hjn7z6[9] & Ivz8v6));
assign Efz8v6 = (Vdz8v6 & K309v6);
assign Qez8v6 = (~(Ryyet6 & Cez8v6));
assign Jez8v6 = (~(Zqtet6 & I209v6));
assign Xez8v6 = (Qez8v6 & Jez8v6);
assign Txret6 = (~(Efz8v6 & Xez8v6));
assign Zfz8v6 = (~(Hjn7z6[5] & Xzz8v6));
assign E009v6 = (P209v6 | Lfz8v6);
assign Sfz8v6 = (~(Vitet6 & E009v6));
assign Ngz8v6 = (Zfz8v6 & Sfz8v6);
assign Ggz8v6 = (~(Hjn7z6[10] & Ivz8v6));
assign Svret6 = (~(Ngz8v6 & Ggz8v6));
assign Bhz8v6 = (~(Hjn7z6[6] & Xzz8v6));
assign Ugz8v6 = (~(Ugtet6 & E009v6));
assign Phz8v6 = (Bhz8v6 & Ugz8v6);
assign Ihz8v6 = (~(Hjn7z6[11] & Ivz8v6));
assign Rtret6 = (~(Phz8v6 & Ihz8v6));
assign Diz8v6 = (~(Hjn7z6[7] & Xzz8v6));
assign Whz8v6 = (~(Tetet6 & E009v6));
assign Riz8v6 = (Diz8v6 & Whz8v6);
assign Kiz8v6 = (~(Hjn7z6[12] & Ivz8v6));
assign Qrret6 = (~(Riz8v6 & Kiz8v6));
assign Fjz8v6 = (~(Hjn7z6[8] & Xzz8v6));
assign Yiz8v6 = (~(Sctet6 & E009v6));
assign Tjz8v6 = (Fjz8v6 & Yiz8v6);
assign Mjz8v6 = (~(Hjn7z6[13] & Ivz8v6));
assign Ppret6 = (~(Tjz8v6 & Mjz8v6));
assign Hkz8v6 = (~(Hjn7z6[9] & Xzz8v6));
assign Akz8v6 = (~(Ratet6 & E009v6));
assign Vkz8v6 = (Hkz8v6 & Akz8v6);
assign Okz8v6 = (~(Hjn7z6[14] & Ivz8v6));
assign Onret6 = (~(Vkz8v6 & Okz8v6));
assign Jlz8v6 = (~(Hjn7z6[10] & Xzz8v6));
assign Clz8v6 = (~(Q8tet6 & E009v6));
assign Xlz8v6 = (Jlz8v6 & Clz8v6);
assign Qlz8v6 = (~(Hjn7z6[15] & Ivz8v6));
assign Nlret6 = (~(Xlz8v6 & Qlz8v6));
assign Lmz8v6 = (~(Hjn7z6[11] & Xzz8v6));
assign Emz8v6 = (~(P6tet6 & E009v6));
assign Zmz8v6 = (Lmz8v6 & Emz8v6);
assign Smz8v6 = (~(Hjn7z6[16] & Ivz8v6));
assign Mjret6 = (~(Zmz8v6 & Smz8v6));
assign Nnz8v6 = (~(Hjn7z6[12] & Xzz8v6));
assign Gnz8v6 = (~(O4tet6 & E009v6));
assign Boz8v6 = (Nnz8v6 & Gnz8v6);
assign Unz8v6 = (~(Hjn7z6[17] & Ivz8v6));
assign Lhret6 = (~(Boz8v6 & Unz8v6));
assign Poz8v6 = (~(Hjn7z6[13] & Xzz8v6));
assign Ioz8v6 = (~(N2tet6 & E009v6));
assign Dpz8v6 = (Poz8v6 & Ioz8v6);
assign Woz8v6 = (~(Hjn7z6[18] & Ivz8v6));
assign Kfret6 = (~(Dpz8v6 & Woz8v6));
assign Rpz8v6 = (~(Hjn7z6[14] & Xzz8v6));
assign Kpz8v6 = (~(M0tet6 & E009v6));
assign Fqz8v6 = (Rpz8v6 & Kpz8v6);
assign Ypz8v6 = (~(Hjn7z6[19] & Ivz8v6));
assign Jdret6 = (~(Fqz8v6 & Ypz8v6));
assign Tqz8v6 = (~(Hjn7z6[15] & Xzz8v6));
assign Mqz8v6 = (~(Lyset6 & E009v6));
assign Hrz8v6 = (Tqz8v6 & Mqz8v6);
assign Arz8v6 = (~(Hjn7z6[20] & Ivz8v6));
assign Ibret6 = (~(Hrz8v6 & Arz8v6));
assign Vrz8v6 = (~(Hjn7z6[16] & Xzz8v6));
assign Orz8v6 = (~(Kwset6 & E009v6));
assign Jsz8v6 = (Vrz8v6 & Orz8v6);
assign Csz8v6 = (~(Hjn7z6[21] & Ivz8v6));
assign H9ret6 = (~(Jsz8v6 & Csz8v6));
assign Xsz8v6 = (~(Hjn7z6[17] & Xzz8v6));
assign Qsz8v6 = (~(Juset6 & E009v6));
assign Ltz8v6 = (Xsz8v6 & Qsz8v6);
assign Etz8v6 = (~(Hjn7z6[22] & Ivz8v6));
assign G7ret6 = (~(Ltz8v6 & Etz8v6));
assign Ztz8v6 = (~(Hjn7z6[18] & Xzz8v6));
assign Stz8v6 = (~(Isset6 & E009v6));
assign Nuz8v6 = (Ztz8v6 & Stz8v6);
assign Guz8v6 = (~(Hjn7z6[23] & Ivz8v6));
assign F5ret6 = (~(Nuz8v6 & Guz8v6));
assign Bvz8v6 = (~(Hjn7z6[19] & Xzz8v6));
assign Uuz8v6 = (~(Hqset6 & E009v6));
assign Wvz8v6 = (Bvz8v6 & Uuz8v6);
assign Pvz8v6 = (~(Hjn7z6[24] & Ivz8v6));
assign E3ret6 = (~(Wvz8v6 & Pvz8v6));
assign Kwz8v6 = (~(Hjn7z6[20] & Xzz8v6));
assign Dwz8v6 = (~(Goset6 & E009v6));
assign D1ret6 = (~(Kwz8v6 & Dwz8v6));
assign Ywz8v6 = (~(Hjn7z6[21] & Xzz8v6));
assign Rwz8v6 = (~(Fmset6 & E009v6));
assign Czqet6 = (~(Ywz8v6 & Rwz8v6));
assign Mxz8v6 = (~(Hjn7z6[22] & Xzz8v6));
assign Fxz8v6 = (~(Ekset6 & E009v6));
assign Bxqet6 = (~(Mxz8v6 & Fxz8v6));
assign Ayz8v6 = (~(Hjn7z6[23] & Xzz8v6));
assign Txz8v6 = (~(Diset6 & E009v6));
assign Avqet6 = (~(Ayz8v6 & Txz8v6));
assign Oyz8v6 = (~(Hjn7z6[24] & Xzz8v6));
assign Hyz8v6 = (~(Cgset6 & E009v6));
assign Zsqet6 = (~(Oyz8v6 & Hyz8v6));
assign Czz8v6 = (~(Hjn7z6[25] & Xzz8v6));
assign Vyz8v6 = (~(Beset6 & E009v6));
assign Yqqet6 = (~(Czz8v6 & Vyz8v6));
assign Qzz8v6 = (~(Hjn7z6[26] & Xzz8v6));
assign Jzz8v6 = (~(Acset6 & E009v6));
assign Xoqet6 = (~(Qzz8v6 & Jzz8v6));
assign S009v6 = (~(Hjn7z6[27] & Xzz8v6));
assign L009v6 = (~(Z9set6 & E009v6));
assign Wmqet6 = (~(S009v6 & L009v6));
assign N109v6 = (G109v6 | Z009v6);
assign B209v6 = (~(Hjn7z6[28] & N109v6));
assign U109v6 = (Sr97z6 | N109v6);
assign Vkqet6 = (~(B209v6 & U109v6));
assign W209v6 = (P209v6 | I209v6);
assign Uiqet6 = (W209v6 | Hjn7z6[29]);
assign Tgqet6 = (Hjn7z6[30] & Y309v6);
assign Seqet6 = (Hjn7z6[31] & Y309v6);
assign D309v6 = (!Znn7z6[3]);
assign K309v6 = (!P209v6);
assign R309v6 = (!Znn7z6[2]);
assign Y309v6 = (!W209v6);
assign F409v6 = (!Znn7z6[1]);
assign Ra09v6 = (~(Gf09v6 | Yo37v6));
assign T409v6 = (~(Iuvmz6[5] & Ra09v6));
assign Ya09v6 = (~(M6s7z6[1] | Yo37v6));
assign M409v6 = (~(Iuvmz6[7] & Ya09v6));
assign Jd09v6 = (T409v6 & M409v6);
assign V509v6 = (Ze09v6 | Jd09v6);
assign H509v6 = (~(Iuvmz6[6] & Ra09v6));
assign A509v6 = (~(Iuvmz6[8] & Ya09v6));
assign L709v6 = (H509v6 & A509v6);
assign O509v6 = (L709v6 | M6s7z6[0]);
assign Q609v6 = (V509v6 & O509v6);
assign C609v6 = (~(M6s7z6[0] | M6s7z6[1]));
assign Ee09v6 = (C609v6 & Yo37v6);
assign J609v6 = (~(Ee09v6 & Iuvmz6[4]));
assign Nks7z6[0] = (~(Q609v6 & J609v6));
assign E709v6 = (~(Iuvmz6[7] & Ra09v6));
assign X609v6 = (~(Iuvmz6[4] & Ya09v6));
assign I909v6 = (E709v6 & X609v6);
assign Z709v6 = (I909v6 | M6s7z6[0]);
assign S709v6 = (L709v6 | Ze09v6);
assign N809v6 = (Z709v6 & S709v6);
assign G809v6 = (~(Ee09v6 & Iuvmz6[5]));
assign Nks7z6[1] = (~(N809v6 & G809v6));
assign B909v6 = (~(Iuvmz6[8] & Ra09v6));
assign U809v6 = (~(Iuvmz6[5] & Ya09v6));
assign Tb09v6 = (B909v6 & U809v6);
assign W909v6 = (Tb09v6 | M6s7z6[0]);
assign P909v6 = (I909v6 | Ze09v6);
assign Ka09v6 = (W909v6 & P909v6);
assign Da09v6 = (~(Ee09v6 & Iuvmz6[6]));
assign Nks7z6[2] = (~(Ka09v6 & Da09v6));
assign Mb09v6 = (~(Iuvmz6[4] & Ra09v6));
assign Fb09v6 = (~(Iuvmz6[6] & Ya09v6));
assign Cd09v6 = (Mb09v6 & Fb09v6);
assign Hc09v6 = (Cd09v6 | M6s7z6[0]);
assign Ac09v6 = (Tb09v6 | Ze09v6);
assign Vc09v6 = (Hc09v6 & Ac09v6);
assign Oc09v6 = (~(Ee09v6 & Iuvmz6[7]));
assign Nks7z6[3] = (~(Vc09v6 & Oc09v6));
assign Xd09v6 = (Ze09v6 | Cd09v6);
assign Qd09v6 = (Jd09v6 | M6s7z6[0]);
assign Se09v6 = (Xd09v6 & Qd09v6);
assign Le09v6 = (~(Iuvmz6[8] & Ee09v6));
assign Nks7z6[4] = (~(Se09v6 & Le09v6));
assign Ze09v6 = (!M6s7z6[0]);
assign Gf09v6 = (!M6s7z6[1]);
assign Fkwmv6 = (~(Vzwmv6 | Fqxmz6[3]));
assign Xmwmv6 = (~(K3a7z6 | Fqxmz6[4]));
assign Nf09v6 = (Fqxmz6[2] | Fqxmz6[4]);
assign Bxvmv6 = (I3xmv6 & Nf09v6);
assign Zovmv6 = (~(K3a7z6 | Fqxmz6[2]));
assign Djwmv6 = (Bxvmv6 | Zovmv6);
assign Piwmv6 = (~(G2xmv6 | Q0xmv6));
assign O0wmv6 = (C0xmv6 | Piwmv6);
assign Uf09v6 = (O0wmv6 | Zovmv6);
assign S9wmv6 = (Fqxmz6[5] & Uf09v6);
assign Xuvmv6 = (Djwmv6 & S9wmv6);
assign Qnvmv6 = (~(Fkwmv6 & Xuvmv6));
assign Tkwmv6 = (~(Fqxmz6[0] | E1xmv6));
assign Xnvmv6 = (~(Uia7z6 | Q0xmv6));
assign Bg09v6 = (C0xmv6 | Z1xmv6);
assign Ig09v6 = (~(Fqxmz6[5] & Bg09v6));
assign Oswmv6 = (~(Piwmv6 & Fqxmz6[4]));
assign Lgwmv6 = (Ig09v6 & Oswmv6);
assign Pg09v6 = (SWDITMS | Q0xmv6);
assign Cnvmv6 = (~(Pg09v6 & K4xmv6));
assign Alwmv6 = (~(C0xmv6 & Cnvmv6));
assign Jnvmv6 = (~(Lgwmv6 & Alwmv6));
assign Wbwmv6 = (~(Tkwmv6 & Jnvmv6));
assign Fsvmv6 = (Qnvmv6 & Wbwmv6);
assign K5wmv6 = (~(Fqxmz6[3] | Fqxmz6[0]));
assign Lovmv6 = (~(S1xmv6 | Zovmv6));
assign Eovmv6 = (Xnvmv6 | Zovmv6);
assign Tsvmv6 = (Fqxmz6[4] & Eovmv6);
assign D5wmv6 = (Lovmv6 & W3xmv6);
assign A0wmv6 = (~(B3xmv6 | D5wmv6));
assign Sovmv6 = (~(Djwmv6 & A0wmv6));
assign Wqvmv6 = (~(K5wmv6 & Sovmv6));
assign Ghwmv6 = (~(Vzwmv6 | E1xmv6));
assign Iqvmv6 = (~(S1xmv6 | L1xmv6));
assign Upvmv6 = (Fqxmz6[4] | SWDITMS);
assign Gpvmv6 = (~(C0xmv6 | Zovmv6));
assign Npvmv6 = (~(Gpvmv6 & Z1xmv6));
assign Bqvmv6 = (~(Upvmv6 & Npvmv6));
assign Pqvmv6 = (~(Iqvmv6 & Bqvmv6));
assign Rrvmv6 = (Wqvmv6 & Pqvmv6);
assign Drvmv6 = (Fkwmv6 | Ghwmv6);
assign Krvmv6 = (~(Drvmv6 & B3xmv6));
assign Yrvmv6 = (Rrvmv6 & Krvmv6);
assign Msvmv6 = (~(Fsvmv6 & Yrvmv6));
assign Nwvmv6 = (~(Msvmv6 & J0xmv6));
assign Atvmv6 = (~(Tsvmv6 | S1xmv6));
assign Suwmv6 = (~(Atvmv6 & Alwmv6));
assign Aewmv6 = (~(Oswmv6 & Suwmv6));
assign Cuvmv6 = (~(Aewmv6 & Fkwmv6));
assign Otvmv6 = (~(Alwmv6 & E1xmv6));
assign Htvmv6 = (E1xmv6 | Xmwmv6);
assign Bwwmv6 = (Otvmv6 & Htvmv6);
assign Uwvmv6 = (U2xmv6 | Bwwmv6);
assign Vtvmv6 = (~(Uwvmv6 & Vzwmv6));
assign Zvvmv6 = (Cuvmv6 & Vtvmv6);
assign Aswmv6 = (~(Q0xmv6 | Fqxmz6[4]));
assign Juvmv6 = (~(Us47v6 & Aswmv6));
assign Quvmv6 = (~(Juvmv6 & Oswmv6));
assign Evvmv6 = (~(S1xmv6 & Quvmv6));
assign Lvvmv6 = (~(Evvmv6 & D4xmv6));
assign Svvmv6 = (~(Ghwmv6 & Lvvmv6));
assign Gwvmv6 = (Zvvmv6 & Svvmv6);
assign Mzvmv6 = (Gwvmv6 | J0xmv6);
assign Woxmz6[0] = (~(Nwvmv6 & Mzvmv6));
assign Dyvmv6 = (~(Fqxmz6[0] & Uwvmv6));
assign Dcwmv6 = (~(Bxvmv6 & O0wmv6));
assign Ixvmv6 = (S1xmv6 | Dcwmv6);
assign Pxvmv6 = (~(Oswmv6 & Ixvmv6));
assign Wxvmv6 = (~(Pxvmv6 & E1xmv6));
assign Ryvmv6 = (Dyvmv6 & Wxvmv6);
assign Kyvmv6 = (~(Aewmv6 & Fqxmz6[3]));
assign Yyvmv6 = (~(Ryvmv6 & Kyvmv6));
assign Fzvmv6 = (~(Yyvmv6 & J0xmv6));
assign Woxmz6[1] = (~(Mzvmv6 & Fzvmv6));
assign Tzvmv6 = (I3xmv6 | Q0xmv6);
assign Hewmv6 = (~(A0wmv6 & Tzvmv6));
assign Z2wmv6 = (~(Hewmv6 & Tkwmv6));
assign Qtwmv6 = (K4xmv6 | Fqxmz6[4]);
assign H0wmv6 = (X0xmv6 | Us47v6);
assign V0wmv6 = (Qtwmv6 & H0wmv6);
assign C1wmv6 = (~(V0wmv6 & O0wmv6));
assign L2wmv6 = (~(C1wmv6 & S1xmv6));
assign X1wmv6 = (~(S1xmv6 | Q0xmv6));
assign J1wmv6 = (C0xmv6 | Uia7z6);
assign Q1wmv6 = (~(I3xmv6 & J1wmv6));
assign E2wmv6 = (~(X1wmv6 & Q1wmv6));
assign S2wmv6 = (L2wmv6 & E2wmv6);
assign Cfwmv6 = (~(S2wmv6 & Ghwmv6));
assign M6wmv6 = (Z2wmv6 & Cfwmv6);
assign I4wmv6 = (I3xmv6 | Fqxmz6[2]);
assign G3wmv6 = (G2xmv6 | C0xmv6);
assign N3wmv6 = (G3wmv6 & I3xmv6);
assign U3wmv6 = (~(N3wmv6 & Fqxmz6[2]));
assign B4wmv6 = (~(U3wmv6 & Fqxmz6[5]));
assign P4wmv6 = (I4wmv6 & B4wmv6);
assign W4wmv6 = (~(P4wmv6 & Oswmv6));
assign Y5wmv6 = (~(W4wmv6 & Fkwmv6));
assign A7wmv6 = (P3xmv6 | D5wmv6);
assign R5wmv6 = (~(K5wmv6 & A7wmv6));
assign F6wmv6 = (Y5wmv6 & R5wmv6);
assign T6wmv6 = (~(M6wmv6 & F6wmv6));
assign Pbwmv6 = (~(T6wmv6 & Fqxmz6[1]));
assign E9wmv6 = (~(Hewmv6 & Ghwmv6));
assign J8wmv6 = (~(A7wmv6 & Fqxmz6[3]));
assign H7wmv6 = (SWDITMS | Fqxmz6[5]);
assign O7wmv6 = (~(H7wmv6 & Aswmv6));
assign V7wmv6 = (~(Oswmv6 & O7wmv6));
assign C8wmv6 = (~(V7wmv6 & E1xmv6));
assign Q8wmv6 = (~(J8wmv6 & C8wmv6));
assign X8wmv6 = (~(Q8wmv6 & Vzwmv6));
assign Uawmv6 = (E9wmv6 & X8wmv6);
assign L9wmv6 = (Fqxmz6[2] | SWDITMS);
assign Z9wmv6 = (~(S9wmv6 & L9wmv6));
assign Gawmv6 = (~(Z9wmv6 & Dcwmv6));
assign Nawmv6 = (~(Fkwmv6 & Gawmv6));
assign Bbwmv6 = (~(Uawmv6 & Nawmv6));
assign Ibwmv6 = (~(Bbwmv6 & J0xmv6));
assign Woxmz6[2] = (~(Pbwmv6 & Ibwmv6));
assign Mdwmv6 = (Wbwmv6 & Oswmv6);
assign Ycwmv6 = (Vzwmv6 | D4xmv6);
assign Kcwmv6 = (~(Dcwmv6 | Fqxmz6[0]));
assign Rcwmv6 = (~(Kcwmv6 & Fqxmz6[5]));
assign Fdwmv6 = (Ycwmv6 & Rcwmv6);
assign Tdwmv6 = (~(Mdwmv6 & Fdwmv6));
assign Egwmv6 = (~(Tdwmv6 & J0xmv6));
assign Vewmv6 = (~(Aewmv6 & Vzwmv6));
assign Oewmv6 = (~(Hewmv6 & Fkwmv6));
assign Jfwmv6 = (Vewmv6 & Oewmv6);
assign Qfwmv6 = (~(Jfwmv6 & Cfwmv6));
assign Xfwmv6 = (~(Qfwmv6 & Fqxmz6[1]));
assign Iiwmv6 = (Egwmv6 & Xfwmv6);
assign Zgwmv6 = (Tkwmv6 | J0xmv6);
assign Sgwmv6 = (~(Lgwmv6 & I3xmv6));
assign Uhwmv6 = (Zgwmv6 & Sgwmv6);
assign Nhwmv6 = (Ghwmv6 | Fqxmz6[1]);
assign Biwmv6 = (~(Uhwmv6 & Nhwmv6));
assign Woxmz6[3] = (~(Iiwmv6 & Biwmv6));
assign Wiwmv6 = (Cja7z6 & Q0xmv6);
assign Lnwmv6 = (~(Wiwmv6 | Piwmv6));
assign Frwmv6 = (C0xmv6 | Lnwmv6);
assign Kjwmv6 = (~(Djwmv6 & Frwmv6));
assign Rjwmv6 = (~(Kjwmv6 & S1xmv6));
assign Yjwmv6 = (~(D4xmv6 & Rjwmv6));
assign Qmwmv6 = (~(Fkwmv6 & Yjwmv6));
assign Uvwmv6 = (~(S1xmv6 | W3xmv6));
assign Mkwmv6 = (~(C0xmv6 | Fqxmz6[5]));
assign Iwwmv6 = (Mkwmv6 & Lnwmv6);
assign Cmwmv6 = (~(Uvwmv6 | Iwwmv6));
assign Olwmv6 = (L1xmv6 | Xmwmv6);
assign Hlwmv6 = (~(Alwmv6 & Tkwmv6));
assign Vlwmv6 = (~(Olwmv6 & Hlwmv6));
assign Jmwmv6 = (~(Cmwmv6 & Vlwmv6));
assign Ppwmv6 = (Qmwmv6 & Jmwmv6);
assign Enwmv6 = (~(Xmwmv6 | Fqxmz6[3]));
assign Bpwmv6 = (Enwmv6 & Vzwmv6);
assign Znwmv6 = (N2xmv6 | K3a7z6);
assign Snwmv6 = (~(Frwmv6 & X0xmv6));
assign Nowmv6 = (Znwmv6 & Snwmv6);
assign Gowmv6 = (P3xmv6 | S1xmv6);
assign Uowmv6 = (Nowmv6 & Gowmv6);
assign Ipwmv6 = (~(Bpwmv6 & Uowmv6));
assign Wpwmv6 = (~(Ppwmv6 & Ipwmv6));
assign Fywmv6 = (~(Wpwmv6 & J0xmv6));
assign Dqwmv6 = (~(Fqxmz6[4] | SWDITMS));
assign Yqwmv6 = (~(Dqwmv6 & E1xmv6));
assign Kqwmv6 = (Aswmv6 & Fqxmz6[3]);
assign Rqwmv6 = (~(Kqwmv6 & Qr47v6));
assign Mrwmv6 = (Yqwmv6 & Rqwmv6);
assign Trwmv6 = (~(Mrwmv6 & Frwmv6));
assign Luwmv6 = (~(Trwmv6 & S1xmv6));
assign Hswmv6 = (~(Mq47v6 & Aswmv6));
assign Vswmv6 = (Hswmv6 & K4xmv6);
assign Ctwmv6 = (~(Vswmv6 & Oswmv6));
assign Jtwmv6 = (~(Ctwmv6 & Fqxmz6[5]));
assign Xtwmv6 = (~(Qtwmv6 & Jtwmv6));
assign Euwmv6 = (~(Xtwmv6 & Fqxmz6[3]));
assign Gvwmv6 = (Luwmv6 & Euwmv6);
assign Zuwmv6 = (Suwmv6 | Fqxmz6[3]);
assign Nvwmv6 = (~(Gvwmv6 & Zuwmv6));
assign Kxwmv6 = (~(Nvwmv6 & Fqxmz6[0]));
assign Wwwmv6 = (~(Bwwmv6 | Uvwmv6));
assign Pwwmv6 = (~(Iwwmv6 | Fqxmz6[0]));
assign Dxwmv6 = (~(Wwwmv6 & Pwwmv6));
assign Rxwmv6 = (~(Kxwmv6 & Dxwmv6));
assign Yxwmv6 = (~(Rxwmv6 & Fqxmz6[1]));
assign Woxmz6[4] = (~(Fywmv6 & Yxwmv6));
assign Tywmv6 = (~(K3a7z6 | Q0xmv6));
assign Mywmv6 = (~(J0xmv6 | L1xmv6));
assign Azwmv6 = (~(Tywmv6 & Mywmv6));
assign Ozwmv6 = (Azwmv6 ^ Fqxmz6[5]);
assign Hzwmv6 = (C0xmv6 | Q0xmv6);
assign Woxmz6[5] = (~(Ozwmv6 & Hzwmv6));
assign Vzwmv6 = (!Fqxmz6[0]);
assign C0xmv6 = (!Fqxmz6[4]);
assign J0xmv6 = (!Fqxmz6[1]);
assign Q0xmv6 = (!Fqxmz6[2]);
assign X0xmv6 = (!Aswmv6);
assign E1xmv6 = (!Fqxmz6[3]);
assign L1xmv6 = (!Ghwmv6);
assign S1xmv6 = (!Fqxmz6[5]);
assign Z1xmv6 = (!Xnvmv6);
assign G2xmv6 = (!Uia7z6);
assign N2xmv6 = (!Lnwmv6);
assign U2xmv6 = (!Lgwmv6);
assign B3xmv6 = (!Oswmv6);
assign I3xmv6 = (!Xmwmv6);
assign P3xmv6 = (!Dcwmv6);
assign W3xmv6 = (!Tsvmv6);
assign D4xmv6 = (!Xuvmv6);
assign K4xmv6 = (!Zovmv6);
assign Fn0nv6 = (~(O21nv6 | R01nv6));
assign Xw0nv6 = (~(Dwb7z6[3] | Dwb7z6[1]));
assign C6ymv6 = (~(Fn0nv6 | Xw0nv6));
assign Y4xmv6 = (X31nv6 | Y01nv6);
assign Jw0nv6 = (~(Y01nv6 | M11nv6));
assign R4xmv6 = (~(Jjzdt6 & Jw0nv6));
assign F5xmv6 = (Y4xmv6 & R4xmv6);
assign Khymv6 = (~(O21nv6 | Dwb7z6[2]));
assign Ym0nv6 = (~(R01nv6 | J31nv6));
assign X7xmv6 = (F5xmv6 & Q31nv6);
assign Ayxmv6 = (Xw0nv6 & Y01nv6);
assign Hv0nv6 = (Ayxmv6 & Z41nv6);
assign A6xmv6 = (~(Li0et6 & Hv0nv6));
assign Gr0nv6 = (Dwb7z6[3] & O21nv6);
assign Ynzmv6 = (~(Z41nv6 & Gr0nv6));
assign Cp0nv6 = (~(O21nv6 | Dwb7z6[3]));
assign M5xmv6 = (I61nv6 | Cp0nv6);
assign T5xmv6 = (~(M5xmv6 & Iga7z6));
assign J7xmv6 = (A6xmv6 & T5xmv6);
assign W8zmv6 = (~(Y01nv6 | Dwb7z6[0]));
assign Ci0nv6 = (~(Z41nv6 | Dwb7z6[2]));
assign N60nv6 = (W8zmv6 | Ci0nv6);
assign H6xmv6 = (N60nv6 | Gvydt6);
assign V6xmv6 = (~(H6xmv6 & Fn0nv6));
assign Sj0nv6 = (Dwb7z6[0] & Gr0nv6);
assign O6xmv6 = (~(Sj0nv6 & A4zdt6));
assign C7xmv6 = (V6xmv6 & O6xmv6);
assign Q7xmv6 = (J7xmv6 & C7xmv6);
assign E8xmv6 = (~(X7xmv6 & Q7xmv6));
assign Ie0nv6 = (~(K01nv6 | Dwb7z6[5]));
assign Lfxmv6 = (~(E8xmv6 & Ie0nv6));
assign L8xmv6 = (M11nv6 | N60nv6);
assign Syzmv6 = (Dwb7z6[2] & Dwb7z6[1]);
assign Apzmv6 = (Syzmv6 & Dwb7z6[3]);
assign Oa0nv6 = (~(Dwb7z6[0] & Apzmv6));
assign S8xmv6 = (L8xmv6 & Oa0nv6);
assign Z8xmv6 = (~(S8xmv6 & Ynzmv6));
assign N9xmv6 = (~(Ys97z6 & Z8xmv6));
assign Uszmv6 = (Ym0nv6 & Z41nv6);
assign G9xmv6 = (~(If1et6 & Uszmv6));
assign Baxmv6 = (N9xmv6 & G9xmv6);
assign Nr0nv6 = (~(Dwb7z6[3] | J31nv6));
assign U9xmv6 = (~(L32et6 & Nr0nv6));
assign Qexmv6 = (Baxmv6 & U9xmv6);
assign Waxmv6 = (D01nv6 | F11nv6);
assign Kf0nv6 = (~(Y01nv6 & Gr0nv6));
assign W70nv6 = (Dwb7z6[2] & Gr0nv6);
assign Iaxmv6 = (~(C31nv6 | W70nv6));
assign Paxmv6 = (K71nv6 | Iaxmv6);
assign Kbxmv6 = (Waxmv6 & Paxmv6);
assign Dbxmv6 = (~(Hq1et6 & Jw0nv6));
assign Mcxmv6 = (~(Kbxmv6 & Dbxmv6));
assign Ybxmv6 = (~(Mcxmv6 & Dwb7z6[3]));
assign Fhzmv6 = (~(Syzmv6 & R01nv6));
assign Bvxmv6 = (~(Ym0nv6 | A21nv6));
assign Rbxmv6 = (K71nv6 | Bvxmv6);
assign Fcxmv6 = (~(Ybxmv6 & Rbxmv6));
assign Hdxmv6 = (~(Fcxmv6 & Dwb7z6[0]));
assign Tcxmv6 = (~(U51nv6 | Dwb7z6[3]));
assign Adxmv6 = (~(Tcxmv6 & Mcxmv6));
assign Cexmv6 = (Hdxmv6 & Adxmv6);
assign Odxmv6 = (A21nv6 | Apzmv6);
assign Hcymv6 = (~(Odxmv6 & Z41nv6));
assign Vdxmv6 = (D71nv6 | Hcymv6);
assign Jexmv6 = (Cexmv6 & Vdxmv6);
assign Xexmv6 = (~(Qexmv6 & Jexmv6));
assign Wl0nv6 = (~(Dwb7z6[4] | Dwb7z6[5]));
assign Efxmv6 = (~(Xexmv6 & Wl0nv6));
assign Unxmv6 = (Lfxmv6 & Efxmv6);
assign Ufymv6 = (~(Aga7z6 & Hv0nv6));
assign Ov0nv6 = (~(F11nv6 | Z41nv6));
assign Sfxmv6 = (~(Sfydt6 & Ov0nv6));
assign Zfxmv6 = (Ufymv6 & Sfxmv6);
assign Mjxmv6 = (Zfxmv6 & Ynzmv6);
assign Ngxmv6 = (T11nv6 | Kgo7v6);
assign Ggxmv6 = (~(X00et6 & Nr0nv6));
assign Ugxmv6 = (~(Ngxmv6 & Ggxmv6));
assign Phxmv6 = (~(Ugxmv6 & Z41nv6));
assign Bhxmv6 = (~(U51nv6 | Olzdt6));
assign Ihxmv6 = (~(Bhxmv6 & Apzmv6));
assign Yixmv6 = (Phxmv6 & Ihxmv6);
assign Dixmv6 = (E41nv6 | N60nv6);
assign Whxmv6 = (~(Dwb7z6[0] & Nr0nv6));
assign Kixmv6 = (~(Dixmv6 & Whxmv6));
assign Rixmv6 = (~(Kixmv6 & Ys97z6));
assign Fjxmv6 = (Yixmv6 & Rixmv6);
assign Tjxmv6 = (~(Mjxmv6 & Fjxmv6));
assign Av0nv6 = (Dwb7z6[5] & K01nv6);
assign Gnxmv6 = (~(Tjxmv6 & Av0nv6));
assign Qxzmv6 = (~(Dwb7z6[1] | Dwb7z6[2]));
assign R10nv6 = (~(Qxzmv6 | Ci0nv6));
assign Lmxmv6 = (~(Ys97z6 & R10nv6));
assign Akxmv6 = (~(Wxxdt6 & Dwb7z6[1]));
assign Qlxmv6 = (Akxmv6 & Ynzmv6);
assign Hkxmv6 = (~(Dwb7z6[1] | Dwb7z6[0]));
assign Clxmv6 = (~(Hkxmv6 & L32et6));
assign Okxmv6 = (~(M11nv6 | Tnzdt6));
assign Vkxmv6 = (~(Okxmv6 & Dwb7z6[0]));
assign Jlxmv6 = (Clxmv6 & Vkxmv6);
assign Xlxmv6 = (Qlxmv6 & Jlxmv6);
assign Emxmv6 = (Xlxmv6 | R10nv6);
assign Smxmv6 = (~(Lmxmv6 & Emxmv6));
assign Uy0nv6 = (Dwb7z6[5] & Dwb7z6[4]);
assign Zmxmv6 = (~(Smxmv6 & Uy0nv6));
assign Nnxmv6 = (Gnxmv6 & Zmxmv6);
assign Uah7z6[0] = (~(Unxmv6 & Nnxmv6));
assign Ioxmv6 = (~(Ehzdt6 & Jw0nv6));
assign Boxmv6 = (~(Gg0et6 & Hv0nv6));
assign Woxmv6 = (Ioxmv6 & Boxmv6);
assign Ec0nv6 = (Ci0nv6 & Dwb7z6[3]);
assign Poxmv6 = (~(Ec0nv6 & A4zdt6));
assign X6ymv6 = (Q31nv6 & Poxmv6);
assign Csxmv6 = (Woxmv6 & X6ymv6);
assign Dpxmv6 = (Z41nv6 | Btydt6);
assign Ypxmv6 = (~(Dpxmv6 & Fn0nv6));
assign Kpxmv6 = (~(R01nv6 | Tnzdt6));
assign Rpxmv6 = (~(Kpxmv6 & W8zmv6));
assign Orxmv6 = (Ypxmv6 & Rpxmv6);
assign Arxmv6 = (~(Cp0nv6 & Dwb7z6[0]));
assign Fqxmv6 = (R01nv6 | Dwb7z6[2]);
assign Mqxmv6 = (~(J31nv6 & Fqxmv6));
assign Tqxmv6 = (~(Mqxmv6 & Z41nv6));
assign S7ymv6 = (Arxmv6 & Tqxmv6);
assign Hrxmv6 = (S7ymv6 | Iga7z6);
assign Vrxmv6 = (Orxmv6 & Hrxmv6);
assign Jsxmv6 = (~(Csxmv6 & Vrxmv6));
assign Txxmv6 = (~(Jsxmv6 & Ie0nv6));
assign Srzmv6 = (~(Ov0nv6 & Lxydt6));
assign Qsxmv6 = (H21nv6 | Dwb7z6[0]);
assign B2ymv6 = (~(Dwb7z6[3] ^ Z41nv6));
assign Rf0nv6 = (Dwb7z6[2] & O21nv6);
assign Awzmv6 = (~(B2ymv6 & Rf0nv6));
assign Xsxmv6 = (Qsxmv6 & Awzmv6);
assign Erzmv6 = (~(Xsxmv6 & Oa0nv6));
assign Etxmv6 = (~(Gt97z6 & Erzmv6));
assign Stxmv6 = (Srzmv6 & Etxmv6);
assign Ltxmv6 = (~(G12et6 & Nr0nv6));
assign Ywxmv6 = (Stxmv6 & Ltxmv6);
assign Ptzmv6 = (Jw0nv6 & N51nv6);
assign Uuxmv6 = (~(Co1et6 & Ptzmv6));
assign Zkzmv6 = (~(Z41nv6 | Kf0nv6));
assign Ztxmv6 = (Hcymv6 & G51nv6);
assign Acymv6 = (V21nv6 | B2ymv6);
assign Guxmv6 = (~(Ztxmv6 & Acymv6));
assign Nuxmv6 = (~(Kt0et6 & Guxmv6));
assign Kwxmv6 = (Uuxmv6 & Nuxmv6);
assign Wvxmv6 = (~(Dd1et6 & Uszmv6));
assign Ivxmv6 = (~(Bvxmv6 | Z41nv6));
assign Pvxmv6 = (~(Ivxmv6 & E21et6));
assign Dwxmv6 = (Wvxmv6 & Pvxmv6);
assign Rwxmv6 = (Kwxmv6 & Dwxmv6);
assign Fxxmv6 = (~(Ywxmv6 & Rwxmv6));
assign Mxxmv6 = (~(Fxxmv6 & Wl0nv6));
assign V5ymv6 = (Txxmv6 & Mxxmv6);
assign Oyxmv6 = (~(Mdydt6 & Ayxmv6));
assign Tvzmv6 = (~(C31nv6 | A21nv6));
assign Hyxmv6 = (D01nv6 | Tvzmv6);
assign Vyxmv6 = (Oyxmv6 & Hyxmv6);
assign Rm0nv6 = (~(Fhzmv6 | Dwb7z6[0]));
assign N1ymv6 = (Vyxmv6 & S41nv6);
assign Czxmv6 = (Kgo7v6 | Dwb7z6[0]);
assign L0ymv6 = (~(Czxmv6 & Jw0nv6));
assign Jzxmv6 = (R01nv6 & Y01nv6);
assign Qzxmv6 = (~(Jzxmv6 & Syzdt6));
assign Xzxmv6 = (~(H21nv6 & Qzxmv6));
assign E0ymv6 = (~(Xzxmv6 & N51nv6));
assign Z0ymv6 = (L0ymv6 & E0ymv6);
assign Gzzmv6 = (~(N51nv6 | J31nv6));
assign Pgymv6 = (L41nv6 | Gzzmv6);
assign S0ymv6 = (~(Gt97z6 & Pgymv6));
assign G1ymv6 = (Z0ymv6 & S0ymv6);
assign U1ymv6 = (~(N1ymv6 & G1ymv6));
assign H5ymv6 = (~(U1ymv6 & Av0nv6));
assign P2ymv6 = (~(Gt97z6 & R10nv6));
assign I2ymv6 = (B2ymv6 | Kf0nv6);
assign M4ymv6 = (P2ymv6 & I2ymv6);
assign H30nv6 = (Khymv6 & Dwb7z6[0]);
assign Y3ymv6 = (~(Qvxdt6 & H30nv6));
assign D3ymv6 = (D01nv6 | N51nv6);
assign W2ymv6 = (~(G12et6 & N51nv6));
assign K3ymv6 = (~(D3ymv6 & W2ymv6));
assign R3ymv6 = (~(K3ymv6 & Qxzmv6));
assign F4ymv6 = (Y3ymv6 & R3ymv6);
assign T4ymv6 = (~(M4ymv6 & F4ymv6));
assign A5ymv6 = (~(T4ymv6 & Uy0nv6));
assign O5ymv6 = (H5ymv6 & A5ymv6);
assign Uah7z6[1] = (~(V5ymv6 & O5ymv6));
assign Q6ymv6 = (~(Zezdt6 & Jw0nv6));
assign J6ymv6 = (W8zmv6 & D01nv6);
assign Pnymv6 = (~(J6ymv6 & C6ymv6));
assign E7ymv6 = (Q6ymv6 & Pnymv6);
assign W9ymv6 = (E7ymv6 & X6ymv6);
assign L7ymv6 = (~(Be0et6 & Hv0nv6));
assign Wmzmv6 = (~(Ov0nv6 & Cubdt6));
assign I9ymv6 = (L7ymv6 & Wmzmv6);
assign U8ymv6 = (S7ymv6 | Bfo7v6);
assign Jxzmv6 = (~(Lxydt6 | Dwb7z6[0]));
assign Z7ymv6 = (Wqydt6 & Dwb7z6[0]);
assign G8ymv6 = (Jxzmv6 | Z7ymv6);
assign N8ymv6 = (~(G8ymv6 & Fn0nv6));
assign B9ymv6 = (U8ymv6 & N8ymv6);
assign P9ymv6 = (I9ymv6 & B9ymv6);
assign Daymv6 = (~(W9ymv6 & P9ymv6));
assign Gfymv6 = (~(Daymv6 & Ie0nv6));
assign Raymv6 = (~(Bz1et6 & Nr0nv6));
assign Kaymv6 = (~(Ot97z6 & Erzmv6));
assign Yaymv6 = (Raymv6 & Kaymv6);
assign Qczmv6 = (~(Ov0nv6 & D01nv6));
assign Leymv6 = (Yaymv6 & Qczmv6);
assign Mbymv6 = (~(Xl1et6 & Ptzmv6));
assign Fbymv6 = (~(Ya1et6 & Uszmv6));
assign Xdymv6 = (Mbymv6 & Fbymv6);
assign Tbymv6 = (Z41nv6 | Q31nv6);
assign Lsymv6 = (Acymv6 & Tbymv6);
assign Ocymv6 = (~(Lsymv6 & Hcymv6));
assign Jdymv6 = (~(Fr0et6 & Ocymv6));
assign Vcymv6 = (~(Tvzmv6 | Z41nv6));
assign Cdymv6 = (~(Vcymv6 & Nh1et6));
assign Qdymv6 = (Jdymv6 & Cdymv6);
assign Eeymv6 = (Xdymv6 & Qdymv6);
assign Seymv6 = (~(Leymv6 & Eeymv6));
assign Zeymv6 = (~(Seymv6 & Wl0nv6));
assign Nmymv6 = (Gfymv6 & Zeymv6);
assign Hwzmv6 = (~(N51nv6 & Ym0nv6));
assign Igymv6 = (Hwzmv6 & Awzmv6);
assign Nfymv6 = (~(Kf0nv6 | Dwb7z6[0]));
assign Vjymv6 = (~(Nfymv6 & Tnzdt6));
assign Bgymv6 = (Ufymv6 & Vjymv6);
assign Hjymv6 = (Igymv6 & Bgymv6);
assign Dhymv6 = (~(Gbydt6 & Ov0nv6));
assign Wgymv6 = (~(Pgymv6 & Ot97z6));
assign Tiymv6 = (Dhymv6 & Wgymv6);
assign Lyzmv6 = (Khymv6 & N51nv6);
assign Fiymv6 = (~(Nwzdt6 & Lyzmv6));
assign Rhymv6 = (~(Dwb7z6[0] | Tnzdt6));
assign Yhymv6 = (~(Rhymv6 & Apzmv6));
assign Miymv6 = (Fiymv6 & Yhymv6);
assign Ajymv6 = (Tiymv6 & Miymv6);
assign Ojymv6 = (~(Hjymv6 & Ajymv6));
assign Zlymv6 = (~(Ojymv6 & Av0nv6));
assign Ckymv6 = (~(Bz1et6 & Hv0nv6));
assign Elymv6 = (Ckymv6 & Vjymv6);
assign Qkymv6 = (~(Ot97z6 & R10nv6));
assign Jkymv6 = (~(Ktxdt6 & H30nv6));
assign Xkymv6 = (Qkymv6 & Jkymv6);
assign Llymv6 = (~(Elymv6 & Xkymv6));
assign Slymv6 = (~(Llymv6 & Uy0nv6));
assign Gmymv6 = (Zlymv6 & Slymv6);
assign Uah7z6[2] = (~(Nmymv6 & Gmymv6));
assign Inymv6 = (~(Wb0et6 & Hv0nv6));
assign Bnymv6 = (Q31nv6 | Aga7z6);
assign Umymv6 = (~(R71nv6 & Ov0nv6));
assign Bfzmv6 = (Bnymv6 & Umymv6);
assign Wnymv6 = (Inymv6 & Bfzmv6);
assign Oqymv6 = (Wnymv6 & Pnymv6);
assign Koymv6 = (~(V1zdt6 & Zkzmv6));
assign Fazmv6 = (Syzmv6 & X31nv6);
assign B8zmv6 = (~(Fazmv6 & Z41nv6));
assign Doymv6 = (B8zmv6 | Aga7z6);
assign Aqymv6 = (Koymv6 & Doymv6);
assign Roymv6 = (Rf0nv6 & X31nv6);
assign Mpymv6 = (~(Roymv6 & Uczdt6));
assign Yoymv6 = (Fazmv6 & Dwb7z6[0]);
assign Fpymv6 = (~(Yoymv6 & Qoydt6));
assign Tpymv6 = (Mpymv6 & Fpymv6);
assign Hqymv6 = (Aqymv6 & Tpymv6);
assign Vqymv6 = (~(Oqymv6 & Hqymv6));
assign Rvymv6 = (~(Vqymv6 & Ie0nv6));
assign Jrymv6 = (~(Ww1et6 & Nr0nv6));
assign Crymv6 = (~(Qs97z6 & Erzmv6));
assign Qrymv6 = (Jrymv6 & Crymv6);
assign Wuymv6 = (Qrymv6 & Qczmv6);
assign Esymv6 = (~(Wb0et6 & Ptzmv6));
assign Xrymv6 = (~(Sj1et6 & Rm0nv6));
assign Iuymv6 = (Esymv6 & Xrymv6);
assign Utymv6 = (~(T81et6 & Uszmv6));
assign Ssymv6 = (~(Apzmv6 & Z41nv6));
assign Zsymv6 = (Ssymv6 & Lsymv6);
assign J5zmv6 = (Zsymv6 & G51nv6);
assign Knzmv6 = (Fhzmv6 | Z41nv6);
assign Gtymv6 = (~(J5zmv6 & Knzmv6));
assign Ntymv6 = (~(Ap0et6 & Gtymv6));
assign Buymv6 = (Utymv6 & Ntymv6);
assign Puymv6 = (Iuymv6 & Buymv6);
assign Dvymv6 = (~(Wuymv6 & Puymv6));
assign Kvymv6 = (~(Dvymv6 & Wl0nv6));
assign A4zmv6 = (Rvymv6 & Kvymv6);
assign U7zmv6 = (~(Hv0nv6 & Lxydt6));
assign Yvymv6 = (~(N60nv6 & Gr0nv6));
assign Fwymv6 = (U7zmv6 & Yvymv6);
assign N0zmv6 = (Fwymv6 & Hwzmv6);
assign Cyymv6 = (~(Qs97z6 & Gzzmv6));
assign Twymv6 = (Fhzmv6 | Tnzdt6);
assign Mwymv6 = (~(A9ydt6 & Qxzmv6));
assign Hxymv6 = (Twymv6 & Mwymv6);
assign Axymv6 = (~(Qs97z6 & Fn0nv6));
assign Oxymv6 = (~(Hxymv6 & Axymv6));
assign Vxymv6 = (~(Oxymv6 & Dwb7z6[0]));
assign Zzymv6 = (Cyymv6 & Vxymv6);
assign Lzymv6 = (~(Iuzdt6 & Lyzmv6));
assign Qyymv6 = (Dwb7z6[1] | Yga7z6);
assign Jyymv6 = (~(Olzdt6 & Dwb7z6[3]));
assign Xyymv6 = (~(Qyymv6 & Jyymv6));
assign Ezymv6 = (~(Xyymv6 & W8zmv6));
assign Szymv6 = (Lzymv6 & Ezymv6);
assign G0zmv6 = (Zzymv6 & Szymv6);
assign U0zmv6 = (~(N0zmv6 & G0zmv6));
assign M3zmv6 = (~(U0zmv6 & Av0nv6));
assign B1zmv6 = (~(Ww1et6 & Hv0nv6));
assign R2zmv6 = (B1zmv6 & G51nv6);
assign P1zmv6 = (~(Erxdt6 & H30nv6));
assign F20nv6 = (Qxzmv6 & Dwb7z6[0]);
assign I1zmv6 = (~(F20nv6 & D01nv6));
assign D2zmv6 = (P1zmv6 & I1zmv6);
assign W1zmv6 = (~(Qs97z6 & R10nv6));
assign K2zmv6 = (D2zmv6 & W1zmv6);
assign Y2zmv6 = (~(R2zmv6 & K2zmv6));
assign F3zmv6 = (~(Y2zmv6 & Uy0nv6));
assign T3zmv6 = (M3zmv6 & F3zmv6);
assign Uah7z6[3] = (~(A4zmv6 & T3zmv6));
assign O4zmv6 = (~(Aga7z6 & Ov0nv6));
assign H4zmv6 = (~(Is97z6 & Erzmv6));
assign C5zmv6 = (O4zmv6 & H4zmv6);
assign V4zmv6 = (~(Ru1et6 & Nr0nv6));
assign Z6zmv6 = (C5zmv6 & V4zmv6);
assign Nszmv6 = (~(Fhzmv6 & J5zmv6));
assign X5zmv6 = (~(Vm0et6 & Nszmv6));
assign Q5zmv6 = (~(O61et6 & Uszmv6));
assign L6zmv6 = (X5zmv6 & Q5zmv6);
assign E6zmv6 = (~(R90et6 & Ptzmv6));
assign S6zmv6 = (L6zmv6 & E6zmv6);
assign G7zmv6 = (~(Z6zmv6 & S6zmv6));
assign Jczmv6 = (~(G7zmv6 & Wl0nv6));
assign N7zmv6 = (~(U6ydt6 & Ov0nv6));
assign I8zmv6 = (U7zmv6 & N7zmv6);
assign Obzmv6 = (I8zmv6 & B8zmv6);
assign P8zmv6 = (N51nv6 & Nr0nv6);
assign Y9zmv6 = (~(P8zmv6 & Dszdt6));
assign K9zmv6 = (W8zmv6 & X31nv6);
assign D9zmv6 = (~(Dwb7z6[1] | Kgo7v6));
assign R9zmv6 = (~(K9zmv6 & D9zmv6));
assign Abzmv6 = (Y9zmv6 & R9zmv6);
assign Mazmv6 = (Gzzmv6 | Fazmv6);
assign Tazmv6 = (~(Mazmv6 & Is97z6));
assign Hbzmv6 = (Abzmv6 & Tazmv6);
assign Vbzmv6 = (~(Obzmv6 & Hbzmv6));
assign Cczmv6 = (~(Vbzmv6 & Av0nv6));
assign Skzmv6 = (Jczmv6 & Cczmv6);
assign Xczmv6 = (~(Ru1et6 & Hv0nv6));
assign Nezmv6 = (Xczmv6 & Qczmv6);
assign Zdzmv6 = (~(Yoxdt6 & H30nv6));
assign Edzmv6 = (J31nv6 | Dwb7z6[0]);
assign Ldzmv6 = (~(Y01nv6 & Edzmv6));
assign Sdzmv6 = (~(Ldzmv6 & Is97z6));
assign Gezmv6 = (Zdzmv6 & Sdzmv6);
assign Uezmv6 = (~(Nezmv6 & Gezmv6));
assign Ekzmv6 = (~(Uezmv6 & Uy0nv6));
assign Dgzmv6 = (S41nv6 & Bfzmv6);
assign Pfzmv6 = (~(Pazdt6 & Jw0nv6));
assign Ifzmv6 = (~(R90et6 & Hv0nv6));
assign Wfzmv6 = (Pfzmv6 & Ifzmv6);
assign Jjzmv6 = (Dgzmv6 & Wfzmv6);
assign Rgzmv6 = (~(Kmydt6 & L41nv6));
assign Kgzmv6 = (D01nv6 | V21nv6);
assign Vizmv6 = (Rgzmv6 & Kgzmv6);
assign Ygzmv6 = (Kf0nv6 | Dwb7z6[0]);
assign Mhzmv6 = (~(Fhzmv6 & Ygzmv6));
assign Hizmv6 = (~(Bfo7v6 & Mhzmv6));
assign Thzmv6 = (~(Dwb7z6[0] | Aga7z6));
assign Aizmv6 = (~(Thzmv6 & Syzmv6));
assign Oizmv6 = (Hizmv6 & Aizmv6);
assign Cjzmv6 = (Vizmv6 & Oizmv6);
assign Qjzmv6 = (~(Jjzmv6 & Cjzmv6));
assign Xjzmv6 = (~(Qjzmv6 & Ie0nv6));
assign Lkzmv6 = (Ekzmv6 & Xjzmv6);
assign Uah7z6[4] = (~(Skzmv6 & Lkzmv6));
assign Pmzmv6 = (~(Nr0nv6 | Zkzmv6));
assign Nlzmv6 = (~(K8zdt6 & Jw0nv6));
assign Glzmv6 = (~(M70et6 & Hv0nv6));
assign Bmzmv6 = (Nlzmv6 & Glzmv6);
assign Ulzmv6 = (Lxydt6 | J31nv6);
assign Imzmv6 = (Bmzmv6 & Ulzmv6);
assign Qqzmv6 = (Pmzmv6 & Imzmv6);
assign Dnzmv6 = (~(Ekydt6 & L41nv6));
assign Cqzmv6 = (Dnzmv6 & Wmzmv6);
assign Rnzmv6 = (~(Kf0nv6 & Knzmv6));
assign Tozmv6 = (~(Rnzmv6 & Iga7z6));
assign Fozmv6 = (~(Ynzmv6 | Tnzdt6));
assign Mozmv6 = (~(Fozmv6 & Dwb7z6[2]));
assign Opzmv6 = (Tozmv6 & Mozmv6);
assign Hpzmv6 = (~(Jxzmv6 & Apzmv6));
assign Vpzmv6 = (Opzmv6 & Hpzmv6);
assign Jqzmv6 = (Cqzmv6 & Vpzmv6);
assign Xqzmv6 = (~(Qqzmv6 & Jqzmv6));
assign Mvzmv6 = (~(Xqzmv6 & Ie0nv6));
assign Lrzmv6 = (~(Y4a7z6 & Erzmv6));
assign Gszmv6 = (Srzmv6 & Lrzmv6);
assign Zrzmv6 = (~(Ms1et6 & Nr0nv6));
assign Ruzmv6 = (Gszmv6 & Zrzmv6);
assign Itzmv6 = (~(Qk0et6 & Nszmv6));
assign Btzmv6 = (~(J41et6 & Uszmv6));
assign Duzmv6 = (Itzmv6 & Btzmv6);
assign Wtzmv6 = (~(Ptzmv6 & M70et6));
assign Kuzmv6 = (Duzmv6 & Wtzmv6);
assign Yuzmv6 = (~(Ruzmv6 & Kuzmv6));
assign Fvzmv6 = (~(Yuzmv6 & Wl0nv6));
assign S50nv6 = (Mvzmv6 & Fvzmv6);
assign Cxzmv6 = (Awzmv6 & Tvzmv6);
assign Owzmv6 = (~(Yga7z6 & Jw0nv6));
assign Vwzmv6 = (Owzmv6 & Hwzmv6);
assign D10nv6 = (Cxzmv6 & Vwzmv6);
assign Eyzmv6 = (~(Qxzmv6 & Jxzmv6));
assign Xxzmv6 = (~(O4ydt6 & F20nv6));
assign P00nv6 = (Eyzmv6 & Xxzmv6);
assign B00nv6 = (~(Ypzdt6 & Lyzmv6));
assign Zyzmv6 = (Syzmv6 & Dwb7z6[0]);
assign Nzzmv6 = (Gzzmv6 | Zyzmv6);
assign Uzzmv6 = (~(Nzzmv6 & Y4a7z6));
assign I00nv6 = (B00nv6 & Uzzmv6);
assign W00nv6 = (P00nv6 & I00nv6);
assign K10nv6 = (~(D10nv6 & W00nv6));
assign E50nv6 = (~(K10nv6 & Av0nv6));
assign Y10nv6 = (~(Y4a7z6 & R10nv6));
assign J40nv6 = (Y10nv6 & Kf0nv6);
assign A30nv6 = (~(Tnzdt6 & F20nv6));
assign M20nv6 = (~(H21nv6 | Dwb7z6[0]));
assign T20nv6 = (~(M20nv6 & Ms1et6));
assign V30nv6 = (A30nv6 & T20nv6);
assign O30nv6 = (~(Smxdt6 & H30nv6));
assign C40nv6 = (V30nv6 & O30nv6);
assign Q40nv6 = (~(J40nv6 & C40nv6));
assign X40nv6 = (~(Q40nv6 & Uy0nv6));
assign L50nv6 = (E50nv6 & X40nv6);
assign Uah7z6[5] = (~(S50nv6 & L50nv6));
assign I70nv6 = (~(Ea2et6 & U51nv6));
assign G60nv6 = (~(Jc2et6 & Dwb7z6[0]));
assign Z50nv6 = (~(Gr2et6 & Z41nv6));
assign U60nv6 = (~(G60nv6 & Z50nv6));
assign B70nv6 = (~(U60nv6 & N60nv6));
assign P70nv6 = (~(I70nv6 & B70nv6));
assign K80nv6 = (~(Cp0nv6 & P70nv6));
assign D80nv6 = (~(W70nv6 & Gr2et6));
assign T90nv6 = (K80nv6 & D80nv6);
assign Y80nv6 = (W61nv6 | Y01nv6);
assign R80nv6 = (~(H50et6 & Y01nv6));
assign F90nv6 = (Y80nv6 & R80nv6);
assign Aa0nv6 = (F90nv6 & Dwb7z6[0]);
assign M90nv6 = (F11nv6 | Aa0nv6);
assign Ud0nv6 = (T90nv6 & M90nv6);
assign Ha0nv6 = (Aa0nv6 | M11nv6);
assign Va0nv6 = (~(Oa0nv6 & Ha0nv6));
assign Qb0nv6 = (~(Va0nv6 & O5a7z6));
assign Cb0nv6 = (Jc2et6 | Dwb7z6[2]);
assign Jb0nv6 = (~(Cb0nv6 & I61nv6));
assign Gd0nv6 = (Qb0nv6 & Jb0nv6);
assign Xb0nv6 = (Fn0nv6 & Z41nv6);
assign Sc0nv6 = (~(Xb0nv6 & Z72et6));
assign Lc0nv6 = (~(Ec0nv6 & Po2et6));
assign Zc0nv6 = (Sc0nv6 & Lc0nv6);
assign Nd0nv6 = (Gd0nv6 & Zc0nv6);
assign Be0nv6 = (~(Ud0nv6 & Nd0nv6));
assign Km0nv6 = (~(Ie0nv6 & Be0nv6));
assign We0nv6 = (~(Cp0nv6 & Po2et6));
assign Pe0nv6 = (~(Ov0nv6 & Z72et6));
assign Df0nv6 = (We0nv6 & Pe0nv6);
assign Il0nv6 = (Df0nv6 & G51nv6);
assign Vh0nv6 = (~(O5a7z6 | Z41nv6));
assign Oh0nv6 = (T11nv6 | Vh0nv6);
assign Fg0nv6 = (W61nv6 | Kf0nv6);
assign Yf0nv6 = (~(Zz0et6 & Rf0nv6));
assign Tg0nv6 = (Fg0nv6 & Yf0nv6);
assign Mg0nv6 = (~(Nj2et6 & Xw0nv6));
assign Ah0nv6 = (~(Tg0nv6 & Mg0nv6));
assign Hh0nv6 = (~(Ah0nv6 & Z41nv6));
assign Uk0nv6 = (Oh0nv6 & Hh0nv6);
assign Qi0nv6 = (Y01nv6 | P61nv6);
assign Ji0nv6 = (B61nv6 | Po2et6);
assign Lj0nv6 = (Qi0nv6 & Ji0nv6);
assign Xi0nv6 = (E41nv6 | W61nv6);
assign Ej0nv6 = (~(Q31nv6 & Xi0nv6));
assign Gk0nv6 = (~(Lj0nv6 & Ej0nv6));
assign Zj0nv6 = (~(Sj0nv6 & Gr2et6));
assign Nk0nv6 = (Gk0nv6 & Zj0nv6);
assign Bl0nv6 = (Uk0nv6 & Nk0nv6);
assign Pl0nv6 = (~(Il0nv6 & Bl0nv6));
assign Dm0nv6 = (~(Wl0nv6 & Pl0nv6));
assign Wz0nv6 = (Km0nv6 & Dm0nv6);
assign Ho0nv6 = (~(Ym0nv6 | Rm0nv6));
assign Tn0nv6 = (~(Fn0nv6 & Po2et6));
assign Mn0nv6 = (~(Qzydt6 & Hv0nv6));
assign Ao0nv6 = (Tn0nv6 & Mn0nv6);
assign Mu0nv6 = (Ho0nv6 & Ao0nv6);
assign Vo0nv6 = (~(C0ydt6 & A21nv6));
assign Oo0nv6 = (~(Yhydt6 & Ov0nv6));
assign Yt0nv6 = (Vo0nv6 & Oo0nv6);
assign Qp0nv6 = (~(F6zdt6 & Jw0nv6));
assign Jp0nv6 = (~(C30et6 & Cp0nv6));
assign Xp0nv6 = (~(Qp0nv6 & Jp0nv6));
assign Sq0nv6 = (~(Xp0nv6 & Z41nv6));
assign Eq0nv6 = (Gr2et6 | Y01nv6);
assign Lq0nv6 = (~(Eq0nv6 & I61nv6));
assign Kt0nv6 = (Sq0nv6 & Lq0nv6);
assign Zq0nv6 = (~(I2ydt6 & Jw0nv6));
assign Ps0nv6 = (Zq0nv6 & E41nv6);
assign Bs0nv6 = (~(O5a7z6 & Gr0nv6));
assign Ur0nv6 = (~(Hbo7v6 & Nr0nv6));
assign Is0nv6 = (Bs0nv6 & Ur0nv6);
assign Ws0nv6 = (~(Ps0nv6 & Is0nv6));
assign Dt0nv6 = (~(Ws0nv6 & Dwb7z6[0]));
assign Rt0nv6 = (Kt0nv6 & Dt0nv6);
assign Fu0nv6 = (Yt0nv6 & Rt0nv6);
assign Tu0nv6 = (~(Mu0nv6 & Fu0nv6));
assign Iz0nv6 = (~(Av0nv6 & Tu0nv6));
assign Cw0nv6 = (~(Hv0nv6 & Po2et6));
assign Vv0nv6 = (~(Mkxdt6 & Ov0nv6));
assign Gy0nv6 = (Cw0nv6 & Vv0nv6);
assign Qw0nv6 = (Dwb7z6[2] | Jw0nv6);
assign Sx0nv6 = (~(Qw0nv6 & Gr2et6));
assign Ex0nv6 = (~(Xw0nv6 | Dwb7z6[2]));
assign Lx0nv6 = (~(Ex0nv6 & P61nv6));
assign Zx0nv6 = (Sx0nv6 & Lx0nv6);
assign Ny0nv6 = (~(Gy0nv6 & Zx0nv6));
assign Bz0nv6 = (~(Uy0nv6 & Ny0nv6));
assign Pz0nv6 = (Iz0nv6 & Bz0nv6);
assign Q52et6 = (~(Wz0nv6 & Pz0nv6));
assign D01nv6 = (!Tnzdt6);
assign K01nv6 = (!Dwb7z6[4]);
assign R01nv6 = (!Dwb7z6[3]);
assign Y01nv6 = (!Dwb7z6[2]);
assign F11nv6 = (!Ayxmv6);
assign M11nv6 = (!Xw0nv6);
assign T11nv6 = (!Jw0nv6);
assign A21nv6 = (!Fhzmv6);
assign H21nv6 = (!Qxzmv6);
assign O21nv6 = (!Dwb7z6[1]);
assign V21nv6 = (!W70nv6);
assign C31nv6 = (!Kf0nv6);
assign J31nv6 = (!Khymv6);
assign Q31nv6 = (!Ym0nv6);
assign X31nv6 = (!C6ymv6);
assign E41nv6 = (!Fn0nv6);
assign L41nv6 = (!Oa0nv6);
assign S41nv6 = (!Rm0nv6);
assign Z41nv6 = (!Dwb7z6[0]);
assign G51nv6 = (!Zkzmv6);
assign N51nv6 = (!B2ymv6);
assign U51nv6 = (!N60nv6);
assign B61nv6 = (!Ci0nv6);
assign I61nv6 = (!Ynzmv6);
assign P61nv6 = (!Vh0nv6);
assign W61nv6 = (!O5a7z6);
assign D71nv6 = (!Pv0et6);
assign K71nv6 = (!Ux0et6);
assign R71nv6 = (!Cubdt6);
assign Zpe7v6 = (~(Y71nv6 & F81nv6));
assign F81nv6 = (~(M81nv6 & T81nv6));
assign Y71nv6 = (A91nv6 & H91nv6);
assign A91nv6 = (~(Xre7v6 & O91nv6));
assign O91nv6 = (~(V91nv6 & Ca1nv6));
assign Rte7v6 = (L9e7v6 | Ja1nv6);
assign Ja1nv6 = (I6e7v6 & H91nv6);
assign H91nv6 = (~(Qa1nv6 & Xa1nv6));
assign Xa1nv6 = (Eb1nv6 ? T81nv6 : V91nv6);
assign Qa1nv6 = (Lb1nv6 & I6e7v6);
assign Ame7v6 = (~(Y097z6 & Sb1nv6));
assign Sb1nv6 = (~(Xzd7v6 & Lkh7v6));
assign Boe7v6 = (~(Zb1nv6 & Gc1nv6));
assign Gc1nv6 = (~(G1e7v6 & Ekh7v6));
assign Mq47v6 = (~(Nc1nv6 & SWDITMS));
assign Qr47v6 = (~(Uc1nv6 & SWDITMS));
assign Us47v6 = (Uia7z6 & SWDITMS);
assign Jv47v6 = (~(Bd1nv6 & Id1nv6));
assign Id1nv6 = (~(Pd1nv6 & Wd1nv6));
assign Pd1nv6 = (~(De1nv6 & Ke1nv6));
assign Bd1nv6 = (~(Re1nv6 | Ye1nv6));
assign Vw47v6 = (~(Ff1nv6 & Mf1nv6));
assign Mf1nv6 = (Tf1nv6 & Ag1nv6);
assign Ag1nv6 = (~(Uj57v6 & Ye1nv6));
assign Ye1nv6 = (Hg1nv6 & Uzxmz6[4]);
assign Hg1nv6 = (Uzxmz6[1] & Og1nv6);
assign Tf1nv6 = (Vg1nv6 & Ch1nv6);
assign Ch1nv6 = (~(Jh1nv6 & Qh1nv6));
assign Jh1nv6 = (Hf57v6 ? Ei1nv6 : Xh1nv6);
assign Vg1nv6 = (~(Cxxmz6[0] & Re1nv6));
assign Re1nv6 = (Li1nv6 & Uzxmz6[0]);
assign Ff1nv6 = (Si1nv6 & Zi1nv6);
assign Zi1nv6 = (Ke1nv6 | Gj1nv6);
assign Si1nv6 = (De1nv6 ? Nj1nv6 : Wd1nv6);
assign De1nv6 = (~(Xh1nv6 | Ei1nv6));
assign Nj1nv6 = (~(Uj1nv6 & Ke1nv6));
assign Lt57v6 = (Bk1nv6 | Ik1nv6);
assign Ik1nv6 = (R9ymz6[3] ? G8ymz6[0] : Pk1nv6);
assign Pk1nv6 = (Wk1nv6 & Dl1nv6);
assign Dl1nv6 = (Kl1nv6 | L5ymz6[34]);
assign Kl1nv6 = (Rl1nv6 & W6ymz6[3]);
assign Rl1nv6 = (Yl1nv6 & Fm1nv6);
assign Fm1nv6 = (Mm1nv6 | Tm1nv6);
assign Yl1nv6 = (~(W6ymz6[0] & An1nv6));
assign Wk1nv6 = (Hn1nv6 & On1nv6);
assign On1nv6 = (~(Vn1nv6 & Co1nv6));
assign Vn1nv6 = (Jo1nv6 & Qo1nv6);
assign Hn1nv6 = (~(Xo1nv6 & Ep1nv6));
assign Ep1nv6 = (Mm1nv6 ? Qo1nv6 : Lp1nv6);
assign Lp1nv6 = (~(W6ymz6[0] | L5ymz6[3]));
assign Xo1nv6 = (W6ymz6[1] & W6ymz6[3]);
assign Bk1nv6 = (~(Sp1nv6 & Zp1nv6));
assign Sp1nv6 = (Gq1nv6 ^ Nq1nv6);
assign Z3ymz6[3] = (~(Uq1nv6 & Br1nv6));
assign Br1nv6 = (Ir1nv6 & Pr1nv6);
assign Ir1nv6 = (~(Wr1nv6 & Ds1nv6));
assign Uq1nv6 = (Ks1nv6 & Rs1nv6);
assign Rs1nv6 = (~(Ys1nv6 & Gq1nv6));
assign Ys1nv6 = (!Ft1nv6);
assign Ks1nv6 = (~(R9ymz6[3] & Zp1nv6));
assign Z3ymz6[2] = (~(Mt1nv6 & Tt1nv6));
assign Tt1nv6 = (~(R9ymz6[2] & Au1nv6));
assign Au1nv6 = (~(R9ymz6[1] & Nq1nv6));
assign Mt1nv6 = (~(Hu1nv6 & Gq1nv6));
assign Z3ymz6[1] = (Ou1nv6 | Vu1nv6);
assign Ou1nv6 = (Wr1nv6 ? Cv1nv6 : Ds1nv6);
assign Cv1nv6 = (~(Jv1nv6 & Qv1nv6));
assign Jv1nv6 = (Xv1nv6 & Ew1nv6);
assign Ew1nv6 = (Lw1nv6 | R9ymz6[3]);
assign Xv1nv6 = (Pr1nv6 | R9ymz6[0]);
assign Ds1nv6 = (R9ymz6[2] & Gq1nv6);
assign Z3ymz6[0] = (Vu1nv6 | Sw1nv6);
assign Sw1nv6 = (Zw1nv6 & Hu1nv6);
assign Hu1nv6 = (!Wr1nv6);
assign Zw1nv6 = (~(Gx1nv6 & Qv1nv6));
assign Qv1nv6 = (~(Nx1nv6 | Ux1nv6));
assign Ux1nv6 = (~(R9ymz6[1] | R9ymz6[2]));
assign Gx1nv6 = (~(Nq1nv6 | By1nv6));
assign Vu1nv6 = (Wr1nv6 ? Py1nv6 : Iy1nv6);
assign Wr1nv6 = (JTAGNSW & K3a7z6);
assign Py1nv6 = (R9ymz6[0] & Zp1nv6);
assign Oa67v6 = (Dz1nv6 ? Wy1nv6 : Esf8v6);
assign G967v6 = (JTAGNSW ? Rz1nv6 : Kz1nv6);
assign Rz1nv6 = (Hw57v6 & Esf8v6);
assign Kz1nv6 = (Uz47v6 & Wy1nv6);
assign O667v6 = (Dz1nv6 ? Sl47v6 : Mg47v6);
assign X767v6 = (Dz1nv6 ? Qm47v6 : Kh47v6);
assign Ddeet6 = (~(Yz1nv6 | Ffeet6));
assign Yz1nv6 = (Dgo7v6 & F02nv6);
assign X8eet6 = (M02nv6 & T02nv6);
assign T02nv6 = (Dgo7v6 ? Cbeet6 : Ffeet6);
assign M02nv6 = (A12nv6 & F02nv6);
assign T9fet6 = (H12nv6 & O12nv6);
assign O12nv6 = (V12nv6 & C22nv6);
assign C22nv6 = (J22nv6 & Q22nv6);
assign J22nv6 = (X22nv6 & E32nv6);
assign H12nv6 = (L32nv6 & S32nv6);
assign S32nv6 = (Z32nv6 & G42nv6);
assign L32nv6 = (Toi7z6[9] & N42nv6);
assign Hbfet6 = (Q22nv6 & U42nv6);
assign Vcfet6 = (Q22nv6 & B52nv6);
assign Jefet6 = (Q22nv6 & I52nv6);
assign Xffet6 = (Q22nv6 & P52nv6);
assign Lhfet6 = (Q22nv6 & W52nv6);
assign Zifet6 = (Q22nv6 & D62nv6);
assign Nkfet6 = (Q22nv6 & K62nv6);
assign Bmfet6 = (Q22nv6 & R62nv6);
assign P3m8v6 = (Sja7z6 & Kja7z6);
assign Gpfet6 = (Y62nv6 & F72nv6);
assign F72nv6 = (M72nv6 & T72nv6);
assign T72nv6 = (~(A82nv6 & H82nv6));
assign H82nv6 = (O82nv6 & V82nv6);
assign O82nv6 = (~(C92nv6 & J92nv6));
assign A82nv6 = (Nmadt6 & Q92nv6);
assign Q92nv6 = (~(Fjadt6 & Inadt6));
assign M72nv6 = (~(Ovfet6 | Qtfet6));
assign Y62nv6 = (X92nv6 & D5cet6);
assign X92nv6 = (Ea2nv6 & La2nv6);
assign La2nv6 = (~(Sa2nv6 & Za2nv6));
assign Ozfet6 = (~(Gb2nv6 & Nb2nv6));
assign Nb2nv6 = (~(Ub2nv6 & Bc2nv6));
assign Gb2nv6 = (~(Ic2nv6 & Pc2nv6));
assign Pc2nv6 = (Wc2nv6 & Dd2nv6);
assign Dd2nv6 = (~(Kd2nv6 & Rd2nv6));
assign Wc2nv6 = (~(Yd2nv6 | Fe2nv6));
assign Ic2nv6 = (Me2nv6 & E1cet6);
assign Me2nv6 = (Te2nv6 & Nmadt6);
assign Qtfet6 = (Af2nv6 & Hf2nv6);
assign Hf2nv6 = (Of2nv6 & Vf2nv6);
assign Vf2nv6 = (Cg2nv6 & Jg2nv6);
assign Cg2nv6 = (Qg2nv6 & Xg2nv6);
assign Of2nv6 = (Eh2nv6 & Lh2nv6);
assign Eh2nv6 = (Sh2nv6 & SLEEPHOLDACKn);
assign Af2nv6 = (Zh2nv6 & Gi2nv6);
assign Gi2nv6 = (Ni2nv6 & Ui2nv6);
assign Ni2nv6 = (Za2nv6 & Bj2nv6);
assign Zh2nv6 = (Ij2nv6 & Ub2nv6);
assign Ij2nv6 = (Pj2nv6 & Wj2nv6);
assign Wj2nv6 = (~(Dk2nv6 & Kk2nv6));
assign Kk2nv6 = (Rk2nv6 & Yk2nv6);
assign Yk2nv6 = (Fl2nv6 & Ml2nv6);
assign Ml2nv6 = (Tl2nv6 & Am2nv6);
assign Am2nv6 = (Hm2nv6 & Om2nv6);
assign Hm2nv6 = (Vm2nv6 & Cn2nv6);
assign Tl2nv6 = (Jn2nv6 & Qn2nv6);
assign Jn2nv6 = (~(Z3j7z6[11] | Z3j7z6[3]));
assign Fl2nv6 = (Xn2nv6 & Eo2nv6);
assign Eo2nv6 = (Lo2nv6 & So2nv6);
assign Lo2nv6 = (Zo2nv6 & Gp2nv6);
assign Xn2nv6 = (Np2nv6 & Up2nv6);
assign Np2nv6 = (Bq2nv6 & Iq2nv6);
assign Rk2nv6 = (Pq2nv6 & Wq2nv6);
assign Wq2nv6 = (Dr2nv6 & Kr2nv6);
assign Kr2nv6 = (Rr2nv6 & Yr2nv6);
assign Rr2nv6 = (Fs2nv6 & Ms2nv6);
assign Dr2nv6 = (~(Ts2nv6 | G5j7z6[18]));
assign Ts2nv6 = (G5j7z6[19] | G5j7z6[48]);
assign Pq2nv6 = (At2nv6 & Ht2nv6);
assign Ht2nv6 = (Ot2nv6 & Vt2nv6);
assign Ot2nv6 = (Cu2nv6 & Ju2nv6);
assign At2nv6 = (Qu2nv6 & Xu2nv6);
assign Qu2nv6 = (Ev2nv6 & Lv2nv6);
assign Dk2nv6 = (Sv2nv6 & Zv2nv6);
assign Zv2nv6 = (Gw2nv6 & Nw2nv6);
assign Nw2nv6 = (Uw2nv6 & Bx2nv6);
assign Bx2nv6 = (Ix2nv6 & Px2nv6);
assign Ix2nv6 = (~(Wx2nv6 | Dy2nv6));
assign Uw2nv6 = (Ky2nv6 & Ry2nv6);
assign Ky2nv6 = (~(Yy2nv6 | Fz2nv6));
assign Gw2nv6 = (Mz2nv6 & Tz2nv6);
assign Tz2nv6 = (A03nv6 & H03nv6);
assign A03nv6 = (~(O03nv6 | V03nv6));
assign Mz2nv6 = (C13nv6 & J13nv6);
assign C13nv6 = (Q13nv6 & X13nv6);
assign Sv2nv6 = (E23nv6 & L23nv6);
assign L23nv6 = (S23nv6 & Z23nv6);
assign Z23nv6 = (G33nv6 & N33nv6);
assign G33nv6 = (U33nv6 & B43nv6);
assign S23nv6 = (I43nv6 & P43nv6);
assign I43nv6 = (W43nv6 & D53nv6);
assign E23nv6 = (K53nv6 & R53nv6);
assign R53nv6 = (Y53nv6 & F63nv6);
assign Y53nv6 = (~(M63nv6 | T63nv6));
assign K53nv6 = (A73nv6 & H73nv6);
assign A73nv6 = (O73nv6 & V73nv6);
assign S1get6 = (Ea2nv6 & Za2nv6);
assign Lrfet6 = (~(C83nv6 & J83nv6));
assign J83nv6 = (~(Q83nv6 & X83nv6));
assign Q83nv6 = (E93nv6 & L93nv6);
assign E93nv6 = (~(S93nv6 & Z93nv6));
assign Z93nv6 = (~(Ga3nv6 & Qg2nv6));
assign C83nv6 = (~(Na3nv6 & Tnzdt6));
assign Ovfet6 = (Ua3nv6 & Pj2nv6);
assign Pj2nv6 = (~(Sa2nv6 & S93nv6));
assign Ua3nv6 = (L93nv6 & Bb3nv6);
assign Bb3nv6 = (!Ib3nv6);
assign L93nv6 = (~(Pb3nv6 & Oreet6));
assign Pb3nv6 = (Wb3nv6 & S93nv6);
assign Wb3nv6 = (~(Dc3nv6 & Kc3nv6));
assign Kc3nv6 = (~(Rc3nv6 & P2j7z6[1]));
assign Pnmet6 = (~(Yc3nv6 & Fd3nv6));
assign Fd3nv6 = (Md3nv6 & Td3nv6);
assign Td3nv6 = (Oe3nv6 ? He3nv6 : Ae3nv6);
assign He3nv6 = (~(HADDRI[28] & Ve3nv6));
assign Ae3nv6 = (~(Cf3nv6 & HADDRI[25]));
assign Cf3nv6 = (!Jf3nv6);
assign Md3nv6 = (Qf3nv6 & Xf3nv6);
assign Xf3nv6 = (Ve3nv6 | Eg3nv6);
assign Qf3nv6 = (Zg3nv6 ? Sg3nv6 : Lg3nv6);
assign Sg3nv6 = (~(Gh3nv6 & HADDRI[19]));
assign Lg3nv6 = (~(HADDRI[22] & Jf3nv6));
assign Yc3nv6 = (Nh3nv6 & Uh3nv6);
assign Uh3nv6 = (Pi3nv6 ? Ii3nv6 : Bi3nv6);
assign Ii3nv6 = (~(HADDRI[10] & Wi3nv6));
assign Bi3nv6 = (Dj3nv6 | Kj3nv6);
assign Nh3nv6 = (Fk3nv6 ? Yj3nv6 : Rj3nv6);
assign Yj3nv6 = (~(HADDRI[16] & Mk3nv6));
assign Rj3nv6 = (~(Tk3nv6 & HADDRI[13]));
assign Crmet6 = (~(Al3nv6 & Hl3nv6));
assign Hl3nv6 = (Ol3nv6 & Vl3nv6);
assign Vl3nv6 = (Qm3nv6 ? Jm3nv6 : Cm3nv6);
assign Jm3nv6 = (~(Xm3nv6 & HADDRI[24]));
assign Cm3nv6 = (~(HADDRI[27] & En3nv6));
assign Ol3nv6 = (Ln3nv6 & Sn3nv6);
assign Sn3nv6 = (Zn3nv6 | En3nv6);
assign Ln3nv6 = (Uo3nv6 ? No3nv6 : Go3nv6);
assign No3nv6 = (~(HADDRI[21] & Bp3nv6));
assign Go3nv6 = (~(Ip3nv6 & HADDRI[18]));
assign Al3nv6 = (Pp3nv6 & Wp3nv6);
assign Wp3nv6 = (Rq3nv6 ? Kq3nv6 : Dq3nv6);
assign Kq3nv6 = (Yq3nv6 | Fr3nv6);
assign Dq3nv6 = (~(HADDRI[9] & Mr3nv6));
assign Pp3nv6 = (Hs3nv6 ? As3nv6 : Tr3nv6);
assign As3nv6 = (~(Os3nv6 & HADDRI[12]));
assign Tr3nv6 = (~(HADDRI[15] & Vs3nv6));
assign Pumet6 = (~(Ct3nv6 & Jt3nv6));
assign Jt3nv6 = (Qt3nv6 & Xt3nv6);
assign Xt3nv6 = (Su3nv6 ? Lu3nv6 : Eu3nv6);
assign Lu3nv6 = (~(Zu3nv6 & HADDRI[23]));
assign Eu3nv6 = (~(HADDRI[26] & Gv3nv6));
assign Qt3nv6 = (Nv3nv6 & Uv3nv6);
assign Uv3nv6 = (Gv3nv6 | Bw3nv6);
assign Nv3nv6 = (Ww3nv6 ? Pw3nv6 : Iw3nv6);
assign Pw3nv6 = (~(Dx3nv6 & HADDRI[17]));
assign Iw3nv6 = (~(HADDRI[20] & Kx3nv6));
assign Ct3nv6 = (Rx3nv6 & Yx3nv6);
assign Yx3nv6 = (Ty3nv6 ? My3nv6 : Fy3nv6);
assign My3nv6 = (Az3nv6 | Hz3nv6);
assign Fy3nv6 = (~(HADDRI[8] & Oz3nv6));
assign Rx3nv6 = (J04nv6 ? C04nv6 : Vz3nv6);
assign C04nv6 = (~(Q04nv6 & HADDRI[11]));
assign Vz3nv6 = (~(HADDRI[14] & X04nv6));
assign P1net6 = (~(E14nv6 & L14nv6));
assign L14nv6 = (S14nv6 & Z14nv6);
assign Z14nv6 = (Oe3nv6 ? N24nv6 : G24nv6);
assign N24nv6 = (~(U24nv6 & Ve3nv6));
assign G24nv6 = (Jf3nv6 | B34nv6);
assign S14nv6 = (I34nv6 & P34nv6);
assign P34nv6 = (Ve3nv6 | W34nv6);
assign I34nv6 = (Zg3nv6 ? K44nv6 : D44nv6);
assign K44nv6 = (~(Gh3nv6 & R44nv6));
assign D44nv6 = (~(Y44nv6 & Jf3nv6));
assign E14nv6 = (F54nv6 & M54nv6);
assign M54nv6 = (Pi3nv6 ? A64nv6 : T54nv6);
assign A64nv6 = (~(H64nv6 & Wi3nv6));
assign T54nv6 = (Dj3nv6 | O64nv6);
assign F54nv6 = (Fk3nv6 ? C74nv6 : V64nv6);
assign C74nv6 = (J74nv6 | Gh3nv6);
assign V64nv6 = (~(Tk3nv6 & Q74nv6));
assign C5net6 = (~(X74nv6 & E84nv6));
assign E84nv6 = (L84nv6 & S84nv6);
assign S84nv6 = (Qm3nv6 ? G94nv6 : Z84nv6);
assign G94nv6 = (~(Xm3nv6 & N94nv6));
assign Z84nv6 = (~(U94nv6 & En3nv6));
assign L84nv6 = (Ba4nv6 & Ia4nv6);
assign Ia4nv6 = (En3nv6 | Pa4nv6);
assign Ba4nv6 = (Uo3nv6 ? Db4nv6 : Wa4nv6);
assign Db4nv6 = (Kb4nv6 | Xm3nv6);
assign Wa4nv6 = (~(Ip3nv6 & Rb4nv6));
assign X74nv6 = (Yb4nv6 & Fc4nv6);
assign Fc4nv6 = (Rq3nv6 ? Tc4nv6 : Mc4nv6);
assign Tc4nv6 = (Ad4nv6 | Fr3nv6);
assign Mc4nv6 = (~(Hd4nv6 & Mr3nv6));
assign Yb4nv6 = (Hs3nv6 ? Vd4nv6 : Od4nv6);
assign Vd4nv6 = (~(Os3nv6 & Ce4nv6));
assign Od4nv6 = (~(Je4nv6 & Vs3nv6));
assign P8net6 = (~(Qe4nv6 & Xe4nv6));
assign Xe4nv6 = (Ef4nv6 & Lf4nv6);
assign Lf4nv6 = (Su3nv6 ? Zf4nv6 : Sf4nv6);
assign Zf4nv6 = (Kx3nv6 | Gg4nv6);
assign Sf4nv6 = (Ng4nv6 | Ug4nv6);
assign Ug4nv6 = (!Gv3nv6);
assign Ef4nv6 = (Bh4nv6 & Ih4nv6);
assign Ih4nv6 = (Gv3nv6 | Ph4nv6);
assign Bh4nv6 = (Ww3nv6 ? Di4nv6 : Wh4nv6);
assign Di4nv6 = (X04nv6 | Ki4nv6);
assign Wh4nv6 = (Ri4nv6 | Zu3nv6);
assign Qe4nv6 = (Yi4nv6 & Fj4nv6);
assign Fj4nv6 = (Ty3nv6 ? Tj4nv6 : Mj4nv6);
assign Tj4nv6 = (Ak4nv6 | Hz3nv6);
assign Mj4nv6 = (~(Hk4nv6 & Oz3nv6));
assign Yi4nv6 = (J04nv6 ? Vk4nv6 : Ok4nv6);
assign Vk4nv6 = (~(Q04nv6 & Cl4nv6));
assign Ok4nv6 = (~(Jl4nv6 & X04nv6));
assign L8m7z6[7] = (Vbm7z6[13] & Ql4nv6);
assign L8m7z6[6] = (~(Xl4nv6 & Em4nv6));
assign Em4nv6 = (~(Vbm7z6[11] & Lm4nv6));
assign Xl4nv6 = (Sm4nv6 & Zm4nv6);
assign Zm4nv6 = (~(Vbm7z6[9] & Gn4nv6));
assign Sm4nv6 = (~(Vbm7z6[12] & Nn4nv6));
assign L8m7z6[5] = (~(Un4nv6 & Bo4nv6));
assign Bo4nv6 = (~(Vbm7z6[9] & Lm4nv6));
assign Un4nv6 = (Io4nv6 & Po4nv6);
assign Po4nv6 = (~(Vbm7z6[12] & Gn4nv6));
assign Io4nv6 = (~(Vbm7z6[11] & Nn4nv6));
assign L8m7z6[4] = (~(Wo4nv6 & Dp4nv6));
assign Dp4nv6 = (~(Vbm7z6[7] & Lm4nv6));
assign Wo4nv6 = (Kp4nv6 & Rp4nv6);
assign Rp4nv6 = (~(Vbm7z6[8] & Gn4nv6));
assign Kp4nv6 = (~(Vbm7z6[10] & Nn4nv6));
assign L8m7z6[3] = (~(Yp4nv6 & Fq4nv6));
assign Fq4nv6 = (~(Vbm7z6[12] & Lm4nv6));
assign Yp4nv6 = (Mq4nv6 & Tq4nv6);
assign Tq4nv6 = (~(Vbm7z6[11] & Gn4nv6));
assign Mq4nv6 = (~(Vbm7z6[9] & Nn4nv6));
assign L8m7z6[2] = (~(Ar4nv6 & Hr4nv6));
assign Hr4nv6 = (~(Vbm7z6[10] & Lm4nv6));
assign Ar4nv6 = (Or4nv6 & Vr4nv6);
assign Vr4nv6 = (~(Vbm7z6[7] & Gn4nv6));
assign Or4nv6 = (~(Vbm7z6[8] & Nn4nv6));
assign L8m7z6[1] = (~(Cs4nv6 & Js4nv6));
assign Js4nv6 = (~(Vbm7z6[8] & Lm4nv6));
assign Lm4nv6 = (!Qs4nv6);
assign Cs4nv6 = (Xs4nv6 & Et4nv6);
assign Et4nv6 = (~(Vbm7z6[10] & Gn4nv6));
assign Gn4nv6 = (!Lt4nv6);
assign Xs4nv6 = (~(Vbm7z6[7] & Nn4nv6));
assign Nn4nv6 = (!St4nv6);
assign L8m7z6[0] = (Vbm7z6[6] & Ql4nv6);
assign Ql4nv6 = (~(Zt4nv6 & Qs4nv6));
assign Qs4nv6 = (Vbm7z6[3] ? Nu4nv6 : Gu4nv6);
assign Zt4nv6 = (Lt4nv6 & St4nv6);
assign St4nv6 = (Vbm7z6[3] ? Bv4nv6 : Uu4nv6);
assign Bv4nv6 = (Gu4nv6 & Iv4nv6);
assign Iv4nv6 = (~(Pv4nv6 & Wv4nv6));
assign Pv4nv6 = (Vbm7z6[1] & Vbm7z6[2]);
assign Gu4nv6 = (Vbm7z6[5] ? Kw4nv6 : Dw4nv6);
assign Kw4nv6 = (!Rw4nv6);
assign Rw4nv6 = (Vbm7z6[4] ? Fx4nv6 : Yw4nv6);
assign Dw4nv6 = (~(Mx4nv6 & Vbm7z6[1]));
assign Mx4nv6 = (Vbm7z6[4] & Tx4nv6);
assign Lt4nv6 = (Vbm7z6[3] ? Uu4nv6 : Nu4nv6);
assign Uu4nv6 = (Vbm7z6[5] ? Hy4nv6 : Ay4nv6);
assign Hy4nv6 = (!Oy4nv6);
assign Oy4nv6 = (Vbm7z6[4] ? Vy4nv6 : Fx4nv6);
assign Ay4nv6 = (~(Yw4nv6 & Vbm7z6[4]));
assign Nu4nv6 = (Vbm7z6[5] ? Jz4nv6 : Cz4nv6);
assign Jz4nv6 = (!Qz4nv6);
assign Qz4nv6 = (Vbm7z6[4] ? Yw4nv6 : Vy4nv6);
assign Yw4nv6 = (Vbm7z6[2] & Xz4nv6);
assign Xz4nv6 = (!Vbm7z6[1]);
assign Vy4nv6 = (Vbm7z6[1] & Tx4nv6);
assign Cz4nv6 = (~(Vbm7z6[4] & Fx4nv6));
assign Fx4nv6 = (Vbm7z6[1] ^ Tx4nv6);
assign Tx4nv6 = (!Vbm7z6[2]);
assign Pvlet6 = (~(E05nv6 & L05nv6));
assign L05nv6 = (S05nv6 & Z05nv6);
assign Z05nv6 = (U15nv6 ? N15nv6 : G15nv6);
assign N15nv6 = (~(HADDRI[28] & B25nv6));
assign G15nv6 = (~(I25nv6 & HADDRI[25]));
assign S05nv6 = (P25nv6 & W25nv6);
assign W25nv6 = (B25nv6 | Eg3nv6);
assign P25nv6 = (R35nv6 ? K35nv6 : D35nv6);
assign K35nv6 = (~(HADDRI[22] & Y35nv6));
assign D35nv6 = (~(F45nv6 & HADDRI[19]));
assign E05nv6 = (M45nv6 & T45nv6);
assign T45nv6 = (O55nv6 ? H55nv6 : A55nv6);
assign H55nv6 = (~(HADDRI[10] & V55nv6));
assign A55nv6 = (C65nv6 | Kj3nv6);
assign M45nv6 = (X65nv6 ? Q65nv6 : J65nv6);
assign Q65nv6 = (~(HADDRI[16] & E75nv6));
assign J65nv6 = (~(L75nv6 & HADDRI[13]));
assign Czlet6 = (~(S75nv6 & Z75nv6));
assign Z75nv6 = (G85nv6 & N85nv6);
assign N85nv6 = (I95nv6 ? B95nv6 : U85nv6);
assign B95nv6 = (~(HADDRI[27] & P95nv6));
assign U85nv6 = (~(W95nv6 & HADDRI[24]));
assign G85nv6 = (Da5nv6 & Ka5nv6);
assign Ka5nv6 = (Zn3nv6 | P95nv6);
assign Da5nv6 = (Fb5nv6 ? Ya5nv6 : Ra5nv6);
assign Ya5nv6 = (~(HADDRI[21] & Mb5nv6));
assign Ra5nv6 = (~(Tb5nv6 & HADDRI[18]));
assign S75nv6 = (Ac5nv6 & Hc5nv6);
assign Hc5nv6 = (Cd5nv6 ? Vc5nv6 : Oc5nv6);
assign Vc5nv6 = (~(HADDRI[9] & Jd5nv6));
assign Oc5nv6 = (Yq3nv6 | Qd5nv6);
assign Ac5nv6 = (Le5nv6 ? Ee5nv6 : Xd5nv6);
assign Ee5nv6 = (~(HADDRI[15] & Se5nv6));
assign Xd5nv6 = (~(Ze5nv6 & HADDRI[12]));
assign P2met6 = (~(Gf5nv6 & Nf5nv6));
assign Nf5nv6 = (Uf5nv6 & Bg5nv6);
assign Bg5nv6 = (Wg5nv6 ? Pg5nv6 : Ig5nv6);
assign Pg5nv6 = (~(HADDRI[26] & Dh5nv6));
assign Ig5nv6 = (~(Kh5nv6 & HADDRI[23]));
assign Uf5nv6 = (Rh5nv6 & Yh5nv6);
assign Yh5nv6 = (Dh5nv6 | Bw3nv6);
assign Rh5nv6 = (Ti5nv6 ? Mi5nv6 : Fi5nv6);
assign Mi5nv6 = (~(HADDRI[20] & Aj5nv6));
assign Fi5nv6 = (~(Hj5nv6 & HADDRI[17]));
assign Gf5nv6 = (Oj5nv6 & Vj5nv6);
assign Vj5nv6 = (Qk5nv6 ? Jk5nv6 : Ck5nv6);
assign Jk5nv6 = (Az3nv6 | Xk5nv6);
assign Ck5nv6 = (~(HADDRI[8] & El5nv6));
assign Oj5nv6 = (Zl5nv6 ? Sl5nv6 : Ll5nv6);
assign Sl5nv6 = (~(HADDRI[14] & Gm5nv6));
assign Ll5nv6 = (~(Nm5nv6 & HADDRI[11]));
assign P9met6 = (~(Um5nv6 & Bn5nv6));
assign Bn5nv6 = (In5nv6 & Pn5nv6);
assign Pn5nv6 = (F45nv6 ? Do5nv6 : Wn5nv6);
assign Do5nv6 = (~(R44nv6 & Ko5nv6));
assign Wn5nv6 = (Ro5nv6 | J74nv6);
assign In5nv6 = (Yo5nv6 & Fp5nv6);
assign Fp5nv6 = (Mp5nv6 | C65nv6);
assign Mp5nv6 = (~(Tp5nv6 & Aq5nv6));
assign Yo5nv6 = (I25nv6 ? Oq5nv6 : Hq5nv6);
assign Oq5nv6 = (B34nv6 | U15nv6);
assign Hq5nv6 = (~(R35nv6 & Y44nv6));
assign R35nv6 = (!Ko5nv6);
assign Um5nv6 = (Vq5nv6 & Cr5nv6);
assign Cr5nv6 = (L75nv6 ? Qr5nv6 : Jr5nv6);
assign Qr5nv6 = (~(Q74nv6 & Ro5nv6));
assign Jr5nv6 = (~(O55nv6 & H64nv6));
assign Vq5nv6 = (Es5nv6 ? W34nv6 : Xr5nv6);
assign Xr5nv6 = (~(U15nv6 & U24nv6));
assign Cdmet6 = (~(Ls5nv6 & Ss5nv6));
assign Ss5nv6 = (Zs5nv6 & Gt5nv6);
assign Gt5nv6 = (Tb5nv6 ? Ut5nv6 : Nt5nv6);
assign Ut5nv6 = (~(Rb4nv6 & Bu5nv6));
assign Nt5nv6 = (~(Le5nv6 & Je4nv6));
assign Le5nv6 = (!Iu5nv6);
assign Zs5nv6 = (Pu5nv6 & Wu5nv6);
assign Wu5nv6 = (~(Dv5nv6 & Kv5nv6));
assign Dv5nv6 = (~(Qd5nv6 | Cd5nv6));
assign Pu5nv6 = (W95nv6 ? Yv5nv6 : Rv5nv6);
assign Yv5nv6 = (~(N94nv6 & Fw5nv6));
assign Rv5nv6 = (Bu5nv6 | Kb4nv6);
assign Ls5nv6 = (Mw5nv6 & Tw5nv6);
assign Tw5nv6 = (Ze5nv6 ? Hx5nv6 : Ax5nv6);
assign Hx5nv6 = (~(Ce4nv6 & Iu5nv6));
assign Ax5nv6 = (~(Cd5nv6 & Hd4nv6));
assign Mw5nv6 = (Vx5nv6 ? Pa4nv6 : Ox5nv6);
assign Ox5nv6 = (~(I95nv6 & U94nv6));
assign Pgmet6 = (~(Cy5nv6 & Jy5nv6));
assign Jy5nv6 = (Qy5nv6 & Xy5nv6);
assign Xy5nv6 = (Hj5nv6 ? Lz5nv6 : Ez5nv6);
assign Lz5nv6 = (Ki4nv6 | Ti5nv6);
assign Ez5nv6 = (~(Zl5nv6 & Jl4nv6));
assign Zl5nv6 = (!Sz5nv6);
assign Qy5nv6 = (Zz5nv6 & G06nv6);
assign G06nv6 = (~(N06nv6 & Qk5nv6));
assign N06nv6 = (~(Ak4nv6 | Xk5nv6));
assign Zz5nv6 = (Kh5nv6 ? B16nv6 : U06nv6);
assign B16nv6 = (Gg4nv6 | Wg5nv6);
assign U06nv6 = (I16nv6 | Ri4nv6);
assign Cy5nv6 = (P16nv6 & W16nv6);
assign W16nv6 = (Nm5nv6 ? K26nv6 : D26nv6);
assign K26nv6 = (~(Cl4nv6 & Sz5nv6));
assign D26nv6 = (~(Hk4nv6 & R26nv6));
assign P16nv6 = (F36nv6 ? Ph4nv6 : Y26nv6);
assign Y26nv6 = (M36nv6 | Ng4nv6);
assign Dyl7z6[7] = (N1m7z6[13] & T36nv6);
assign Dyl7z6[6] = (~(A46nv6 & H46nv6));
assign H46nv6 = (~(N1m7z6[11] & O46nv6));
assign A46nv6 = (V46nv6 & C56nv6);
assign C56nv6 = (~(N1m7z6[9] & J56nv6));
assign V46nv6 = (~(N1m7z6[12] & Q56nv6));
assign Dyl7z6[5] = (~(X56nv6 & E66nv6));
assign E66nv6 = (~(N1m7z6[9] & O46nv6));
assign X56nv6 = (L66nv6 & S66nv6);
assign S66nv6 = (~(N1m7z6[12] & J56nv6));
assign L66nv6 = (~(N1m7z6[11] & Q56nv6));
assign Dyl7z6[4] = (~(Z66nv6 & G76nv6));
assign G76nv6 = (~(N1m7z6[7] & O46nv6));
assign Z66nv6 = (N76nv6 & U76nv6);
assign U76nv6 = (~(N1m7z6[8] & J56nv6));
assign N76nv6 = (~(N1m7z6[10] & Q56nv6));
assign Dyl7z6[3] = (~(B86nv6 & I86nv6));
assign I86nv6 = (~(N1m7z6[12] & O46nv6));
assign B86nv6 = (P86nv6 & W86nv6);
assign W86nv6 = (~(N1m7z6[11] & J56nv6));
assign P86nv6 = (~(N1m7z6[9] & Q56nv6));
assign Dyl7z6[2] = (~(D96nv6 & K96nv6));
assign K96nv6 = (~(N1m7z6[10] & O46nv6));
assign D96nv6 = (R96nv6 & Y96nv6);
assign Y96nv6 = (~(N1m7z6[7] & J56nv6));
assign R96nv6 = (~(N1m7z6[8] & Q56nv6));
assign Dyl7z6[1] = (~(Fa6nv6 & Ma6nv6));
assign Ma6nv6 = (~(N1m7z6[8] & O46nv6));
assign O46nv6 = (!Ta6nv6);
assign Fa6nv6 = (Ab6nv6 & Hb6nv6);
assign Hb6nv6 = (~(N1m7z6[10] & J56nv6));
assign J56nv6 = (!Ob6nv6);
assign Ab6nv6 = (~(N1m7z6[7] & Q56nv6));
assign Q56nv6 = (!Vb6nv6);
assign Dyl7z6[0] = (N1m7z6[6] & T36nv6);
assign T36nv6 = (~(Cc6nv6 & Ta6nv6));
assign Ta6nv6 = (N1m7z6[3] ? Qc6nv6 : Jc6nv6);
assign Cc6nv6 = (Ob6nv6 & Vb6nv6);
assign Vb6nv6 = (N1m7z6[3] ? Ed6nv6 : Xc6nv6);
assign Ed6nv6 = (Jc6nv6 & Ld6nv6);
assign Ld6nv6 = (~(Sd6nv6 & Zd6nv6));
assign Sd6nv6 = (N1m7z6[2] & N1m7z6[1]);
assign Jc6nv6 = (N1m7z6[5] ? Ne6nv6 : Ge6nv6);
assign Ne6nv6 = (!Ue6nv6);
assign Ue6nv6 = (N1m7z6[4] ? If6nv6 : Bf6nv6);
assign Ge6nv6 = (~(Pf6nv6 & N1m7z6[4]));
assign Ob6nv6 = (N1m7z6[3] ? Xc6nv6 : Qc6nv6);
assign Xc6nv6 = (N1m7z6[5] ? Dg6nv6 : Wf6nv6);
assign Dg6nv6 = (!Kg6nv6);
assign Kg6nv6 = (N1m7z6[4] ? Pf6nv6 : If6nv6);
assign Wf6nv6 = (~(Bf6nv6 & N1m7z6[4]));
assign Qc6nv6 = (N1m7z6[5] ? Yg6nv6 : Rg6nv6);
assign Yg6nv6 = (!Fh6nv6);
assign Fh6nv6 = (N1m7z6[4] ? Bf6nv6 : Pf6nv6);
assign Bf6nv6 = (N1m7z6[2] & Mh6nv6);
assign Mh6nv6 = (!N1m7z6[1]);
assign Pf6nv6 = (N1m7z6[1] & Th6nv6);
assign Rg6nv6 = (~(N1m7z6[4] & If6nv6));
assign If6nv6 = (N1m7z6[1] ^ Th6nv6);
assign Th6nv6 = (!N1m7z6[2]);
assign P3let6 = (~(Ai6nv6 & Hi6nv6));
assign Hi6nv6 = (Oi6nv6 & Vi6nv6);
assign Vi6nv6 = (Qj6nv6 ? Jj6nv6 : Cj6nv6);
assign Jj6nv6 = (~(HADDRI[28] & Xj6nv6));
assign Cj6nv6 = (~(Ek6nv6 & HADDRI[25]));
assign Oi6nv6 = (Lk6nv6 & Sk6nv6);
assign Sk6nv6 = (Xj6nv6 | Eg3nv6);
assign Lk6nv6 = (Nl6nv6 ? Gl6nv6 : Zk6nv6);
assign Gl6nv6 = (~(HADDRI[22] & Ul6nv6));
assign Zk6nv6 = (~(Bm6nv6 & HADDRI[19]));
assign Ai6nv6 = (Im6nv6 & Pm6nv6);
assign Pm6nv6 = (Kn6nv6 ? Dn6nv6 : Wm6nv6);
assign Dn6nv6 = (~(HADDRI[10] & Rn6nv6));
assign Wm6nv6 = (Yn6nv6 | Kj3nv6);
assign Im6nv6 = (To6nv6 ? Mo6nv6 : Fo6nv6);
assign Mo6nv6 = (~(HADDRI[16] & Ap6nv6));
assign Fo6nv6 = (~(Hp6nv6 & HADDRI[13]));
assign C7let6 = (~(Op6nv6 & Vp6nv6));
assign Vp6nv6 = (Cq6nv6 & Jq6nv6);
assign Jq6nv6 = (Er6nv6 ? Xq6nv6 : Qq6nv6);
assign Xq6nv6 = (~(HADDRI[27] & Lr6nv6));
assign Qq6nv6 = (~(Sr6nv6 & HADDRI[24]));
assign Cq6nv6 = (Zr6nv6 & Gs6nv6);
assign Gs6nv6 = (Zn3nv6 | Lr6nv6);
assign Zr6nv6 = (Bt6nv6 ? Us6nv6 : Ns6nv6);
assign Us6nv6 = (~(HADDRI[21] & It6nv6));
assign Ns6nv6 = (~(Pt6nv6 & HADDRI[18]));
assign Op6nv6 = (Wt6nv6 & Du6nv6);
assign Du6nv6 = (Yu6nv6 ? Ru6nv6 : Ku6nv6);
assign Ru6nv6 = (~(HADDRI[9] & Fv6nv6));
assign Ku6nv6 = (Yq3nv6 | Mv6nv6);
assign Wt6nv6 = (Hw6nv6 ? Aw6nv6 : Tv6nv6);
assign Aw6nv6 = (~(HADDRI[15] & Ow6nv6));
assign Tv6nv6 = (~(Vw6nv6 & HADDRI[12]));
assign Palet6 = (~(Cx6nv6 & Jx6nv6));
assign Jx6nv6 = (Qx6nv6 & Xx6nv6);
assign Xx6nv6 = (Sy6nv6 ? Ly6nv6 : Ey6nv6);
assign Ly6nv6 = (~(HADDRI[26] & Zy6nv6));
assign Ey6nv6 = (~(Gz6nv6 & HADDRI[23]));
assign Qx6nv6 = (Nz6nv6 & Uz6nv6);
assign Uz6nv6 = (Zy6nv6 | Bw3nv6);
assign Nz6nv6 = (P07nv6 ? I07nv6 : B07nv6);
assign I07nv6 = (~(HADDRI[20] & W07nv6));
assign B07nv6 = (~(D17nv6 & HADDRI[17]));
assign Cx6nv6 = (K17nv6 & R17nv6);
assign R17nv6 = (M27nv6 ? F27nv6 : Y17nv6);
assign F27nv6 = (Az3nv6 | T27nv6);
assign Y17nv6 = (~(HADDRI[8] & A37nv6));
assign K17nv6 = (V37nv6 ? O37nv6 : H37nv6);
assign O37nv6 = (~(HADDRI[14] & C47nv6));
assign H37nv6 = (~(J47nv6 & HADDRI[11]));
assign Phlet6 = (~(Q47nv6 & X47nv6));
assign X47nv6 = (E57nv6 & L57nv6);
assign L57nv6 = (Bm6nv6 ? Z57nv6 : S57nv6);
assign Z57nv6 = (~(R44nv6 & G67nv6));
assign S57nv6 = (N67nv6 | J74nv6);
assign E57nv6 = (U67nv6 & B77nv6);
assign B77nv6 = (I77nv6 | Yn6nv6);
assign I77nv6 = (~(Tp5nv6 & P77nv6));
assign U67nv6 = (Ek6nv6 ? D87nv6 : W77nv6);
assign D87nv6 = (B34nv6 | Qj6nv6);
assign W77nv6 = (~(Nl6nv6 & Y44nv6));
assign Nl6nv6 = (!G67nv6);
assign Q47nv6 = (K87nv6 & R87nv6);
assign R87nv6 = (Hp6nv6 ? F97nv6 : Y87nv6);
assign F97nv6 = (~(Q74nv6 & N67nv6));
assign Y87nv6 = (~(Kn6nv6 & H64nv6));
assign K87nv6 = (T97nv6 ? W34nv6 : M97nv6);
assign M97nv6 = (~(Qj6nv6 & U24nv6));
assign Cllet6 = (~(Aa7nv6 & Ha7nv6));
assign Ha7nv6 = (Oa7nv6 & Va7nv6);
assign Va7nv6 = (Pt6nv6 ? Jb7nv6 : Cb7nv6);
assign Jb7nv6 = (~(Rb4nv6 & Qb7nv6));
assign Cb7nv6 = (~(Hw6nv6 & Je4nv6));
assign Hw6nv6 = (!Xb7nv6);
assign Oa7nv6 = (Ec7nv6 & Lc7nv6);
assign Lc7nv6 = (~(Sc7nv6 & Kv5nv6));
assign Sc7nv6 = (~(Mv6nv6 | Yu6nv6));
assign Ec7nv6 = (Sr6nv6 ? Gd7nv6 : Zc7nv6);
assign Gd7nv6 = (~(N94nv6 & Nd7nv6));
assign Zc7nv6 = (Qb7nv6 | Kb4nv6);
assign Aa7nv6 = (Ud7nv6 & Be7nv6);
assign Be7nv6 = (Vw6nv6 ? Pe7nv6 : Ie7nv6);
assign Pe7nv6 = (~(Ce4nv6 & Xb7nv6));
assign Ie7nv6 = (~(Yu6nv6 & Hd4nv6));
assign Ud7nv6 = (Df7nv6 ? Pa4nv6 : We7nv6);
assign We7nv6 = (~(Er6nv6 & U94nv6));
assign Polet6 = (~(Kf7nv6 & Rf7nv6));
assign Rf7nv6 = (Yf7nv6 & Fg7nv6);
assign Fg7nv6 = (D17nv6 ? Tg7nv6 : Mg7nv6);
assign Tg7nv6 = (Ki4nv6 | P07nv6);
assign Mg7nv6 = (~(V37nv6 & Jl4nv6));
assign V37nv6 = (!Ah7nv6);
assign Yf7nv6 = (Hh7nv6 & Oh7nv6);
assign Oh7nv6 = (~(Vh7nv6 & Ci7nv6));
assign Vh7nv6 = (~(Ji7nv6 | T27nv6));
assign Hh7nv6 = (Gz6nv6 ? Xi7nv6 : Qi7nv6);
assign Xi7nv6 = (Gg4nv6 | Sy6nv6);
assign Qi7nv6 = (Ej7nv6 | Ri4nv6);
assign Kf7nv6 = (Lj7nv6 & Sj7nv6);
assign Sj7nv6 = (J47nv6 ? Gk7nv6 : Zj7nv6);
assign Gk7nv6 = (~(Cl4nv6 & Ah7nv6));
assign Zj7nv6 = (~(Hk4nv6 & Ji7nv6));
assign Lj7nv6 = (Uk7nv6 ? Ph4nv6 : Nk7nv6);
assign Nk7nv6 = (Bl7nv6 | Ng4nv6);
assign Vnl7z6[7] = (Frl7z6[13] & Il7nv6);
assign Vnl7z6[6] = (~(Pl7nv6 & Wl7nv6));
assign Wl7nv6 = (~(Frl7z6[11] & Dm7nv6));
assign Pl7nv6 = (Km7nv6 & Rm7nv6);
assign Rm7nv6 = (~(Frl7z6[9] & Ym7nv6));
assign Km7nv6 = (~(Frl7z6[12] & Fn7nv6));
assign Vnl7z6[5] = (~(Mn7nv6 & Tn7nv6));
assign Tn7nv6 = (~(Frl7z6[9] & Dm7nv6));
assign Mn7nv6 = (Ao7nv6 & Ho7nv6);
assign Ho7nv6 = (~(Frl7z6[12] & Ym7nv6));
assign Ao7nv6 = (~(Frl7z6[11] & Fn7nv6));
assign Vnl7z6[4] = (~(Oo7nv6 & Vo7nv6));
assign Vo7nv6 = (~(Frl7z6[7] & Dm7nv6));
assign Oo7nv6 = (Cp7nv6 & Jp7nv6);
assign Jp7nv6 = (~(Frl7z6[8] & Ym7nv6));
assign Cp7nv6 = (~(Frl7z6[10] & Fn7nv6));
assign Vnl7z6[3] = (~(Qp7nv6 & Xp7nv6));
assign Xp7nv6 = (~(Frl7z6[12] & Dm7nv6));
assign Qp7nv6 = (Eq7nv6 & Lq7nv6);
assign Lq7nv6 = (~(Frl7z6[11] & Ym7nv6));
assign Eq7nv6 = (~(Frl7z6[9] & Fn7nv6));
assign Vnl7z6[2] = (~(Sq7nv6 & Zq7nv6));
assign Zq7nv6 = (~(Frl7z6[10] & Dm7nv6));
assign Sq7nv6 = (Gr7nv6 & Nr7nv6);
assign Nr7nv6 = (~(Frl7z6[7] & Ym7nv6));
assign Gr7nv6 = (~(Frl7z6[8] & Fn7nv6));
assign Vnl7z6[1] = (~(Ur7nv6 & Bs7nv6));
assign Bs7nv6 = (~(Frl7z6[8] & Dm7nv6));
assign Dm7nv6 = (!Is7nv6);
assign Ur7nv6 = (Ps7nv6 & Ws7nv6);
assign Ws7nv6 = (~(Frl7z6[10] & Ym7nv6));
assign Ym7nv6 = (!Dt7nv6);
assign Ps7nv6 = (~(Frl7z6[7] & Fn7nv6));
assign Fn7nv6 = (!Kt7nv6);
assign Vnl7z6[0] = (Frl7z6[6] & Il7nv6);
assign Il7nv6 = (~(Rt7nv6 & Is7nv6));
assign Is7nv6 = (Frl7z6[3] ? Fu7nv6 : Yt7nv6);
assign Rt7nv6 = (Dt7nv6 & Kt7nv6);
assign Kt7nv6 = (Frl7z6[3] ? Tu7nv6 : Mu7nv6);
assign Tu7nv6 = (Yt7nv6 & Av7nv6);
assign Av7nv6 = (~(Hv7nv6 & Ov7nv6));
assign Hv7nv6 = (Frl7z6[1] & Frl7z6[2]);
assign Yt7nv6 = (Frl7z6[5] ? Cw7nv6 : Vv7nv6);
assign Cw7nv6 = (!Jw7nv6);
assign Jw7nv6 = (Frl7z6[4] ? Xw7nv6 : Qw7nv6);
assign Vv7nv6 = (~(Ex7nv6 & Frl7z6[1]));
assign Ex7nv6 = (Frl7z6[4] & Lx7nv6);
assign Dt7nv6 = (Frl7z6[3] ? Mu7nv6 : Fu7nv6);
assign Mu7nv6 = (Frl7z6[5] ? Zx7nv6 : Sx7nv6);
assign Zx7nv6 = (!Gy7nv6);
assign Gy7nv6 = (Frl7z6[4] ? Ny7nv6 : Xw7nv6);
assign Sx7nv6 = (~(Qw7nv6 & Frl7z6[4]));
assign Fu7nv6 = (Frl7z6[5] ? Bz7nv6 : Uy7nv6);
assign Bz7nv6 = (!Iz7nv6);
assign Iz7nv6 = (Frl7z6[4] ? Qw7nv6 : Ny7nv6);
assign Qw7nv6 = (Frl7z6[2] & Pz7nv6);
assign Pz7nv6 = (!Frl7z6[1]);
assign Ny7nv6 = (Frl7z6[1] & Lx7nv6);
assign Uy7nv6 = (~(Frl7z6[4] & Xw7nv6));
assign Xw7nv6 = (Frl7z6[1] ^ Lx7nv6);
assign Lx7nv6 = (!Frl7z6[2]);
assign Pbket6 = (~(Wz7nv6 & D08nv6));
assign D08nv6 = (K08nv6 & R08nv6);
assign R08nv6 = (M18nv6 ? F18nv6 : Y08nv6);
assign F18nv6 = (~(HADDRI[28] & T18nv6));
assign Y08nv6 = (~(A28nv6 & HADDRI[25]));
assign K08nv6 = (H28nv6 & O28nv6);
assign O28nv6 = (T18nv6 | Eg3nv6);
assign H28nv6 = (J38nv6 ? C38nv6 : V28nv6);
assign C38nv6 = (~(HADDRI[22] & Q38nv6));
assign V28nv6 = (~(X38nv6 & HADDRI[19]));
assign Wz7nv6 = (E48nv6 & L48nv6);
assign L48nv6 = (G58nv6 ? Z48nv6 : S48nv6);
assign Z48nv6 = (~(HADDRI[10] & N58nv6));
assign S48nv6 = (U58nv6 | Kj3nv6);
assign E48nv6 = (P68nv6 ? I68nv6 : B68nv6);
assign I68nv6 = (~(HADDRI[16] & W68nv6));
assign B68nv6 = (~(D78nv6 & HADDRI[13]));
assign Cfket6 = (~(K78nv6 & R78nv6));
assign R78nv6 = (Y78nv6 & F88nv6);
assign F88nv6 = (A98nv6 ? T88nv6 : M88nv6);
assign T88nv6 = (~(HADDRI[27] & H98nv6));
assign M88nv6 = (~(O98nv6 & HADDRI[24]));
assign Y78nv6 = (V98nv6 & Ca8nv6);
assign Ca8nv6 = (Zn3nv6 | H98nv6);
assign V98nv6 = (Xa8nv6 ? Qa8nv6 : Ja8nv6);
assign Qa8nv6 = (~(HADDRI[21] & Eb8nv6));
assign Ja8nv6 = (~(Lb8nv6 & HADDRI[18]));
assign K78nv6 = (Sb8nv6 & Zb8nv6);
assign Zb8nv6 = (Uc8nv6 ? Nc8nv6 : Gc8nv6);
assign Nc8nv6 = (~(HADDRI[9] & Bd8nv6));
assign Gc8nv6 = (Yq3nv6 | Id8nv6);
assign Sb8nv6 = (De8nv6 ? Wd8nv6 : Pd8nv6);
assign Wd8nv6 = (~(HADDRI[15] & Ke8nv6));
assign Pd8nv6 = (~(Re8nv6 & HADDRI[12]));
assign Piket6 = (~(Ye8nv6 & Ff8nv6));
assign Ff8nv6 = (Mf8nv6 & Tf8nv6);
assign Tf8nv6 = (Og8nv6 ? Hg8nv6 : Ag8nv6);
assign Hg8nv6 = (~(HADDRI[26] & Vg8nv6));
assign Ag8nv6 = (~(Ch8nv6 & HADDRI[23]));
assign Mf8nv6 = (Jh8nv6 & Qh8nv6);
assign Qh8nv6 = (Vg8nv6 | Bw3nv6);
assign Jh8nv6 = (Li8nv6 ? Ei8nv6 : Xh8nv6);
assign Ei8nv6 = (~(HADDRI[20] & Si8nv6));
assign Xh8nv6 = (~(Zi8nv6 & HADDRI[17]));
assign Ye8nv6 = (Gj8nv6 & Nj8nv6);
assign Nj8nv6 = (Ik8nv6 ? Bk8nv6 : Uj8nv6);
assign Bk8nv6 = (Az3nv6 | Pk8nv6);
assign Uj8nv6 = (~(HADDRI[8] & Wk8nv6));
assign Gj8nv6 = (Rl8nv6 ? Kl8nv6 : Dl8nv6);
assign Kl8nv6 = (~(HADDRI[14] & Yl8nv6));
assign Dl8nv6 = (~(Fm8nv6 & HADDRI[11]));
assign Ppket6 = (~(Mm8nv6 & Tm8nv6));
assign Tm8nv6 = (An8nv6 & Hn8nv6);
assign Hn8nv6 = (X38nv6 ? Vn8nv6 : On8nv6);
assign Vn8nv6 = (~(R44nv6 & Co8nv6));
assign On8nv6 = (Jo8nv6 | J74nv6);
assign An8nv6 = (Qo8nv6 & Xo8nv6);
assign Xo8nv6 = (Ep8nv6 | U58nv6);
assign Ep8nv6 = (~(Tp5nv6 & Lp8nv6));
assign Qo8nv6 = (A28nv6 ? Zp8nv6 : Sp8nv6);
assign Zp8nv6 = (B34nv6 | M18nv6);
assign Sp8nv6 = (~(J38nv6 & Y44nv6));
assign J38nv6 = (!Co8nv6);
assign Mm8nv6 = (Gq8nv6 & Nq8nv6);
assign Nq8nv6 = (D78nv6 ? Br8nv6 : Uq8nv6);
assign Br8nv6 = (~(Q74nv6 & Jo8nv6));
assign Uq8nv6 = (~(G58nv6 & H64nv6));
assign Gq8nv6 = (Pr8nv6 ? W34nv6 : Ir8nv6);
assign Ir8nv6 = (~(M18nv6 & U24nv6));
assign Ctket6 = (~(Wr8nv6 & Ds8nv6));
assign Ds8nv6 = (Ks8nv6 & Rs8nv6);
assign Rs8nv6 = (Lb8nv6 ? Ft8nv6 : Ys8nv6);
assign Ft8nv6 = (~(Rb4nv6 & Mt8nv6));
assign Ys8nv6 = (~(De8nv6 & Je4nv6));
assign De8nv6 = (!Tt8nv6);
assign Ks8nv6 = (Au8nv6 & Hu8nv6);
assign Hu8nv6 = (~(Ou8nv6 & Kv5nv6));
assign Ou8nv6 = (~(Id8nv6 | Uc8nv6));
assign Au8nv6 = (O98nv6 ? Cv8nv6 : Vu8nv6);
assign Cv8nv6 = (~(N94nv6 & Jv8nv6));
assign Vu8nv6 = (Mt8nv6 | Kb4nv6);
assign Wr8nv6 = (Qv8nv6 & Xv8nv6);
assign Xv8nv6 = (Re8nv6 ? Lw8nv6 : Ew8nv6);
assign Lw8nv6 = (~(Ce4nv6 & Tt8nv6));
assign Ew8nv6 = (~(Uc8nv6 & Hd4nv6));
assign Qv8nv6 = (Zw8nv6 ? Pa4nv6 : Sw8nv6);
assign Sw8nv6 = (~(A98nv6 & U94nv6));
assign Pwket6 = (~(Gx8nv6 & Nx8nv6));
assign Nx8nv6 = (Ux8nv6 & By8nv6);
assign By8nv6 = (Zi8nv6 ? Py8nv6 : Iy8nv6);
assign Py8nv6 = (Ki4nv6 | Li8nv6);
assign Iy8nv6 = (~(Rl8nv6 & Jl4nv6));
assign Rl8nv6 = (!Wy8nv6);
assign Ux8nv6 = (Dz8nv6 & Kz8nv6);
assign Kz8nv6 = (~(Rz8nv6 & Ik8nv6));
assign Rz8nv6 = (~(Ak4nv6 | Pk8nv6));
assign Dz8nv6 = (Ch8nv6 ? F09nv6 : Yz8nv6);
assign F09nv6 = (Gg4nv6 | Og8nv6);
assign Yz8nv6 = (M09nv6 | Ri4nv6);
assign Gx8nv6 = (T09nv6 & A19nv6);
assign A19nv6 = (Fm8nv6 ? O19nv6 : H19nv6);
assign O19nv6 = (~(Cl4nv6 & Wy8nv6));
assign H19nv6 = (~(Hk4nv6 & V19nv6));
assign T09nv6 = (J29nv6 ? Ph4nv6 : C29nv6);
assign C29nv6 = (Q29nv6 | Ng4nv6);
assign Ndl7z6[7] = (Xgl7z6[13] & X29nv6);
assign Ndl7z6[6] = (~(E39nv6 & L39nv6));
assign L39nv6 = (~(Xgl7z6[11] & S39nv6));
assign E39nv6 = (Z39nv6 & G49nv6);
assign G49nv6 = (~(Xgl7z6[9] & N49nv6));
assign Z39nv6 = (~(Xgl7z6[12] & U49nv6));
assign Ndl7z6[5] = (~(B59nv6 & I59nv6));
assign I59nv6 = (~(Xgl7z6[9] & S39nv6));
assign B59nv6 = (P59nv6 & W59nv6);
assign W59nv6 = (~(Xgl7z6[12] & N49nv6));
assign P59nv6 = (~(Xgl7z6[11] & U49nv6));
assign Ndl7z6[4] = (~(D69nv6 & K69nv6));
assign K69nv6 = (~(Xgl7z6[7] & S39nv6));
assign D69nv6 = (R69nv6 & Y69nv6);
assign Y69nv6 = (~(Xgl7z6[8] & N49nv6));
assign R69nv6 = (~(Xgl7z6[10] & U49nv6));
assign Ndl7z6[3] = (~(F79nv6 & M79nv6));
assign M79nv6 = (~(Xgl7z6[12] & S39nv6));
assign F79nv6 = (T79nv6 & A89nv6);
assign A89nv6 = (~(Xgl7z6[11] & N49nv6));
assign T79nv6 = (~(Xgl7z6[9] & U49nv6));
assign Ndl7z6[2] = (~(H89nv6 & O89nv6));
assign O89nv6 = (~(Xgl7z6[10] & S39nv6));
assign H89nv6 = (V89nv6 & C99nv6);
assign C99nv6 = (~(Xgl7z6[7] & N49nv6));
assign V89nv6 = (~(Xgl7z6[8] & U49nv6));
assign Ndl7z6[1] = (~(J99nv6 & Q99nv6));
assign Q99nv6 = (~(Xgl7z6[8] & S39nv6));
assign S39nv6 = (!X99nv6);
assign J99nv6 = (Ea9nv6 & La9nv6);
assign La9nv6 = (~(Xgl7z6[10] & N49nv6));
assign N49nv6 = (!Sa9nv6);
assign Ea9nv6 = (~(Xgl7z6[7] & U49nv6));
assign U49nv6 = (!Za9nv6);
assign Ndl7z6[0] = (Xgl7z6[6] & X29nv6);
assign X29nv6 = (~(Gb9nv6 & X99nv6));
assign X99nv6 = (Xgl7z6[3] ? Ub9nv6 : Nb9nv6);
assign Gb9nv6 = (Sa9nv6 & Za9nv6);
assign Za9nv6 = (Xgl7z6[3] ? Ic9nv6 : Bc9nv6);
assign Ic9nv6 = (Nb9nv6 & Pc9nv6);
assign Pc9nv6 = (~(Wc9nv6 & Dd9nv6));
assign Wc9nv6 = (Xgl7z6[2] & Xgl7z6[1]);
assign Nb9nv6 = (Xgl7z6[5] ? Rd9nv6 : Kd9nv6);
assign Rd9nv6 = (!Yd9nv6);
assign Yd9nv6 = (Xgl7z6[4] ? Me9nv6 : Fe9nv6);
assign Kd9nv6 = (~(Te9nv6 & Xgl7z6[4]));
assign Sa9nv6 = (Xgl7z6[3] ? Bc9nv6 : Ub9nv6);
assign Bc9nv6 = (Xgl7z6[5] ? Hf9nv6 : Af9nv6);
assign Hf9nv6 = (!Of9nv6);
assign Of9nv6 = (Xgl7z6[4] ? Te9nv6 : Me9nv6);
assign Af9nv6 = (~(Fe9nv6 & Xgl7z6[4]));
assign Ub9nv6 = (Xgl7z6[5] ? Cg9nv6 : Vf9nv6);
assign Cg9nv6 = (!Jg9nv6);
assign Jg9nv6 = (Xgl7z6[4] ? Fe9nv6 : Te9nv6);
assign Fe9nv6 = (Xgl7z6[2] & Qg9nv6);
assign Qg9nv6 = (!Xgl7z6[1]);
assign Te9nv6 = (Xgl7z6[1] & Xg9nv6);
assign Vf9nv6 = (~(Xgl7z6[4] & Me9nv6));
assign Me9nv6 = (Xgl7z6[1] ^ Xg9nv6);
assign Xg9nv6 = (!Xgl7z6[2]);
assign Pjjet6 = (~(Eh9nv6 & Lh9nv6));
assign Lh9nv6 = (Sh9nv6 & Zh9nv6);
assign Zh9nv6 = (Ui9nv6 ? Ni9nv6 : Gi9nv6);
assign Ni9nv6 = (~(HADDRI[28] & Bj9nv6));
assign Gi9nv6 = (~(Ij9nv6 & HADDRI[25]));
assign Sh9nv6 = (Pj9nv6 & Wj9nv6);
assign Wj9nv6 = (Bj9nv6 | Eg3nv6);
assign Pj9nv6 = (Rk9nv6 ? Kk9nv6 : Dk9nv6);
assign Kk9nv6 = (~(HADDRI[22] & Yk9nv6));
assign Dk9nv6 = (~(Fl9nv6 & HADDRI[19]));
assign Eh9nv6 = (Ml9nv6 & Tl9nv6);
assign Tl9nv6 = (Om9nv6 ? Hm9nv6 : Am9nv6);
assign Hm9nv6 = (~(HADDRI[10] & Vm9nv6));
assign Am9nv6 = (Cn9nv6 | Kj3nv6);
assign Ml9nv6 = (Xn9nv6 ? Qn9nv6 : Jn9nv6);
assign Qn9nv6 = (~(HADDRI[16] & Eo9nv6));
assign Jn9nv6 = (~(Lo9nv6 & HADDRI[13]));
assign Cnjet6 = (~(So9nv6 & Zo9nv6));
assign Zo9nv6 = (Gp9nv6 & Np9nv6);
assign Np9nv6 = (Iq9nv6 ? Bq9nv6 : Up9nv6);
assign Bq9nv6 = (~(HADDRI[27] & Pq9nv6));
assign Up9nv6 = (~(Wq9nv6 & HADDRI[24]));
assign Gp9nv6 = (Dr9nv6 & Kr9nv6);
assign Kr9nv6 = (Zn3nv6 | Pq9nv6);
assign Dr9nv6 = (Fs9nv6 ? Yr9nv6 : Rr9nv6);
assign Yr9nv6 = (~(HADDRI[21] & Ms9nv6));
assign Rr9nv6 = (~(Ts9nv6 & HADDRI[18]));
assign So9nv6 = (At9nv6 & Ht9nv6);
assign Ht9nv6 = (Cu9nv6 ? Vt9nv6 : Ot9nv6);
assign Vt9nv6 = (~(HADDRI[9] & Ju9nv6));
assign Ot9nv6 = (Yq3nv6 | Qu9nv6);
assign At9nv6 = (Lv9nv6 ? Ev9nv6 : Xu9nv6);
assign Ev9nv6 = (~(HADDRI[15] & Sv9nv6));
assign Xu9nv6 = (~(Zv9nv6 & HADDRI[12]));
assign Pqjet6 = (~(Gw9nv6 & Nw9nv6));
assign Nw9nv6 = (Uw9nv6 & Bx9nv6);
assign Bx9nv6 = (Wx9nv6 ? Px9nv6 : Ix9nv6);
assign Px9nv6 = (~(HADDRI[26] & Dy9nv6));
assign Ix9nv6 = (~(Ky9nv6 & HADDRI[23]));
assign Uw9nv6 = (Ry9nv6 & Yy9nv6);
assign Yy9nv6 = (Dy9nv6 | Bw3nv6);
assign Ry9nv6 = (Tz9nv6 ? Mz9nv6 : Fz9nv6);
assign Mz9nv6 = (~(HADDRI[20] & A0anv6));
assign Fz9nv6 = (~(H0anv6 & HADDRI[17]));
assign Gw9nv6 = (O0anv6 & V0anv6);
assign V0anv6 = (Q1anv6 ? J1anv6 : C1anv6);
assign J1anv6 = (Az3nv6 | X1anv6);
assign C1anv6 = (~(HADDRI[8] & E2anv6));
assign O0anv6 = (Z2anv6 ? S2anv6 : L2anv6);
assign S2anv6 = (~(HADDRI[14] & G3anv6));
assign L2anv6 = (~(N3anv6 & HADDRI[11]));
assign Pxjet6 = (~(U3anv6 & B4anv6));
assign B4anv6 = (I4anv6 & P4anv6);
assign P4anv6 = (Fl9nv6 ? D5anv6 : W4anv6);
assign D5anv6 = (~(R44nv6 & K5anv6));
assign W4anv6 = (R5anv6 | J74nv6);
assign I4anv6 = (Y5anv6 & F6anv6);
assign F6anv6 = (M6anv6 | Cn9nv6);
assign M6anv6 = (~(Tp5nv6 & T6anv6));
assign Y5anv6 = (Ij9nv6 ? H7anv6 : A7anv6);
assign H7anv6 = (B34nv6 | Ui9nv6);
assign A7anv6 = (~(Rk9nv6 & Y44nv6));
assign Rk9nv6 = (!K5anv6);
assign U3anv6 = (O7anv6 & V7anv6);
assign V7anv6 = (Lo9nv6 ? J8anv6 : C8anv6);
assign J8anv6 = (~(Q74nv6 & R5anv6));
assign C8anv6 = (~(Om9nv6 & H64nv6));
assign O7anv6 = (X8anv6 ? W34nv6 : Q8anv6);
assign Q8anv6 = (~(Ui9nv6 & U24nv6));
assign C1ket6 = (~(E9anv6 & L9anv6));
assign L9anv6 = (S9anv6 & Z9anv6);
assign Z9anv6 = (Ts9nv6 ? Naanv6 : Gaanv6);
assign Naanv6 = (~(Rb4nv6 & Uaanv6));
assign Gaanv6 = (~(Lv9nv6 & Je4nv6));
assign Lv9nv6 = (!Bbanv6);
assign S9anv6 = (Ibanv6 & Pbanv6);
assign Pbanv6 = (~(Wbanv6 & Kv5nv6));
assign Wbanv6 = (~(Qu9nv6 | Cu9nv6));
assign Ibanv6 = (Wq9nv6 ? Kcanv6 : Dcanv6);
assign Kcanv6 = (~(N94nv6 & Rcanv6));
assign Dcanv6 = (Uaanv6 | Kb4nv6);
assign E9anv6 = (Ycanv6 & Fdanv6);
assign Fdanv6 = (Zv9nv6 ? Tdanv6 : Mdanv6);
assign Tdanv6 = (~(Ce4nv6 & Bbanv6));
assign Mdanv6 = (~(Cu9nv6 & Hd4nv6));
assign Ycanv6 = (Heanv6 ? Pa4nv6 : Aeanv6);
assign Aeanv6 = (~(Iq9nv6 & U94nv6));
assign P4ket6 = (~(Oeanv6 & Veanv6));
assign Veanv6 = (Cfanv6 & Jfanv6);
assign Jfanv6 = (H0anv6 ? Xfanv6 : Qfanv6);
assign Xfanv6 = (Ki4nv6 | Tz9nv6);
assign Qfanv6 = (~(Z2anv6 & Jl4nv6));
assign Z2anv6 = (!Eganv6);
assign Cfanv6 = (Lganv6 & Sganv6);
assign Sganv6 = (~(Zganv6 & Q1anv6));
assign Zganv6 = (~(Ak4nv6 | X1anv6));
assign Lganv6 = (Ky9nv6 ? Nhanv6 : Ghanv6);
assign Nhanv6 = (Gg4nv6 | Wx9nv6);
assign Ghanv6 = (Uhanv6 | Ri4nv6);
assign Oeanv6 = (Bianv6 & Iianv6);
assign Iianv6 = (N3anv6 ? Wianv6 : Pianv6);
assign Wianv6 = (~(Cl4nv6 & Eganv6));
assign Pianv6 = (~(Hk4nv6 & Djanv6));
assign Bianv6 = (Rjanv6 ? Ph4nv6 : Kjanv6);
assign Kjanv6 = (Yjanv6 | Ng4nv6);
assign F3l7z6[7] = (P6l7z6[13] & Fkanv6);
assign F3l7z6[6] = (~(Mkanv6 & Tkanv6));
assign Tkanv6 = (~(P6l7z6[11] & Alanv6));
assign Mkanv6 = (Hlanv6 & Olanv6);
assign Olanv6 = (~(P6l7z6[9] & Vlanv6));
assign Hlanv6 = (~(P6l7z6[12] & Cmanv6));
assign F3l7z6[5] = (~(Jmanv6 & Qmanv6));
assign Qmanv6 = (~(P6l7z6[9] & Alanv6));
assign Jmanv6 = (Xmanv6 & Enanv6);
assign Enanv6 = (~(P6l7z6[12] & Vlanv6));
assign Xmanv6 = (~(P6l7z6[11] & Cmanv6));
assign F3l7z6[4] = (~(Lnanv6 & Snanv6));
assign Snanv6 = (~(P6l7z6[7] & Alanv6));
assign Lnanv6 = (Znanv6 & Goanv6);
assign Goanv6 = (~(P6l7z6[8] & Vlanv6));
assign Znanv6 = (~(P6l7z6[10] & Cmanv6));
assign F3l7z6[3] = (~(Noanv6 & Uoanv6));
assign Uoanv6 = (~(P6l7z6[12] & Alanv6));
assign Noanv6 = (Bpanv6 & Ipanv6);
assign Ipanv6 = (~(P6l7z6[11] & Vlanv6));
assign Bpanv6 = (~(P6l7z6[9] & Cmanv6));
assign F3l7z6[2] = (~(Ppanv6 & Wpanv6));
assign Wpanv6 = (~(P6l7z6[10] & Alanv6));
assign Ppanv6 = (Dqanv6 & Kqanv6);
assign Kqanv6 = (~(P6l7z6[7] & Vlanv6));
assign Dqanv6 = (~(P6l7z6[8] & Cmanv6));
assign F3l7z6[1] = (~(Rqanv6 & Yqanv6));
assign Yqanv6 = (~(P6l7z6[8] & Alanv6));
assign Alanv6 = (!Franv6);
assign Rqanv6 = (Mranv6 & Tranv6);
assign Tranv6 = (~(P6l7z6[10] & Vlanv6));
assign Vlanv6 = (!Asanv6);
assign Mranv6 = (~(P6l7z6[7] & Cmanv6));
assign Cmanv6 = (!Hsanv6);
assign F3l7z6[0] = (P6l7z6[6] & Fkanv6);
assign Fkanv6 = (~(Osanv6 & Franv6));
assign Franv6 = (P6l7z6[3] ? Ctanv6 : Vsanv6);
assign Osanv6 = (Asanv6 & Hsanv6);
assign Hsanv6 = (P6l7z6[3] ? Qtanv6 : Jtanv6);
assign Qtanv6 = (Vsanv6 & Xtanv6);
assign Xtanv6 = (~(Euanv6 & Luanv6));
assign Euanv6 = (P6l7z6[1] & P6l7z6[2]);
assign Vsanv6 = (P6l7z6[5] ? Zuanv6 : Suanv6);
assign Zuanv6 = (!Gvanv6);
assign Gvanv6 = (P6l7z6[4] ? Uvanv6 : Nvanv6);
assign Suanv6 = (~(Bwanv6 & P6l7z6[1]));
assign Bwanv6 = (P6l7z6[4] & Iwanv6);
assign Asanv6 = (P6l7z6[3] ? Jtanv6 : Ctanv6);
assign Jtanv6 = (P6l7z6[5] ? Wwanv6 : Pwanv6);
assign Wwanv6 = (!Dxanv6);
assign Dxanv6 = (P6l7z6[4] ? Kxanv6 : Uvanv6);
assign Pwanv6 = (~(Nvanv6 & P6l7z6[4]));
assign Ctanv6 = (P6l7z6[5] ? Yxanv6 : Rxanv6);
assign Yxanv6 = (!Fyanv6);
assign Fyanv6 = (P6l7z6[4] ? Nvanv6 : Kxanv6);
assign Nvanv6 = (P6l7z6[2] & Myanv6);
assign Myanv6 = (!P6l7z6[1]);
assign Kxanv6 = (P6l7z6[1] & Iwanv6);
assign Rxanv6 = (~(P6l7z6[4] & Uvanv6));
assign Uvanv6 = (P6l7z6[1] ^ Iwanv6);
assign Iwanv6 = (!P6l7z6[2]);
assign Priet6 = (~(Tyanv6 & Azanv6));
assign Azanv6 = (Hzanv6 & Ozanv6);
assign Ozanv6 = (J0bnv6 ? C0bnv6 : Vzanv6);
assign C0bnv6 = (~(HADDRI[28] & Q0bnv6));
assign Vzanv6 = (~(X0bnv6 & HADDRI[25]));
assign Hzanv6 = (E1bnv6 & L1bnv6);
assign L1bnv6 = (Q0bnv6 | Eg3nv6);
assign E1bnv6 = (G2bnv6 ? Z1bnv6 : S1bnv6);
assign Z1bnv6 = (~(HADDRI[22] & N2bnv6));
assign S1bnv6 = (~(U2bnv6 & HADDRI[19]));
assign Tyanv6 = (B3bnv6 & I3bnv6);
assign I3bnv6 = (D4bnv6 ? W3bnv6 : P3bnv6);
assign W3bnv6 = (~(HADDRI[10] & K4bnv6));
assign P3bnv6 = (R4bnv6 | Kj3nv6);
assign B3bnv6 = (M5bnv6 ? F5bnv6 : Y4bnv6);
assign F5bnv6 = (~(HADDRI[16] & T5bnv6));
assign Y4bnv6 = (~(A6bnv6 & HADDRI[13]));
assign Cviet6 = (~(H6bnv6 & O6bnv6));
assign O6bnv6 = (V6bnv6 & C7bnv6);
assign C7bnv6 = (X7bnv6 ? Q7bnv6 : J7bnv6);
assign Q7bnv6 = (~(HADDRI[27] & E8bnv6));
assign J7bnv6 = (~(L8bnv6 & HADDRI[24]));
assign V6bnv6 = (S8bnv6 & Z8bnv6);
assign Z8bnv6 = (Zn3nv6 | E8bnv6);
assign S8bnv6 = (U9bnv6 ? N9bnv6 : G9bnv6);
assign N9bnv6 = (~(HADDRI[21] & Babnv6));
assign G9bnv6 = (~(Iabnv6 & HADDRI[18]));
assign H6bnv6 = (Pabnv6 & Wabnv6);
assign Wabnv6 = (Rbbnv6 ? Kbbnv6 : Dbbnv6);
assign Kbbnv6 = (~(HADDRI[9] & Ybbnv6));
assign Dbbnv6 = (Yq3nv6 | Fcbnv6);
assign Pabnv6 = (Adbnv6 ? Tcbnv6 : Mcbnv6);
assign Tcbnv6 = (~(HADDRI[15] & Hdbnv6));
assign Mcbnv6 = (~(Odbnv6 & HADDRI[12]));
assign Pyiet6 = (~(Vdbnv6 & Cebnv6));
assign Cebnv6 = (Jebnv6 & Qebnv6);
assign Qebnv6 = (Lfbnv6 ? Efbnv6 : Xebnv6);
assign Efbnv6 = (~(HADDRI[26] & Sfbnv6));
assign Xebnv6 = (~(Zfbnv6 & HADDRI[23]));
assign Jebnv6 = (Ggbnv6 & Ngbnv6);
assign Ngbnv6 = (Sfbnv6 | Bw3nv6);
assign Ggbnv6 = (Ihbnv6 ? Bhbnv6 : Ugbnv6);
assign Bhbnv6 = (~(HADDRI[20] & Phbnv6));
assign Ugbnv6 = (~(Whbnv6 & HADDRI[17]));
assign Vdbnv6 = (Dibnv6 & Kibnv6);
assign Kibnv6 = (Fjbnv6 ? Yibnv6 : Ribnv6);
assign Yibnv6 = (Az3nv6 | Mjbnv6);
assign Ribnv6 = (~(HADDRI[8] & Tjbnv6));
assign Dibnv6 = (Okbnv6 ? Hkbnv6 : Akbnv6);
assign Hkbnv6 = (~(HADDRI[14] & Vkbnv6));
assign Akbnv6 = (~(Clbnv6 & HADDRI[11]));
assign P5jet6 = (~(Jlbnv6 & Qlbnv6));
assign Qlbnv6 = (Xlbnv6 & Embnv6);
assign Embnv6 = (U2bnv6 ? Smbnv6 : Lmbnv6);
assign Smbnv6 = (~(R44nv6 & Zmbnv6));
assign Lmbnv6 = (Gnbnv6 | J74nv6);
assign Xlbnv6 = (Nnbnv6 & Unbnv6);
assign Unbnv6 = (Bobnv6 | R4bnv6);
assign Bobnv6 = (~(Tp5nv6 & Iobnv6));
assign Nnbnv6 = (X0bnv6 ? Wobnv6 : Pobnv6);
assign Wobnv6 = (B34nv6 | J0bnv6);
assign Pobnv6 = (~(G2bnv6 & Y44nv6));
assign G2bnv6 = (!Zmbnv6);
assign Jlbnv6 = (Dpbnv6 & Kpbnv6);
assign Kpbnv6 = (A6bnv6 ? Ypbnv6 : Rpbnv6);
assign Ypbnv6 = (~(Q74nv6 & Gnbnv6));
assign Rpbnv6 = (~(D4bnv6 & H64nv6));
assign Dpbnv6 = (Mqbnv6 ? W34nv6 : Fqbnv6);
assign Fqbnv6 = (~(J0bnv6 & U24nv6));
assign C9jet6 = (~(Tqbnv6 & Arbnv6));
assign Arbnv6 = (Hrbnv6 & Orbnv6);
assign Orbnv6 = (Iabnv6 ? Csbnv6 : Vrbnv6);
assign Csbnv6 = (~(Rb4nv6 & Jsbnv6));
assign Vrbnv6 = (~(Adbnv6 & Je4nv6));
assign Adbnv6 = (!Qsbnv6);
assign Hrbnv6 = (Xsbnv6 & Etbnv6);
assign Etbnv6 = (~(Ltbnv6 & Kv5nv6));
assign Ltbnv6 = (~(Fcbnv6 | Rbbnv6));
assign Xsbnv6 = (L8bnv6 ? Ztbnv6 : Stbnv6);
assign Ztbnv6 = (~(N94nv6 & Gubnv6));
assign Stbnv6 = (Jsbnv6 | Kb4nv6);
assign Tqbnv6 = (Nubnv6 & Uubnv6);
assign Uubnv6 = (Odbnv6 ? Ivbnv6 : Bvbnv6);
assign Ivbnv6 = (~(Ce4nv6 & Qsbnv6));
assign Bvbnv6 = (~(Rbbnv6 & Hd4nv6));
assign Nubnv6 = (Wvbnv6 ? Pa4nv6 : Pvbnv6);
assign Pvbnv6 = (~(X7bnv6 & U94nv6));
assign Pcjet6 = (~(Dwbnv6 & Kwbnv6));
assign Kwbnv6 = (Rwbnv6 & Ywbnv6);
assign Ywbnv6 = (Whbnv6 ? Mxbnv6 : Fxbnv6);
assign Mxbnv6 = (Ki4nv6 | Ihbnv6);
assign Fxbnv6 = (~(Okbnv6 & Jl4nv6));
assign Okbnv6 = (!Txbnv6);
assign Rwbnv6 = (Aybnv6 & Hybnv6);
assign Hybnv6 = (~(Oybnv6 & Fjbnv6));
assign Oybnv6 = (~(Ak4nv6 | Mjbnv6));
assign Aybnv6 = (Zfbnv6 ? Czbnv6 : Vybnv6);
assign Czbnv6 = (Gg4nv6 | Lfbnv6);
assign Vybnv6 = (Jzbnv6 | Ri4nv6);
assign Dwbnv6 = (Qzbnv6 & Xzbnv6);
assign Xzbnv6 = (Clbnv6 ? L0cnv6 : E0cnv6);
assign L0cnv6 = (~(Cl4nv6 & Txbnv6));
assign E0cnv6 = (~(Hk4nv6 & S0cnv6));
assign Qzbnv6 = (G1cnv6 ? Ph4nv6 : Z0cnv6);
assign Z0cnv6 = (N1cnv6 | Ng4nv6);
assign Xsk7z6[7] = (Hwk7z6[13] & U1cnv6);
assign Xsk7z6[6] = (~(B2cnv6 & I2cnv6));
assign I2cnv6 = (~(Hwk7z6[11] & P2cnv6));
assign B2cnv6 = (W2cnv6 & D3cnv6);
assign D3cnv6 = (~(Hwk7z6[9] & K3cnv6));
assign W2cnv6 = (~(Hwk7z6[12] & R3cnv6));
assign Xsk7z6[5] = (~(Y3cnv6 & F4cnv6));
assign F4cnv6 = (~(Hwk7z6[9] & P2cnv6));
assign Y3cnv6 = (M4cnv6 & T4cnv6);
assign T4cnv6 = (~(Hwk7z6[12] & K3cnv6));
assign M4cnv6 = (~(Hwk7z6[11] & R3cnv6));
assign Xsk7z6[4] = (~(A5cnv6 & H5cnv6));
assign H5cnv6 = (~(Hwk7z6[7] & P2cnv6));
assign A5cnv6 = (O5cnv6 & V5cnv6);
assign V5cnv6 = (~(Hwk7z6[8] & K3cnv6));
assign O5cnv6 = (~(Hwk7z6[10] & R3cnv6));
assign Xsk7z6[3] = (~(C6cnv6 & J6cnv6));
assign J6cnv6 = (~(Hwk7z6[12] & P2cnv6));
assign C6cnv6 = (Q6cnv6 & X6cnv6);
assign X6cnv6 = (~(Hwk7z6[11] & K3cnv6));
assign Q6cnv6 = (~(Hwk7z6[9] & R3cnv6));
assign Xsk7z6[2] = (~(E7cnv6 & L7cnv6));
assign L7cnv6 = (~(Hwk7z6[10] & P2cnv6));
assign E7cnv6 = (S7cnv6 & Z7cnv6);
assign Z7cnv6 = (~(Hwk7z6[7] & K3cnv6));
assign S7cnv6 = (~(Hwk7z6[8] & R3cnv6));
assign Xsk7z6[1] = (~(G8cnv6 & N8cnv6));
assign N8cnv6 = (~(Hwk7z6[8] & P2cnv6));
assign P2cnv6 = (!U8cnv6);
assign G8cnv6 = (B9cnv6 & I9cnv6);
assign I9cnv6 = (~(Hwk7z6[10] & K3cnv6));
assign K3cnv6 = (!P9cnv6);
assign B9cnv6 = (~(Hwk7z6[7] & R3cnv6));
assign R3cnv6 = (!W9cnv6);
assign Xsk7z6[0] = (Hwk7z6[6] & U1cnv6);
assign U1cnv6 = (~(Dacnv6 & U8cnv6));
assign U8cnv6 = (Hwk7z6[3] ? Racnv6 : Kacnv6);
assign Dacnv6 = (P9cnv6 & W9cnv6);
assign W9cnv6 = (Hwk7z6[3] ? Fbcnv6 : Yacnv6);
assign Fbcnv6 = (Kacnv6 & Mbcnv6);
assign Mbcnv6 = (~(Tbcnv6 & Accnv6));
assign Tbcnv6 = (Hwk7z6[2] & Hwk7z6[1]);
assign Kacnv6 = (Hwk7z6[5] ? Occnv6 : Hccnv6);
assign Occnv6 = (!Vccnv6);
assign Vccnv6 = (Hwk7z6[4] ? Jdcnv6 : Cdcnv6);
assign Hccnv6 = (~(Qdcnv6 & Hwk7z6[4]));
assign P9cnv6 = (Hwk7z6[3] ? Yacnv6 : Racnv6);
assign Yacnv6 = (Hwk7z6[5] ? Eecnv6 : Xdcnv6);
assign Eecnv6 = (!Lecnv6);
assign Lecnv6 = (Hwk7z6[4] ? Qdcnv6 : Jdcnv6);
assign Xdcnv6 = (~(Cdcnv6 & Hwk7z6[4]));
assign Racnv6 = (Hwk7z6[5] ? Zecnv6 : Secnv6);
assign Zecnv6 = (!Gfcnv6);
assign Gfcnv6 = (Hwk7z6[4] ? Cdcnv6 : Qdcnv6);
assign Cdcnv6 = (Hwk7z6[2] & Nfcnv6);
assign Nfcnv6 = (!Hwk7z6[1]);
assign Qdcnv6 = (Hwk7z6[1] & Ufcnv6);
assign Secnv6 = (~(Hwk7z6[4] & Jdcnv6));
assign Jdcnv6 = (Hwk7z6[1] ^ Ufcnv6);
assign Ufcnv6 = (!Hwk7z6[2]);
assign Pzhet6 = (~(Bgcnv6 & Igcnv6));
assign Igcnv6 = (Pgcnv6 & Wgcnv6);
assign Wgcnv6 = (Rhcnv6 ? Khcnv6 : Dhcnv6);
assign Khcnv6 = (~(HADDRI[28] & Yhcnv6));
assign Dhcnv6 = (~(Ficnv6 & HADDRI[25]));
assign Pgcnv6 = (Micnv6 & Ticnv6);
assign Ticnv6 = (Yhcnv6 | Eg3nv6);
assign Micnv6 = (Ojcnv6 ? Hjcnv6 : Ajcnv6);
assign Hjcnv6 = (~(HADDRI[22] & Vjcnv6));
assign Ajcnv6 = (~(Ckcnv6 & HADDRI[19]));
assign Bgcnv6 = (Jkcnv6 & Qkcnv6);
assign Qkcnv6 = (Llcnv6 ? Elcnv6 : Xkcnv6);
assign Elcnv6 = (~(HADDRI[10] & Slcnv6));
assign Xkcnv6 = (Zlcnv6 | Kj3nv6);
assign Jkcnv6 = (Umcnv6 ? Nmcnv6 : Gmcnv6);
assign Nmcnv6 = (~(HADDRI[16] & Bncnv6));
assign Gmcnv6 = (~(Incnv6 & HADDRI[13]));
assign C3iet6 = (~(Pncnv6 & Wncnv6));
assign Wncnv6 = (Docnv6 & Kocnv6);
assign Kocnv6 = (Fpcnv6 ? Yocnv6 : Rocnv6);
assign Yocnv6 = (~(HADDRI[27] & Mpcnv6));
assign Rocnv6 = (~(Tpcnv6 & HADDRI[24]));
assign Docnv6 = (Aqcnv6 & Hqcnv6);
assign Hqcnv6 = (Zn3nv6 | Mpcnv6);
assign Aqcnv6 = (Crcnv6 ? Vqcnv6 : Oqcnv6);
assign Vqcnv6 = (~(HADDRI[21] & Jrcnv6));
assign Oqcnv6 = (~(Qrcnv6 & HADDRI[18]));
assign Pncnv6 = (Xrcnv6 & Escnv6);
assign Escnv6 = (Zscnv6 ? Sscnv6 : Lscnv6);
assign Sscnv6 = (~(HADDRI[9] & Gtcnv6));
assign Lscnv6 = (Yq3nv6 | Ntcnv6);
assign Xrcnv6 = (Iucnv6 ? Bucnv6 : Utcnv6);
assign Bucnv6 = (~(HADDRI[15] & Pucnv6));
assign Utcnv6 = (~(Wucnv6 & HADDRI[12]));
assign P6iet6 = (~(Dvcnv6 & Kvcnv6));
assign Kvcnv6 = (Rvcnv6 & Yvcnv6);
assign Yvcnv6 = (Twcnv6 ? Mwcnv6 : Fwcnv6);
assign Mwcnv6 = (~(HADDRI[26] & Axcnv6));
assign Fwcnv6 = (~(Hxcnv6 & HADDRI[23]));
assign Rvcnv6 = (Oxcnv6 & Vxcnv6);
assign Vxcnv6 = (Axcnv6 | Bw3nv6);
assign Oxcnv6 = (Qycnv6 ? Jycnv6 : Cycnv6);
assign Jycnv6 = (~(HADDRI[20] & Xycnv6));
assign Cycnv6 = (~(Ezcnv6 & HADDRI[17]));
assign Dvcnv6 = (Lzcnv6 & Szcnv6);
assign Szcnv6 = (N0dnv6 ? G0dnv6 : Zzcnv6);
assign G0dnv6 = (Az3nv6 | U0dnv6);
assign Zzcnv6 = (~(HADDRI[8] & B1dnv6));
assign Lzcnv6 = (W1dnv6 ? P1dnv6 : I1dnv6);
assign P1dnv6 = (~(HADDRI[14] & D2dnv6));
assign I1dnv6 = (~(K2dnv6 & HADDRI[11]));
assign Pdiet6 = (~(R2dnv6 & Y2dnv6));
assign Y2dnv6 = (F3dnv6 & M3dnv6);
assign M3dnv6 = (Ckcnv6 ? A4dnv6 : T3dnv6);
assign A4dnv6 = (~(R44nv6 & H4dnv6));
assign T3dnv6 = (O4dnv6 | J74nv6);
assign F3dnv6 = (V4dnv6 & C5dnv6);
assign C5dnv6 = (J5dnv6 | Zlcnv6);
assign J5dnv6 = (~(Tp5nv6 & Q5dnv6));
assign V4dnv6 = (Ficnv6 ? E6dnv6 : X5dnv6);
assign E6dnv6 = (B34nv6 | Rhcnv6);
assign X5dnv6 = (~(Ojcnv6 & Y44nv6));
assign Ojcnv6 = (!H4dnv6);
assign R2dnv6 = (L6dnv6 & S6dnv6);
assign S6dnv6 = (Incnv6 ? G7dnv6 : Z6dnv6);
assign G7dnv6 = (~(Q74nv6 & O4dnv6));
assign Z6dnv6 = (~(Llcnv6 & H64nv6));
assign L6dnv6 = (U7dnv6 ? W34nv6 : N7dnv6);
assign N7dnv6 = (~(Rhcnv6 & U24nv6));
assign Chiet6 = (~(B8dnv6 & I8dnv6));
assign I8dnv6 = (P8dnv6 & W8dnv6);
assign W8dnv6 = (Qrcnv6 ? K9dnv6 : D9dnv6);
assign K9dnv6 = (~(Rb4nv6 & R9dnv6));
assign D9dnv6 = (~(Iucnv6 & Je4nv6));
assign Iucnv6 = (!Y9dnv6);
assign P8dnv6 = (Fadnv6 & Madnv6);
assign Madnv6 = (~(Tadnv6 & Kv5nv6));
assign Tadnv6 = (~(Ntcnv6 | Zscnv6));
assign Fadnv6 = (Tpcnv6 ? Hbdnv6 : Abdnv6);
assign Hbdnv6 = (~(N94nv6 & Obdnv6));
assign Abdnv6 = (R9dnv6 | Kb4nv6);
assign B8dnv6 = (Vbdnv6 & Ccdnv6);
assign Ccdnv6 = (Wucnv6 ? Qcdnv6 : Jcdnv6);
assign Qcdnv6 = (~(Ce4nv6 & Y9dnv6));
assign Jcdnv6 = (~(Zscnv6 & Hd4nv6));
assign Vbdnv6 = (Eddnv6 ? Pa4nv6 : Xcdnv6);
assign Xcdnv6 = (~(Fpcnv6 & U94nv6));
assign Pkiet6 = (~(Lddnv6 & Sddnv6));
assign Sddnv6 = (Zddnv6 & Gednv6);
assign Gednv6 = (Ezcnv6 ? Uednv6 : Nednv6);
assign Uednv6 = (Ki4nv6 | Qycnv6);
assign Nednv6 = (~(W1dnv6 & Jl4nv6));
assign W1dnv6 = (!Bfdnv6);
assign Zddnv6 = (Ifdnv6 & Pfdnv6);
assign Pfdnv6 = (~(Wfdnv6 & N0dnv6));
assign Wfdnv6 = (~(Ak4nv6 | U0dnv6));
assign Ifdnv6 = (Hxcnv6 ? Kgdnv6 : Dgdnv6);
assign Kgdnv6 = (Gg4nv6 | Twcnv6);
assign Dgdnv6 = (Rgdnv6 | Ri4nv6);
assign Lddnv6 = (Ygdnv6 & Fhdnv6);
assign Fhdnv6 = (K2dnv6 ? Thdnv6 : Mhdnv6);
assign Thdnv6 = (~(Cl4nv6 & Bfdnv6));
assign Mhdnv6 = (~(Hk4nv6 & Aidnv6));
assign Ygdnv6 = (Oidnv6 ? Ph4nv6 : Hidnv6);
assign Hidnv6 = (Vidnv6 | Ng4nv6);
assign Pik7z6[7] = (Zlk7z6[13] & Cjdnv6);
assign Pik7z6[6] = (~(Jjdnv6 & Qjdnv6));
assign Qjdnv6 = (~(Zlk7z6[11] & Xjdnv6));
assign Jjdnv6 = (Ekdnv6 & Lkdnv6);
assign Lkdnv6 = (~(Zlk7z6[9] & Skdnv6));
assign Ekdnv6 = (~(Zlk7z6[12] & Zkdnv6));
assign Pik7z6[5] = (~(Gldnv6 & Nldnv6));
assign Nldnv6 = (~(Zlk7z6[9] & Xjdnv6));
assign Gldnv6 = (Uldnv6 & Bmdnv6);
assign Bmdnv6 = (~(Zlk7z6[12] & Skdnv6));
assign Uldnv6 = (~(Zlk7z6[11] & Zkdnv6));
assign Pik7z6[4] = (~(Imdnv6 & Pmdnv6));
assign Pmdnv6 = (~(Zlk7z6[7] & Xjdnv6));
assign Imdnv6 = (Wmdnv6 & Dndnv6);
assign Dndnv6 = (~(Zlk7z6[8] & Skdnv6));
assign Wmdnv6 = (~(Zlk7z6[10] & Zkdnv6));
assign Pik7z6[3] = (~(Kndnv6 & Rndnv6));
assign Rndnv6 = (~(Zlk7z6[12] & Xjdnv6));
assign Kndnv6 = (Yndnv6 & Fodnv6);
assign Fodnv6 = (~(Zlk7z6[11] & Skdnv6));
assign Yndnv6 = (~(Zlk7z6[9] & Zkdnv6));
assign Pik7z6[2] = (~(Modnv6 & Todnv6));
assign Todnv6 = (~(Zlk7z6[10] & Xjdnv6));
assign Modnv6 = (Apdnv6 & Hpdnv6);
assign Hpdnv6 = (~(Zlk7z6[7] & Skdnv6));
assign Apdnv6 = (~(Zlk7z6[8] & Zkdnv6));
assign Pik7z6[1] = (~(Opdnv6 & Vpdnv6));
assign Vpdnv6 = (~(Zlk7z6[8] & Xjdnv6));
assign Xjdnv6 = (!Cqdnv6);
assign Opdnv6 = (Jqdnv6 & Qqdnv6);
assign Qqdnv6 = (~(Zlk7z6[10] & Skdnv6));
assign Skdnv6 = (!Xqdnv6);
assign Jqdnv6 = (~(Zlk7z6[7] & Zkdnv6));
assign Zkdnv6 = (!Erdnv6);
assign Pik7z6[0] = (Zlk7z6[6] & Cjdnv6);
assign Cjdnv6 = (~(Lrdnv6 & Cqdnv6));
assign Cqdnv6 = (Zlk7z6[3] ? Zrdnv6 : Srdnv6);
assign Lrdnv6 = (Xqdnv6 & Erdnv6);
assign Erdnv6 = (Zlk7z6[3] ? Nsdnv6 : Gsdnv6);
assign Nsdnv6 = (Srdnv6 & Usdnv6);
assign Usdnv6 = (~(Btdnv6 & Itdnv6));
assign Btdnv6 = (Zlk7z6[1] & Zlk7z6[2]);
assign Srdnv6 = (Zlk7z6[5] ? Wtdnv6 : Ptdnv6);
assign Wtdnv6 = (!Dudnv6);
assign Dudnv6 = (Zlk7z6[4] ? Rudnv6 : Kudnv6);
assign Ptdnv6 = (~(Yudnv6 & Zlk7z6[1]));
assign Yudnv6 = (Zlk7z6[4] & Fvdnv6);
assign Xqdnv6 = (Zlk7z6[3] ? Gsdnv6 : Zrdnv6);
assign Gsdnv6 = (Zlk7z6[5] ? Tvdnv6 : Mvdnv6);
assign Tvdnv6 = (!Awdnv6);
assign Awdnv6 = (Zlk7z6[4] ? Hwdnv6 : Rudnv6);
assign Mvdnv6 = (~(Kudnv6 & Zlk7z6[4]));
assign Zrdnv6 = (Zlk7z6[5] ? Vwdnv6 : Owdnv6);
assign Vwdnv6 = (!Cxdnv6);
assign Cxdnv6 = (Zlk7z6[4] ? Kudnv6 : Hwdnv6);
assign Kudnv6 = (Zlk7z6[2] & Jxdnv6);
assign Jxdnv6 = (!Zlk7z6[1]);
assign Hwdnv6 = (Zlk7z6[1] & Fvdnv6);
assign Owdnv6 = (~(Zlk7z6[4] & Rudnv6));
assign Rudnv6 = (Zlk7z6[1] ^ Fvdnv6);
assign Fvdnv6 = (!Zlk7z6[2]);
assign P7het6 = (~(Qxdnv6 & Xxdnv6));
assign Xxdnv6 = (Eydnv6 & Lydnv6);
assign Lydnv6 = (Gzdnv6 ? Zydnv6 : Sydnv6);
assign Zydnv6 = (~(HADDRI[28] & Nzdnv6));
assign Sydnv6 = (~(Uzdnv6 & HADDRI[25]));
assign Eydnv6 = (B0env6 & I0env6);
assign I0env6 = (Nzdnv6 | Eg3nv6);
assign B0env6 = (D1env6 ? W0env6 : P0env6);
assign W0env6 = (~(HADDRI[22] & K1env6));
assign P0env6 = (~(R1env6 & HADDRI[19]));
assign Qxdnv6 = (Y1env6 & F2env6);
assign F2env6 = (A3env6 ? T2env6 : M2env6);
assign T2env6 = (~(HADDRI[10] & H3env6));
assign M2env6 = (O3env6 | Kj3nv6);
assign Y1env6 = (J4env6 ? C4env6 : V3env6);
assign C4env6 = (~(HADDRI[16] & Q4env6));
assign V3env6 = (~(X4env6 & HADDRI[13]));
assign Cbhet6 = (~(E5env6 & L5env6));
assign L5env6 = (S5env6 & Z5env6);
assign Z5env6 = (U6env6 ? N6env6 : G6env6);
assign N6env6 = (~(HADDRI[27] & B7env6));
assign G6env6 = (~(I7env6 & HADDRI[24]));
assign S5env6 = (P7env6 & W7env6);
assign W7env6 = (Zn3nv6 | B7env6);
assign P7env6 = (R8env6 ? K8env6 : D8env6);
assign K8env6 = (~(HADDRI[21] & Y8env6));
assign D8env6 = (~(F9env6 & HADDRI[18]));
assign E5env6 = (M9env6 & T9env6);
assign T9env6 = (Oaenv6 ? Haenv6 : Aaenv6);
assign Haenv6 = (~(HADDRI[9] & Vaenv6));
assign Aaenv6 = (Yq3nv6 | Cbenv6);
assign M9env6 = (Xbenv6 ? Qbenv6 : Jbenv6);
assign Qbenv6 = (~(HADDRI[15] & Ecenv6));
assign Jbenv6 = (~(Lcenv6 & HADDRI[12]));
assign Pehet6 = (~(Scenv6 & Zcenv6));
assign Zcenv6 = (Gdenv6 & Ndenv6);
assign Ndenv6 = (Ieenv6 ? Beenv6 : Udenv6);
assign Beenv6 = (~(HADDRI[26] & Peenv6));
assign Udenv6 = (~(Weenv6 & HADDRI[23]));
assign Gdenv6 = (Dfenv6 & Kfenv6);
assign Kfenv6 = (Peenv6 | Bw3nv6);
assign Dfenv6 = (Fgenv6 ? Yfenv6 : Rfenv6);
assign Yfenv6 = (~(HADDRI[20] & Mgenv6));
assign Rfenv6 = (~(Tgenv6 & HADDRI[17]));
assign Scenv6 = (Ahenv6 & Hhenv6);
assign Hhenv6 = (Cienv6 ? Vhenv6 : Ohenv6);
assign Vhenv6 = (Az3nv6 | Jienv6);
assign Ohenv6 = (~(HADDRI[8] & Qienv6));
assign Ahenv6 = (Ljenv6 ? Ejenv6 : Xienv6);
assign Ejenv6 = (~(HADDRI[14] & Sjenv6));
assign Xienv6 = (~(Zjenv6 & HADDRI[11]));
assign Plhet6 = (~(Gkenv6 & Nkenv6));
assign Nkenv6 = (Ukenv6 & Blenv6);
assign Blenv6 = (R1env6 ? Plenv6 : Ilenv6);
assign Plenv6 = (~(R44nv6 & Wlenv6));
assign Ilenv6 = (Dmenv6 | J74nv6);
assign Ukenv6 = (Kmenv6 & Rmenv6);
assign Rmenv6 = (Ymenv6 | O3env6);
assign Ymenv6 = (~(Tp5nv6 & Fnenv6));
assign Kmenv6 = (Uzdnv6 ? Tnenv6 : Mnenv6);
assign Tnenv6 = (B34nv6 | Gzdnv6);
assign Mnenv6 = (~(D1env6 & Y44nv6));
assign D1env6 = (!Wlenv6);
assign Gkenv6 = (Aoenv6 & Hoenv6);
assign Hoenv6 = (X4env6 ? Voenv6 : Ooenv6);
assign Voenv6 = (~(Q74nv6 & Dmenv6));
assign Ooenv6 = (~(A3env6 & H64nv6));
assign Aoenv6 = (Jpenv6 ? W34nv6 : Cpenv6);
assign Cpenv6 = (~(Gzdnv6 & U24nv6));
assign Cphet6 = (~(Qpenv6 & Xpenv6));
assign Xpenv6 = (Eqenv6 & Lqenv6);
assign Lqenv6 = (F9env6 ? Zqenv6 : Sqenv6);
assign Zqenv6 = (~(Rb4nv6 & Grenv6));
assign Sqenv6 = (~(Xbenv6 & Je4nv6));
assign Xbenv6 = (!Nrenv6);
assign Eqenv6 = (Urenv6 & Bsenv6);
assign Bsenv6 = (~(Isenv6 & Kv5nv6));
assign Isenv6 = (~(Cbenv6 | Oaenv6));
assign Urenv6 = (I7env6 ? Wsenv6 : Psenv6);
assign Wsenv6 = (~(N94nv6 & Dtenv6));
assign Psenv6 = (Grenv6 | Kb4nv6);
assign Qpenv6 = (Ktenv6 & Rtenv6);
assign Rtenv6 = (Lcenv6 ? Fuenv6 : Ytenv6);
assign Fuenv6 = (~(Ce4nv6 & Nrenv6));
assign Ytenv6 = (~(Oaenv6 & Hd4nv6));
assign Ktenv6 = (Tuenv6 ? Pa4nv6 : Muenv6);
assign Muenv6 = (~(U6env6 & U94nv6));
assign Pshet6 = (~(Avenv6 & Hvenv6));
assign Hvenv6 = (Ovenv6 & Vvenv6);
assign Vvenv6 = (Tgenv6 ? Jwenv6 : Cwenv6);
assign Jwenv6 = (Ki4nv6 | Fgenv6);
assign Cwenv6 = (~(Ljenv6 & Jl4nv6));
assign Ljenv6 = (!Qwenv6);
assign Ovenv6 = (Xwenv6 & Exenv6);
assign Exenv6 = (~(Lxenv6 & Cienv6));
assign Lxenv6 = (~(Ak4nv6 | Jienv6));
assign Xwenv6 = (Weenv6 ? Zxenv6 : Sxenv6);
assign Zxenv6 = (Gg4nv6 | Ieenv6);
assign Sxenv6 = (Gyenv6 | Ri4nv6);
assign Avenv6 = (Nyenv6 & Uyenv6);
assign Uyenv6 = (Zjenv6 ? Izenv6 : Bzenv6);
assign Izenv6 = (~(Cl4nv6 & Qwenv6));
assign Bzenv6 = (~(Hk4nv6 & Pzenv6));
assign Nyenv6 = (D0fnv6 ? Ph4nv6 : Wzenv6);
assign Wzenv6 = (K0fnv6 | Ng4nv6);
assign H8k7z6[7] = (Rbk7z6[13] & R0fnv6);
assign H8k7z6[6] = (~(Y0fnv6 & F1fnv6));
assign F1fnv6 = (~(Rbk7z6[11] & M1fnv6));
assign Y0fnv6 = (T1fnv6 & A2fnv6);
assign A2fnv6 = (~(Rbk7z6[9] & H2fnv6));
assign T1fnv6 = (~(Rbk7z6[12] & O2fnv6));
assign H8k7z6[5] = (~(V2fnv6 & C3fnv6));
assign C3fnv6 = (~(Rbk7z6[9] & M1fnv6));
assign V2fnv6 = (J3fnv6 & Q3fnv6);
assign Q3fnv6 = (~(Rbk7z6[12] & H2fnv6));
assign J3fnv6 = (~(Rbk7z6[11] & O2fnv6));
assign H8k7z6[4] = (~(X3fnv6 & E4fnv6));
assign E4fnv6 = (~(Rbk7z6[7] & M1fnv6));
assign X3fnv6 = (L4fnv6 & S4fnv6);
assign S4fnv6 = (~(Rbk7z6[8] & H2fnv6));
assign L4fnv6 = (~(Rbk7z6[10] & O2fnv6));
assign H8k7z6[3] = (~(Z4fnv6 & G5fnv6));
assign G5fnv6 = (~(Rbk7z6[12] & M1fnv6));
assign Z4fnv6 = (N5fnv6 & U5fnv6);
assign U5fnv6 = (~(Rbk7z6[11] & H2fnv6));
assign N5fnv6 = (~(Rbk7z6[9] & O2fnv6));
assign H8k7z6[2] = (~(B6fnv6 & I6fnv6));
assign I6fnv6 = (~(Rbk7z6[10] & M1fnv6));
assign B6fnv6 = (P6fnv6 & W6fnv6);
assign W6fnv6 = (~(Rbk7z6[7] & H2fnv6));
assign P6fnv6 = (~(Rbk7z6[8] & O2fnv6));
assign H8k7z6[1] = (~(D7fnv6 & K7fnv6));
assign K7fnv6 = (~(Rbk7z6[8] & M1fnv6));
assign M1fnv6 = (!R7fnv6);
assign D7fnv6 = (Y7fnv6 & F8fnv6);
assign F8fnv6 = (~(Rbk7z6[10] & H2fnv6));
assign H2fnv6 = (!M8fnv6);
assign Y7fnv6 = (~(Rbk7z6[7] & O2fnv6));
assign O2fnv6 = (!T8fnv6);
assign H8k7z6[0] = (Rbk7z6[6] & R0fnv6);
assign R0fnv6 = (~(A9fnv6 & R7fnv6));
assign R7fnv6 = (Rbk7z6[3] ? O9fnv6 : H9fnv6);
assign A9fnv6 = (M8fnv6 & T8fnv6);
assign T8fnv6 = (Rbk7z6[3] ? Cafnv6 : V9fnv6);
assign Cafnv6 = (H9fnv6 & Jafnv6);
assign Jafnv6 = (~(Qafnv6 & Xafnv6));
assign Qafnv6 = (Rbk7z6[2] & Rbk7z6[1]);
assign H9fnv6 = (Rbk7z6[5] ? Lbfnv6 : Ebfnv6);
assign Lbfnv6 = (!Sbfnv6);
assign Sbfnv6 = (Rbk7z6[4] ? Gcfnv6 : Zbfnv6);
assign Ebfnv6 = (~(Ncfnv6 & Rbk7z6[4]));
assign M8fnv6 = (Rbk7z6[3] ? V9fnv6 : O9fnv6);
assign V9fnv6 = (Rbk7z6[5] ? Bdfnv6 : Ucfnv6);
assign Bdfnv6 = (!Idfnv6);
assign Idfnv6 = (Rbk7z6[4] ? Ncfnv6 : Gcfnv6);
assign Ucfnv6 = (~(Zbfnv6 & Rbk7z6[4]));
assign O9fnv6 = (Rbk7z6[5] ? Wdfnv6 : Pdfnv6);
assign Wdfnv6 = (!Defnv6);
assign Defnv6 = (Rbk7z6[4] ? Zbfnv6 : Ncfnv6);
assign Zbfnv6 = (Rbk7z6[2] & Kefnv6);
assign Kefnv6 = (!Rbk7z6[1]);
assign Ncfnv6 = (Rbk7z6[1] & Refnv6);
assign Pdfnv6 = (~(Rbk7z6[4] & Gcfnv6));
assign Gcfnv6 = (Rbk7z6[1] ^ Refnv6);
assign Refnv6 = (!Rbk7z6[2]);
assign N3k7z6[9] = (Obo7v6 & Cmm7z6[9]);
assign N3k7z6[8] = (Obo7v6 & Cmm7z6[8]);
assign N3k7z6[7] = (Obo7v6 & Cmm7z6[7]);
assign N3k7z6[6] = (Obo7v6 & Cmm7z6[6]);
assign N3k7z6[5] = (Cmm7z6[5] & Obo7v6);
assign N3k7z6[4] = (Cmm7z6[4] & Obo7v6);
assign N3k7z6[3] = (Cmm7z6[3] & Obo7v6);
assign N3k7z6[31] = (Obo7v6 & Cmm7z6[31]);
assign N3k7z6[30] = (Obo7v6 & Cmm7z6[30]);
assign N3k7z6[2] = (Yefnv6 & Obo7v6);
assign N3k7z6[29] = (Obo7v6 & Cmm7z6[29]);
assign N3k7z6[28] = (Obo7v6 & Cmm7z6[28]);
assign N3k7z6[27] = (Obo7v6 & Cmm7z6[27]);
assign N3k7z6[26] = (Obo7v6 & Cmm7z6[26]);
assign N3k7z6[25] = (Obo7v6 & Cmm7z6[25]);
assign N3k7z6[24] = (Obo7v6 & Cmm7z6[24]);
assign N3k7z6[23] = (Obo7v6 & Cmm7z6[23]);
assign N3k7z6[22] = (Obo7v6 & Cmm7z6[22]);
assign N3k7z6[21] = (Obo7v6 & Cmm7z6[21]);
assign N3k7z6[20] = (Obo7v6 & Cmm7z6[20]);
assign N3k7z6[19] = (Obo7v6 & Cmm7z6[19]);
assign N3k7z6[18] = (Obo7v6 & Cmm7z6[18]);
assign N3k7z6[17] = (Obo7v6 & Cmm7z6[17]);
assign N3k7z6[16] = (Obo7v6 & Cmm7z6[16]);
assign N3k7z6[15] = (Obo7v6 & Cmm7z6[15]);
assign N3k7z6[14] = (Obo7v6 & Cmm7z6[14]);
assign N3k7z6[13] = (Obo7v6 & Cmm7z6[13]);
assign N3k7z6[12] = (Obo7v6 & Cmm7z6[12]);
assign N3k7z6[11] = (Obo7v6 & Cmm7z6[11]);
assign N3k7z6[10] = (Obo7v6 & Cmm7z6[10]);
assign D847v6 = (~(Fffnv6 & Mffnv6));
assign Mffnv6 = (Tffnv6 & Agfnv6);
assign Agfnv6 = (~(Hgfnv6 & R8s7z6[0]));
assign Hgfnv6 = (Ogfnv6 & Fho7v6);
assign Ogfnv6 = (Vgfnv6 | R8s7z6[1]);
assign Tffnv6 = (~(Chfnv6 & Jhfnv6));
assign Jhfnv6 = (~(Qhfnv6 & Xhfnv6));
assign Chfnv6 = (~(Eifnv6 | Lifnv6));
assign Fffnv6 = (Sifnv6 & Zifnv6);
assign Zifnv6 = (Gjfnv6 | Ak77z6);
assign Coo7z6[9] = (Zy1ft6 & HADDRI[9]);
assign Coo7z6[8] = (Zy1ft6 & HADDRI[8]);
assign Coo7z6[7] = (Zy1ft6 & HADDRI[7]);
assign Coo7z6[6] = (Zy1ft6 & HADDRI[6]);
assign Coo7z6[5] = (Zy1ft6 & HADDRI[5]);
assign Coo7z6[4] = (Zy1ft6 & HADDRI[4]);
assign Coo7z6[3] = (Zy1ft6 & HADDRI[3]);
assign Coo7z6[31] = (Zy1ft6 & Njfnv6);
assign Coo7z6[30] = (Zy1ft6 & Ujfnv6);
assign Coo7z6[2] = (Zy1ft6 & HADDRI[2]);
assign Coo7z6[29] = (Zy1ft6 & Bkfnv6);
assign Coo7z6[28] = (Zy1ft6 & HADDRI[28]);
assign Coo7z6[27] = (Zy1ft6 & HADDRI[27]);
assign Coo7z6[26] = (Zy1ft6 & HADDRI[26]);
assign Coo7z6[25] = (Zy1ft6 & HADDRI[25]);
assign Coo7z6[24] = (Zy1ft6 & HADDRI[24]);
assign Coo7z6[23] = (Zy1ft6 & HADDRI[23]);
assign Coo7z6[22] = (Zy1ft6 & HADDRI[22]);
assign Coo7z6[21] = (Zy1ft6 & HADDRI[21]);
assign Coo7z6[20] = (Zy1ft6 & HADDRI[20]);
assign Coo7z6[19] = (Zy1ft6 & HADDRI[19]);
assign Coo7z6[18] = (Zy1ft6 & HADDRI[18]);
assign Coo7z6[17] = (Zy1ft6 & HADDRI[17]);
assign Coo7z6[16] = (Zy1ft6 & HADDRI[16]);
assign Coo7z6[15] = (Zy1ft6 & HADDRI[15]);
assign Coo7z6[14] = (Zy1ft6 & HADDRI[14]);
assign Coo7z6[13] = (Zy1ft6 & HADDRI[13]);
assign Coo7z6[12] = (Zy1ft6 & HADDRI[12]);
assign Coo7z6[11] = (Zy1ft6 & HADDRI[11]);
assign Coo7z6[10] = (Zy1ft6 & HADDRI[10]);
assign Zmo7z6[9] = (Zy1ft6 & Cmm7z6[9]);
assign Zmo7z6[8] = (Zy1ft6 & Cmm7z6[8]);
assign Zmo7z6[7] = (Zy1ft6 & Cmm7z6[7]);
assign Zmo7z6[6] = (Zy1ft6 & Cmm7z6[6]);
assign Zmo7z6[5] = (Zy1ft6 & Cmm7z6[5]);
assign Zmo7z6[4] = (Zy1ft6 & Cmm7z6[4]);
assign Zmo7z6[3] = (Zy1ft6 & Cmm7z6[3]);
assign Zmo7z6[31] = (Zy1ft6 & Cmm7z6[31]);
assign Zmo7z6[30] = (Zy1ft6 & Cmm7z6[30]);
assign Zmo7z6[2] = (Zy1ft6 & Yefnv6);
assign Zmo7z6[29] = (Zy1ft6 & Cmm7z6[29]);
assign Zmo7z6[28] = (Zy1ft6 & Cmm7z6[28]);
assign Zmo7z6[27] = (Zy1ft6 & Cmm7z6[27]);
assign Zmo7z6[26] = (Zy1ft6 & Cmm7z6[26]);
assign Zmo7z6[25] = (Zy1ft6 & Cmm7z6[25]);
assign Zmo7z6[24] = (Zy1ft6 & Cmm7z6[24]);
assign Zmo7z6[23] = (Zy1ft6 & Cmm7z6[23]);
assign Zmo7z6[22] = (Zy1ft6 & Cmm7z6[22]);
assign Zmo7z6[21] = (Zy1ft6 & Cmm7z6[21]);
assign Zmo7z6[20] = (Zy1ft6 & Cmm7z6[20]);
assign Zmo7z6[19] = (Zy1ft6 & Cmm7z6[19]);
assign Zmo7z6[18] = (Zy1ft6 & Cmm7z6[18]);
assign Zmo7z6[17] = (Zy1ft6 & Cmm7z6[17]);
assign Zmo7z6[16] = (Zy1ft6 & Cmm7z6[16]);
assign Zmo7z6[15] = (Zy1ft6 & Cmm7z6[15]);
assign Zmo7z6[14] = (Zy1ft6 & Cmm7z6[14]);
assign Zmo7z6[13] = (Zy1ft6 & Cmm7z6[13]);
assign Zmo7z6[12] = (Zy1ft6 & Cmm7z6[12]);
assign Zmo7z6[11] = (Zy1ft6 & Cmm7z6[11]);
assign Zmo7z6[10] = (Zy1ft6 & Cmm7z6[10]);
assign T6r7z6[9] = (Ikfnv6 & Pkfnv6);
assign T6r7z6[8] = (Wkfnv6 & Dlfnv6);
assign T6r7z6[7] = (Klfnv6 & Rlfnv6);
assign T6r7z6[6] = (Ylfnv6 & Fmfnv6);
assign T6r7z6[5] = (Mmfnv6 & Tmfnv6);
assign T6r7z6[4] = (Anfnv6 & Hnfnv6);
assign T6r7z6[3] = (Onfnv6 & Vnfnv6);
assign T6r7z6[31] = (Um77z6 & HTMDHBURST[0]);
assign T6r7z6[30] = (Cn77z6 & HTMDHBURST[0]);
assign T6r7z6[2] = (Cofnv6 & Jofnv6);
assign T6r7z6[29] = (Kn77z6 & HTMDHBURST[0]);
assign T6r7z6[28] = (Sn77z6 & HTMDHBURST[0]);
assign T6r7z6[27] = (Ao77z6 & HTMDHBURST[0]);
assign T6r7z6[26] = (Io77z6 & HTMDHBURST[0]);
assign T6r7z6[25] = (Qo77z6 & HTMDHBURST[0]);
assign T6r7z6[24] = (Yo77z6 & HTMDHBURST[0]);
assign T6r7z6[23] = (Gp77z6 & HTMDHBURST[0]);
assign T6r7z6[22] = (Op77z6 & HTMDHBURST[0]);
assign T6r7z6[21] = (Wp77z6 & HTMDHBURST[0]);
assign T6r7z6[20] = (Eq77z6 & HTMDHBURST[0]);
assign T6r7z6[1] = (Qofnv6 & Xofnv6);
assign T6r7z6[19] = (Mq77z6 & HTMDHBURST[0]);
assign T6r7z6[18] = (Uq77z6 & HTMDHBURST[0]);
assign T6r7z6[17] = (Cr77z6 & HTMDHBURST[0]);
assign T6r7z6[16] = (Kr77z6 & HTMDHBURST[0]);
assign T6r7z6[14] = (Epfnv6 & Lpfnv6);
assign T6r7z6[13] = (Spfnv6 & Zpfnv6);
assign T6r7z6[12] = (Gqfnv6 & Nqfnv6);
assign T6r7z6[11] = (Uqfnv6 & Brfnv6);
assign T6r7z6[10] = (~(Irfnv6 | Prfnv6));
assign S8r7z6[9] = (Mkp7z6[9] & Pkfnv6);
assign S8r7z6[8] = (Mkp7z6[8] & Dlfnv6);
assign S8r7z6[7] = (Mkp7z6[7] & Rlfnv6);
assign S8r7z6[6] = (Mkp7z6[6] & Fmfnv6);
assign S8r7z6[5] = (Mkp7z6[5] & Tmfnv6);
assign S8r7z6[4] = (Mkp7z6[4] & Hnfnv6);
assign S8r7z6[3] = (Mkp7z6[3] & Onfnv6);
assign S8r7z6[2] = (Mkp7z6[2] & Jofnv6);
assign S8r7z6[14] = (Mkp7z6[14] & Lpfnv6);
assign S8r7z6[13] = (Mkp7z6[13] & Zpfnv6);
assign S8r7z6[12] = (Mkp7z6[12] & Nqfnv6);
assign S8r7z6[11] = (Mkp7z6[11] & Brfnv6);
assign S8r7z6[10] = (Mkp7z6[10] & Wrfnv6);
assign Sar7z6[9] = (Dsfnv6 & Pkfnv6);
assign Sar7z6[8] = (Ksfnv6 & Dlfnv6);
assign Sar7z6[7] = (Rsfnv6 & Rlfnv6);
assign Sar7z6[6] = (Ysfnv6 & Fmfnv6);
assign Fmfnv6 = (Tmfnv6 | Ftfnv6);
assign Ftfnv6 = (Mtfnv6 & Rlfnv6);
assign Sar7z6[5] = (Ttfnv6 & Tmfnv6);
assign Tmfnv6 = (Hnfnv6 | Aufnv6);
assign Aufnv6 = (~(Rip7z6[3] | Rip7z6[1]));
assign Sar7z6[4] = (Hufnv6 & Hnfnv6);
assign Hnfnv6 = (Onfnv6 | Oufnv6);
assign Oufnv6 = (Vufnv6 & Mtfnv6);
assign Vufnv6 = (Cvfnv6 & Rlfnv6);
assign Rlfnv6 = (!Rip7z6[3]);
assign Sar7z6[3] = (Jvfnv6 & Onfnv6);
assign Sar7z6[2] = (Qvfnv6 & Jofnv6);
assign Jofnv6 = (~(Xvfnv6 & Ewfnv6));
assign Ewfnv6 = (~(Onfnv6 & Mtfnv6));
assign Xvfnv6 = (!Qofnv6);
assign Sar7z6[1] = (~(Lwfnv6 & Swfnv6));
assign Swfnv6 = (~(S8r7z6[1] & Zwfnv6));
assign S8r7z6[1] = (Mkp7z6[1] & Qofnv6);
assign Lwfnv6 = (~(Gxfnv6 & Qofnv6));
assign Sar7z6[14] = (Nxfnv6 & Lpfnv6);
assign Lpfnv6 = (Mtfnv6 | Zpfnv6);
assign Sar7z6[13] = (Uxfnv6 & Zpfnv6);
assign Zpfnv6 = (Cvfnv6 | Nqfnv6);
assign Sar7z6[12] = (Byfnv6 & Nqfnv6);
assign Nqfnv6 = (Brfnv6 | Iyfnv6);
assign Iyfnv6 = (Mtfnv6 & Cvfnv6);
assign Sar7z6[11] = (Pyfnv6 & Brfnv6);
assign Brfnv6 = (~(Rip7z6[2] & Prfnv6));
assign Prfnv6 = (!Wrfnv6);
assign Sar7z6[10] = (Wyfnv6 & Wrfnv6);
assign Wrfnv6 = (Pkfnv6 | Dzfnv6);
assign Dzfnv6 = (~(Rip7z6[0] | Rip7z6[2]));
assign Pkfnv6 = (Dlfnv6 | Kzfnv6);
assign Dlfnv6 = (~(Rip7z6[3] & Rzfnv6));
assign Rzfnv6 = (~(Kzfnv6 & Mtfnv6));
assign Kzfnv6 = (~(Rip7z6[2] | Rip7z6[1]));
assign Sar7z6[0] = (Zwfnv6 ? S8r7z6[0] : Yzfnv6);
assign Zwfnv6 = (F0gnv6 & M0gnv6);
assign M0gnv6 = (~(T0gnv6 & A1gnv6));
assign A1gnv6 = (~(Mkp7z6[1] & H1gnv6));
assign F0gnv6 = (~(O1gnv6 | V1gnv6));
assign O1gnv6 = (C2gnv6 & J2gnv6);
assign J2gnv6 = (~(Q2gnv6 & X2gnv6));
assign X2gnv6 = (~(Mkp7z6[1] & E3gnv6));
assign E3gnv6 = (L3gnv6 | Mkp7z6[0]);
assign S8r7z6[0] = (S3gnv6 & Mkp7z6[0]);
assign Yzfnv6 = (S3gnv6 & Z3gnv6);
assign S3gnv6 = (Qofnv6 & Mtfnv6);
assign Mtfnv6 = (!Rip7z6[0]);
assign Qofnv6 = (Onfnv6 & Cvfnv6);
assign Cvfnv6 = (!Rip7z6[1]);
assign Onfnv6 = (~(Rip7z6[2] | Rip7z6[3]));
assign Ve5ft6 = (Sr77z6 & HTMDHBURST[0]);
assign P0r7z6[9] = (Ikfnv6 & G4gnv6);
assign P0r7z6[8] = (Wkfnv6 & N4gnv6);
assign P0r7z6[7] = (Klfnv6 & U4gnv6);
assign P0r7z6[6] = (Ylfnv6 & B5gnv6);
assign P0r7z6[5] = (Mmfnv6 & I5gnv6);
assign P0r7z6[4] = (Anfnv6 & P5gnv6);
assign P0r7z6[3] = (W5gnv6 & Vnfnv6);
assign P0r7z6[2] = (Cofnv6 & D6gnv6);
assign P0r7z6[1] = (K6gnv6 & Xofnv6);
assign P0r7z6[14] = (Epfnv6 & R6gnv6);
assign P0r7z6[13] = (Spfnv6 & Y6gnv6);
assign P0r7z6[12] = (Gqfnv6 & F7gnv6);
assign P0r7z6[11] = (Uqfnv6 & M7gnv6);
assign P0r7z6[10] = (~(Irfnv6 | T7gnv6));
assign O2r7z6[9] = (Bqp7z6[9] & G4gnv6);
assign O2r7z6[8] = (Bqp7z6[8] & N4gnv6);
assign O2r7z6[7] = (Bqp7z6[7] & U4gnv6);
assign O2r7z6[6] = (Bqp7z6[6] & B5gnv6);
assign O2r7z6[5] = (Bqp7z6[5] & I5gnv6);
assign O2r7z6[4] = (Bqp7z6[4] & P5gnv6);
assign O2r7z6[3] = (Bqp7z6[3] & W5gnv6);
assign O2r7z6[2] = (Bqp7z6[2] & D6gnv6);
assign O2r7z6[14] = (Bqp7z6[14] & R6gnv6);
assign O2r7z6[13] = (Bqp7z6[13] & Y6gnv6);
assign O2r7z6[12] = (Bqp7z6[12] & F7gnv6);
assign O2r7z6[11] = (Bqp7z6[11] & M7gnv6);
assign O2r7z6[10] = (Bqp7z6[10] & A8gnv6);
assign O4r7z6[9] = (Dsfnv6 & G4gnv6);
assign O4r7z6[8] = (Ksfnv6 & N4gnv6);
assign O4r7z6[7] = (Rsfnv6 & U4gnv6);
assign O4r7z6[6] = (Ysfnv6 & B5gnv6);
assign B5gnv6 = (I5gnv6 | H8gnv6);
assign H8gnv6 = (O8gnv6 & U4gnv6);
assign O4r7z6[5] = (Ttfnv6 & I5gnv6);
assign I5gnv6 = (P5gnv6 | V8gnv6);
assign V8gnv6 = (~(Gop7z6[3] | Gop7z6[1]));
assign O4r7z6[4] = (Hufnv6 & P5gnv6);
assign P5gnv6 = (W5gnv6 | C9gnv6);
assign C9gnv6 = (J9gnv6 & O8gnv6);
assign J9gnv6 = (Q9gnv6 & U4gnv6);
assign U4gnv6 = (!Gop7z6[3]);
assign O4r7z6[3] = (W5gnv6 & Jvfnv6);
assign O4r7z6[2] = (Qvfnv6 & D6gnv6);
assign D6gnv6 = (~(X9gnv6 & Eagnv6));
assign Eagnv6 = (~(W5gnv6 & O8gnv6));
assign X9gnv6 = (!K6gnv6);
assign O4r7z6[1] = (~(Lagnv6 & Sagnv6));
assign Sagnv6 = (~(O2r7z6[1] & Zagnv6));
assign O2r7z6[1] = (Bqp7z6[1] & K6gnv6);
assign Lagnv6 = (~(K6gnv6 & Gxfnv6));
assign O4r7z6[14] = (Nxfnv6 & R6gnv6);
assign R6gnv6 = (O8gnv6 | Y6gnv6);
assign O4r7z6[13] = (Uxfnv6 & Y6gnv6);
assign Y6gnv6 = (Q9gnv6 | F7gnv6);
assign O4r7z6[12] = (Byfnv6 & F7gnv6);
assign F7gnv6 = (M7gnv6 | Gbgnv6);
assign Gbgnv6 = (~(Gop7z6[0] | Gop7z6[1]));
assign O4r7z6[11] = (Pyfnv6 & M7gnv6);
assign M7gnv6 = (~(Gop7z6[2] & T7gnv6));
assign T7gnv6 = (!A8gnv6);
assign O4r7z6[10] = (Wyfnv6 & A8gnv6);
assign A8gnv6 = (G4gnv6 | Nbgnv6);
assign Nbgnv6 = (~(Gop7z6[0] | Gop7z6[2]));
assign G4gnv6 = (N4gnv6 | Ubgnv6);
assign N4gnv6 = (~(Gop7z6[3] & Bcgnv6));
assign Bcgnv6 = (~(Ubgnv6 & O8gnv6));
assign Ubgnv6 = (~(Gop7z6[2] | Gop7z6[1]));
assign O4r7z6[0] = (Zagnv6 ? O2r7z6[0] : Icgnv6);
assign Zagnv6 = (Pcgnv6 & Wcgnv6);
assign Wcgnv6 = (~(T0gnv6 & Ddgnv6));
assign Ddgnv6 = (~(Bqp7z6[1] & H1gnv6));
assign Pcgnv6 = (~(Kdgnv6 | Rdgnv6));
assign Kdgnv6 = (C2gnv6 & Ydgnv6);
assign Ydgnv6 = (~(Q2gnv6 & Fegnv6));
assign Fegnv6 = (~(Bqp7z6[1] & Megnv6));
assign Megnv6 = (L3gnv6 | Bqp7z6[0]);
assign O2r7z6[0] = (Tegnv6 & Bqp7z6[0]);
assign Tegnv6 = (K6gnv6 & O8gnv6);
assign Icgnv6 = (Afgnv6 & K6gnv6);
assign K6gnv6 = (W5gnv6 & Q9gnv6);
assign Q9gnv6 = (!Gop7z6[1]);
assign W5gnv6 = (~(Gop7z6[2] | Gop7z6[3]));
assign Afgnv6 = (Z3gnv6 & O8gnv6);
assign O8gnv6 = (!Gop7z6[0]);
assign Luq7z6[9] = (Ikfnv6 & Hfgnv6);
assign Luq7z6[8] = (Wkfnv6 & Ofgnv6);
assign Luq7z6[7] = (Klfnv6 & Vfgnv6);
assign Luq7z6[6] = (Ylfnv6 & Cggnv6);
assign Luq7z6[5] = (Mmfnv6 & Jggnv6);
assign Luq7z6[4] = (Anfnv6 & Qggnv6);
assign Luq7z6[3] = (Xggnv6 & Vnfnv6);
assign Luq7z6[2] = (Cofnv6 & Ehgnv6);
assign Luq7z6[1] = (Lhgnv6 & Xofnv6);
assign Luq7z6[14] = (Epfnv6 & Shgnv6);
assign Luq7z6[13] = (Spfnv6 & Zhgnv6);
assign Luq7z6[12] = (Gqfnv6 & Gignv6);
assign Luq7z6[11] = (Uqfnv6 & Nignv6);
assign Luq7z6[10] = (~(Irfnv6 | Uignv6));
assign Kwq7z6[9] = (B2q7z6[9] & Hfgnv6);
assign Kwq7z6[8] = (B2q7z6[8] & Ofgnv6);
assign Kwq7z6[7] = (B2q7z6[7] & Vfgnv6);
assign Kwq7z6[6] = (B2q7z6[6] & Cggnv6);
assign Kwq7z6[5] = (B2q7z6[5] & Jggnv6);
assign Kwq7z6[4] = (B2q7z6[4] & Qggnv6);
assign Kwq7z6[3] = (B2q7z6[3] & Xggnv6);
assign Kwq7z6[2] = (B2q7z6[2] & Ehgnv6);
assign Kwq7z6[14] = (B2q7z6[14] & Shgnv6);
assign Kwq7z6[13] = (B2q7z6[13] & Zhgnv6);
assign Kwq7z6[12] = (B2q7z6[12] & Gignv6);
assign Kwq7z6[11] = (B2q7z6[11] & Nignv6);
assign Kwq7z6[10] = (B2q7z6[10] & Bjgnv6);
assign Kyq7z6[9] = (Dsfnv6 & Hfgnv6);
assign Kyq7z6[8] = (Ksfnv6 & Ofgnv6);
assign Kyq7z6[7] = (Rsfnv6 & Vfgnv6);
assign Kyq7z6[6] = (Ysfnv6 & Cggnv6);
assign Cggnv6 = (Jggnv6 | Ijgnv6);
assign Ijgnv6 = (Pjgnv6 & Vfgnv6);
assign Kyq7z6[5] = (Ttfnv6 & Jggnv6);
assign Jggnv6 = (Qggnv6 | Wjgnv6);
assign Wjgnv6 = (~(G0q7z6[1] | G0q7z6[3]));
assign Kyq7z6[4] = (Hufnv6 & Qggnv6);
assign Qggnv6 = (Xggnv6 | Dkgnv6);
assign Dkgnv6 = (Kkgnv6 & Pjgnv6);
assign Kkgnv6 = (Rkgnv6 & Vfgnv6);
assign Vfgnv6 = (!G0q7z6[3]);
assign Kyq7z6[3] = (Xggnv6 & Jvfnv6);
assign Kyq7z6[2] = (Qvfnv6 & Ehgnv6);
assign Ehgnv6 = (~(Ykgnv6 & Flgnv6));
assign Flgnv6 = (~(Xggnv6 & Pjgnv6));
assign Ykgnv6 = (!Lhgnv6);
assign Kyq7z6[1] = (~(Mlgnv6 & Tlgnv6));
assign Tlgnv6 = (~(Kwq7z6[1] & Amgnv6));
assign Kwq7z6[1] = (B2q7z6[1] & Lhgnv6);
assign Mlgnv6 = (~(Lhgnv6 & Gxfnv6));
assign Kyq7z6[14] = (Nxfnv6 & Shgnv6);
assign Shgnv6 = (Pjgnv6 | Zhgnv6);
assign Kyq7z6[13] = (Uxfnv6 & Zhgnv6);
assign Zhgnv6 = (Rkgnv6 | Gignv6);
assign Kyq7z6[12] = (Byfnv6 & Gignv6);
assign Gignv6 = (Nignv6 | Hmgnv6);
assign Hmgnv6 = (Pjgnv6 & Rkgnv6);
assign Kyq7z6[11] = (Pyfnv6 & Nignv6);
assign Nignv6 = (~(G0q7z6[2] & Uignv6));
assign Uignv6 = (!Bjgnv6);
assign Kyq7z6[10] = (Wyfnv6 & Bjgnv6);
assign Bjgnv6 = (Hfgnv6 | Omgnv6);
assign Omgnv6 = (~(G0q7z6[0] | G0q7z6[2]));
assign Hfgnv6 = (~(Vmgnv6 & Cngnv6));
assign Cngnv6 = (G0q7z6[1] | G0q7z6[2]);
assign Vmgnv6 = (!Ofgnv6);
assign Ofgnv6 = (~(G0q7z6[3] & Jngnv6));
assign Jngnv6 = (~(Qngnv6 & Pjgnv6));
assign Qngnv6 = (~(G0q7z6[1] | G0q7z6[2]));
assign Kyq7z6[0] = (Amgnv6 ? Kwq7z6[0] : Xngnv6);
assign Amgnv6 = (Eognv6 & Lognv6);
assign Lognv6 = (~(T0gnv6 & Sognv6));
assign Sognv6 = (~(B2q7z6[1] & H1gnv6));
assign Eognv6 = (~(Zognv6 | Gpgnv6));
assign Zognv6 = (C2gnv6 & Npgnv6);
assign Npgnv6 = (~(Q2gnv6 & Upgnv6));
assign Upgnv6 = (~(B2q7z6[1] & Bqgnv6));
assign Bqgnv6 = (L3gnv6 | B2q7z6[0]);
assign Kwq7z6[0] = (Iqgnv6 & B2q7z6[0]);
assign Iqgnv6 = (Lhgnv6 & Pjgnv6);
assign Xngnv6 = (Pqgnv6 & Lhgnv6);
assign Lhgnv6 = (Xggnv6 & Rkgnv6);
assign Rkgnv6 = (!G0q7z6[1]);
assign Xggnv6 = (~(G0q7z6[2] | G0q7z6[3]));
assign Pqgnv6 = (Z3gnv6 & Pjgnv6);
assign Pjgnv6 = (!G0q7z6[0]);
assign Hoq7z6[9] = (Ikfnv6 & Wqgnv6);
assign Ikfnv6 = (Ot77z6 & HTMDHBURST[0]);
assign Hoq7z6[8] = (Wkfnv6 & Drgnv6);
assign Wkfnv6 = (Wt77z6 & HTMDHBURST[0]);
assign Hoq7z6[7] = (Klfnv6 & Krgnv6);
assign Klfnv6 = (Eu77z6 & HTMDHBURST[0]);
assign Hoq7z6[6] = (Ylfnv6 & Rrgnv6);
assign Ylfnv6 = (Mu77z6 & HTMDHBURST[0]);
assign Hoq7z6[5] = (Mmfnv6 & Yrgnv6);
assign Mmfnv6 = (Uu77z6 & HTMDHBURST[0]);
assign Hoq7z6[4] = (Anfnv6 & Fsgnv6);
assign Anfnv6 = (Cv77z6 & HTMDHBURST[0]);
assign Hoq7z6[3] = (Msgnv6 & Vnfnv6);
assign Vnfnv6 = (Kv77z6 & HTMDHBURST[0]);
assign Hoq7z6[2] = (Cofnv6 & Tsgnv6);
assign Cofnv6 = (Sv77z6 & HTMDHBURST[0]);
assign Hoq7z6[1] = (Atgnv6 & Xofnv6);
assign Xofnv6 = (Aw77z6 & HTMDHBURST[0]);
assign Hoq7z6[14] = (Epfnv6 & Htgnv6);
assign Epfnv6 = (As77z6 & HTMDHBURST[0]);
assign Hoq7z6[13] = (Spfnv6 & Otgnv6);
assign Spfnv6 = (Is77z6 & HTMDHBURST[0]);
assign Hoq7z6[12] = (Gqfnv6 & Vtgnv6);
assign Gqfnv6 = (Qs77z6 & HTMDHBURST[0]);
assign Hoq7z6[11] = (Uqfnv6 & Cugnv6);
assign Uqfnv6 = (Ys77z6 & HTMDHBURST[0]);
assign Hoq7z6[10] = (~(Irfnv6 | Jugnv6));
assign Irfnv6 = (~(Gt77z6 & HTMDHBURST[0]));
assign Gqq7z6[9] = (E6p7z6[9] & Wqgnv6);
assign Gqq7z6[8] = (E6p7z6[8] & Drgnv6);
assign Gqq7z6[7] = (E6p7z6[7] & Krgnv6);
assign Gqq7z6[6] = (E6p7z6[6] & Rrgnv6);
assign Gqq7z6[5] = (E6p7z6[5] & Yrgnv6);
assign Gqq7z6[4] = (E6p7z6[4] & Fsgnv6);
assign Gqq7z6[3] = (E6p7z6[3] & Msgnv6);
assign Gqq7z6[2] = (E6p7z6[2] & Tsgnv6);
assign Gqq7z6[14] = (E6p7z6[14] & Htgnv6);
assign Gqq7z6[13] = (E6p7z6[13] & Otgnv6);
assign Gqq7z6[12] = (E6p7z6[12] & Vtgnv6);
assign Gqq7z6[11] = (E6p7z6[11] & Cugnv6);
assign Gqq7z6[10] = (E6p7z6[10] & Qugnv6);
assign Gsq7z6[9] = (Xugnv6 & Wqgnv6);
assign Xugnv6 = (W22ft6 ? U9p7z6[9] : Dsfnv6);
assign Gsq7z6[8] = (Evgnv6 & Drgnv6);
assign Evgnv6 = (W22ft6 ? U9p7z6[8] : Ksfnv6);
assign Gsq7z6[7] = (Lvgnv6 & Krgnv6);
assign Lvgnv6 = (W22ft6 ? U9p7z6[7] : Rsfnv6);
assign Gsq7z6[6] = (Svgnv6 & Rrgnv6);
assign Rrgnv6 = (Yrgnv6 | Zvgnv6);
assign Zvgnv6 = (Gwgnv6 & Krgnv6);
assign Svgnv6 = (W22ft6 ? U9p7z6[6] : Ysfnv6);
assign Gsq7z6[5] = (Nwgnv6 & Yrgnv6);
assign Yrgnv6 = (Fsgnv6 | Uwgnv6);
assign Uwgnv6 = (~(Q8p7z6[1] | Q8p7z6[3]));
assign Nwgnv6 = (W22ft6 ? U9p7z6[5] : Ttfnv6);
assign Gsq7z6[4] = (Bxgnv6 & Fsgnv6);
assign Fsgnv6 = (Msgnv6 | Ixgnv6);
assign Ixgnv6 = (Pxgnv6 & Gwgnv6);
assign Pxgnv6 = (Wxgnv6 & Krgnv6);
assign Krgnv6 = (!Q8p7z6[3]);
assign Bxgnv6 = (W22ft6 ? U9p7z6[4] : Hufnv6);
assign Gsq7z6[3] = (Dygnv6 & Msgnv6);
assign Dygnv6 = (W22ft6 ? U9p7z6[3] : Jvfnv6);
assign Gsq7z6[31] = (W22ft6 ? U9p7z6[31] : Sar7z6[31]);
assign Sar7z6[31] = (~(Kygnv6 | Rygnv6));
assign Gsq7z6[30] = (W22ft6 ? U9p7z6[30] : Sar7z6[30]);
assign Sar7z6[30] = (~(Kygnv6 | Yygnv6));
assign Gsq7z6[2] = (Fzgnv6 & Tsgnv6);
assign Tsgnv6 = (~(Mzgnv6 & Tzgnv6));
assign Tzgnv6 = (~(Msgnv6 & Gwgnv6));
assign Mzgnv6 = (!Atgnv6);
assign Fzgnv6 = (W22ft6 ? U9p7z6[2] : Qvfnv6);
assign Gsq7z6[29] = (W22ft6 ? U9p7z6[29] : Sar7z6[29]);
assign Sar7z6[29] = (~(Kygnv6 | A0hnv6));
assign Gsq7z6[28] = (W22ft6 ? U9p7z6[28] : Sar7z6[28]);
assign Sar7z6[28] = (~(Kygnv6 | H0hnv6));
assign Gsq7z6[27] = (W22ft6 ? U9p7z6[27] : Sar7z6[27]);
assign Sar7z6[27] = (~(Kygnv6 | O0hnv6));
assign Gsq7z6[26] = (W22ft6 ? U9p7z6[26] : Sar7z6[26]);
assign Sar7z6[26] = (~(Kygnv6 | V0hnv6));
assign Gsq7z6[25] = (W22ft6 ? U9p7z6[25] : Sar7z6[25]);
assign Sar7z6[25] = (~(Kygnv6 | C1hnv6));
assign Gsq7z6[24] = (W22ft6 ? U9p7z6[24] : Sar7z6[24]);
assign Sar7z6[24] = (~(Kygnv6 | J1hnv6));
assign Gsq7z6[23] = (W22ft6 ? U9p7z6[23] : Sar7z6[23]);
assign Sar7z6[23] = (~(Kygnv6 | Q1hnv6));
assign Gsq7z6[22] = (W22ft6 ? U9p7z6[22] : Sar7z6[22]);
assign Sar7z6[22] = (~(Kygnv6 | X1hnv6));
assign Gsq7z6[21] = (W22ft6 ? U9p7z6[21] : Sar7z6[21]);
assign Sar7z6[21] = (~(Kygnv6 | E2hnv6));
assign Gsq7z6[20] = (W22ft6 ? U9p7z6[20] : Sar7z6[20]);
assign Sar7z6[20] = (~(Kygnv6 | L2hnv6));
assign Gsq7z6[1] = (~(S2hnv6 & Z2hnv6));
assign Z2hnv6 = (~(G3hnv6 & Atgnv6));
assign G3hnv6 = (W22ft6 ? U9p7z6[1] : Gxfnv6);
assign S2hnv6 = (~(Gqq7z6[1] & N3hnv6));
assign Gqq7z6[1] = (E6p7z6[1] & Atgnv6);
assign Gsq7z6[19] = (W22ft6 ? U9p7z6[19] : Sar7z6[19]);
assign Sar7z6[19] = (~(Kygnv6 | U3hnv6));
assign U3hnv6 = (!Cmm7z6[19]);
assign Gsq7z6[18] = (W22ft6 ? U9p7z6[18] : Sar7z6[18]);
assign Sar7z6[18] = (~(Kygnv6 | B4hnv6));
assign B4hnv6 = (!Cmm7z6[18]);
assign Gsq7z6[17] = (W22ft6 ? U9p7z6[17] : Sar7z6[17]);
assign Sar7z6[17] = (~(Kygnv6 | I4hnv6));
assign Gsq7z6[16] = (W22ft6 ? U9p7z6[16] : Sar7z6[16]);
assign Sar7z6[16] = (~(Kygnv6 | P4hnv6));
assign Gsq7z6[14] = (W4hnv6 & Htgnv6);
assign Htgnv6 = (Gwgnv6 | Otgnv6);
assign W4hnv6 = (W22ft6 ? U9p7z6[14] : Nxfnv6);
assign Gsq7z6[13] = (D5hnv6 & Otgnv6);
assign Otgnv6 = (Wxgnv6 | Vtgnv6);
assign D5hnv6 = (W22ft6 ? U9p7z6[13] : Uxfnv6);
assign Gsq7z6[12] = (K5hnv6 & Vtgnv6);
assign Vtgnv6 = (Cugnv6 | R5hnv6);
assign R5hnv6 = (Gwgnv6 & Wxgnv6);
assign K5hnv6 = (W22ft6 ? U9p7z6[12] : Byfnv6);
assign Gsq7z6[11] = (Y5hnv6 & Cugnv6);
assign Cugnv6 = (~(Q8p7z6[2] & Jugnv6));
assign Jugnv6 = (!Qugnv6);
assign Y5hnv6 = (W22ft6 ? U9p7z6[11] : Pyfnv6);
assign Gsq7z6[10] = (F6hnv6 & Qugnv6);
assign Qugnv6 = (Wqgnv6 | M6hnv6);
assign M6hnv6 = (~(Q8p7z6[0] | Q8p7z6[2]));
assign Wqgnv6 = (Drgnv6 | T6hnv6);
assign Drgnv6 = (~(Q8p7z6[3] & A7hnv6));
assign A7hnv6 = (~(T6hnv6 & Gwgnv6));
assign T6hnv6 = (~(Q8p7z6[1] | Q8p7z6[2]));
assign F6hnv6 = (W22ft6 ? U9p7z6[10] : Wyfnv6);
assign Gsq7z6[0] = (~(H7hnv6 & O7hnv6));
assign O7hnv6 = (~(V7hnv6 & C8hnv6));
assign C8hnv6 = (W22ft6 ? U9p7z6[0] : J8hnv6);
assign J8hnv6 = (~(L3gnv6 | N3hnv6));
assign H7hnv6 = (~(Gqq7z6[0] & N3hnv6));
assign N3hnv6 = (Q8hnv6 & X8hnv6);
assign X8hnv6 = (~(E9hnv6 | W22ft6));
assign Q8hnv6 = (L9hnv6 & S9hnv6);
assign S9hnv6 = (~(T0gnv6 & Z9hnv6));
assign Z9hnv6 = (~(E6p7z6[1] & H1gnv6));
assign H1gnv6 = (~(Gxfnv6 & Z3gnv6));
assign T0gnv6 = (~(L3gnv6 & Gahnv6));
assign Gahnv6 = (!Gxfnv6);
assign L9hnv6 = (~(C2gnv6 & Nahnv6));
assign Nahnv6 = (~(Q2gnv6 & Uahnv6));
assign Uahnv6 = (~(E6p7z6[1] & Bbhnv6));
assign Bbhnv6 = (L3gnv6 | E6p7z6[0]);
assign L3gnv6 = (!Z3gnv6);
assign Q2gnv6 = (Ibhnv6 & Pbhnv6);
assign Ibhnv6 = (Wbhnv6 & HTMDHBURST[0]);
assign C2gnv6 = (Dchnv6 | Kygnv6);
assign Dchnv6 = (Pbhnv6 ? Kchnv6 : Wbhnv6);
assign Kchnv6 = (~(Gxfnv6 & Wbhnv6));
assign Gqq7z6[0] = (V7hnv6 & E6p7z6[0]);
assign V7hnv6 = (Atgnv6 & Gwgnv6);
assign Gwgnv6 = (!Q8p7z6[0]);
assign Atgnv6 = (Msgnv6 & Wxgnv6);
assign Wxgnv6 = (!Q8p7z6[1]);
assign Msgnv6 = (~(Q8p7z6[2] | Q8p7z6[3]));
assign Bu4ft6 = (W22ft6 ? U9p7z6[15] : Tp5ft6);
assign Zdedt6 = (~(Rchnv6 & Ychnv6));
assign Ofedt6 = (~(Fdhnv6 & Mdhnv6));
assign Dhedt6 = (~(Tdhnv6 & Aehnv6));
assign Tdhnv6 = (Rchnv6 & Hehnv6);
assign Siedt6 = (~(Oehnv6 & Vehnv6));
assign Hkedt6 = (~(Cfhnv6 & Jfhnv6));
assign Cfhnv6 = (Rchnv6 & Qfhnv6);
assign Wledt6 = (~(Fdhnv6 & Qfhnv6));
assign Lnedt6 = (~(Xfhnv6 & Jfhnv6));
assign Xfhnv6 = (Rchnv6 & Eghnv6);
assign Rchnv6 = (~(Lghnv6 | Sghnv6));
assign Apedt6 = (~(Fdhnv6 & Eghnv6));
assign Fdhnv6 = (Oehnv6 & Zghnv6);
assign Oehnv6 = (~(Ghhnv6 | Sghnv6));
assign Sghnv6 = (~(Nhhnv6 | Uhhnv6));
assign Pqedt6 = (~(Bihnv6 & Mdhnv6));
assign Esedt6 = (~(Iihnv6 & Ychnv6));
assign Ychnv6 = (Pihnv6 & Hehnv6);
assign Pihnv6 = (Mdhnv6 & Wihnv6);
assign Ttedt6 = (~(Djhnv6 & Vehnv6));
assign Vehnv6 = (Kjhnv6 & Aehnv6);
assign Kjhnv6 = (Rjhnv6 & Yjhnv6);
assign Ivedt6 = (~(Fkhnv6 & Iihnv6));
assign Fkhnv6 = (Aehnv6 & Hehnv6);
assign Hehnv6 = (Mkhnv6 & Tkhnv6);
assign Tkhnv6 = (~(Alhnv6 & Hlhnv6));
assign Mkhnv6 = (Olhnv6 & Vlhnv6);
assign Aehnv6 = (Cmhnv6 & Jmhnv6);
assign Jmhnv6 = (~(Qmhnv6 & Hlhnv6));
assign Cmhnv6 = (Uhhnv6 ? Eghnv6 : Mdhnv6);
assign Xwedt6 = (~(Bihnv6 & Qfhnv6));
assign Myedt6 = (~(Xmhnv6 & Iihnv6));
assign Xmhnv6 = (Jfhnv6 & Qfhnv6);
assign Qfhnv6 = (Uhhnv6 ? Mdhnv6 : Eghnv6);
assign Mdhnv6 = (~(Enhnv6 & Lnhnv6));
assign Enhnv6 = (Snhnv6 & Znhnv6);
assign B0fdt6 = (~(Bihnv6 & Eghnv6));
assign Bihnv6 = (Djhnv6 & Zghnv6);
assign Zghnv6 = (Gohnv6 & Rjhnv6);
assign Gohnv6 = (Yjhnv6 & Wihnv6);
assign Yjhnv6 = (~(Nohnv6 & Uohnv6));
assign Nohnv6 = (Uhhnv6 & Snhnv6);
assign Djhnv6 = (~(Bphnv6 | Lghnv6));
assign Lghnv6 = (Uhhnv6 & Iphnv6);
assign Iphnv6 = (!Nhhnv6);
assign Nhhnv6 = (~(Pphnv6 & Snhnv6));
assign Pphnv6 = (Wphnv6 & Znhnv6);
assign Q1fdt6 = (~(Dqhnv6 & Iihnv6));
assign Iihnv6 = (~(Bphnv6 | Ghhnv6));
assign Ghhnv6 = (Kqhnv6 & Uhhnv6);
assign Kqhnv6 = (!Rqhnv6);
assign Bphnv6 = (~(Rqhnv6 | Uhhnv6));
assign Rqhnv6 = (~(Yqhnv6 & Wphnv6));
assign Dqhnv6 = (Jfhnv6 & Eghnv6);
assign Eghnv6 = (~(Yqhnv6 & Lnhnv6));
assign Yqhnv6 = (Znhnv6 & Hlhnv6);
assign Jfhnv6 = (Frhnv6 & Rjhnv6);
assign Rjhnv6 = (Mrhnv6 & Olhnv6);
assign Olhnv6 = (~(Alhnv6 & Uhhnv6));
assign Mrhnv6 = (~(Alhnv6 & Snhnv6));
assign Alhnv6 = (~(Znhnv6 | Lnhnv6));
assign Znhnv6 = (!Uohnv6);
assign Frhnv6 = (Vlhnv6 & Wihnv6);
assign Wihnv6 = (~(Qmhnv6 & Snhnv6));
assign Qmhnv6 = (Trhnv6 & Lnhnv6);
assign Lnhnv6 = (!Wphnv6);
assign Wphnv6 = (Ashnv6 ? Ide7z6[2] : Ohe7z6[6]);
assign Trhnv6 = (Uohnv6 & Hshnv6);
assign Hshnv6 = (!Uhhnv6);
assign Vlhnv6 = (~(Oshnv6 & Uohnv6));
assign Uohnv6 = (Ashnv6 ? Ide7z6[3] : Ohe7z6[7]);
assign Oshnv6 = (Uhhnv6 & Hlhnv6);
assign Hlhnv6 = (!Snhnv6);
assign Snhnv6 = (Ashnv6 ? Ide7z6[0] : N0gdt6);
assign Uhhnv6 = (Ashnv6 ? Ide7z6[1] : Ohe7z6[5]);
assign F3fdt6 = (~(Vshnv6 & Cthnv6));
assign U4fdt6 = (~(Jthnv6 & Qthnv6));
assign J6fdt6 = (~(Xthnv6 & Euhnv6));
assign Xthnv6 = (Vshnv6 & Luhnv6);
assign Y7fdt6 = (~(Suhnv6 & Zuhnv6));
assign N9fdt6 = (~(Gvhnv6 & Nvhnv6));
assign Gvhnv6 = (Vshnv6 & Uvhnv6);
assign Cbfdt6 = (~(Jthnv6 & Uvhnv6));
assign Rcfdt6 = (~(Bwhnv6 & Nvhnv6));
assign Bwhnv6 = (Vshnv6 & Iwhnv6);
assign Vshnv6 = (~(Pwhnv6 | Wwhnv6));
assign Gefdt6 = (~(Jthnv6 & Iwhnv6));
assign Jthnv6 = (Suhnv6 & Dxhnv6);
assign Suhnv6 = (~(Wwhnv6 | Kxhnv6));
assign Wwhnv6 = (Rxhnv6 & Yxhnv6);
assign Rxhnv6 = (!Fyhnv6);
assign Vffdt6 = (~(Myhnv6 & Qthnv6));
assign Khfdt6 = (~(Tyhnv6 & Cthnv6));
assign Cthnv6 = (Azhnv6 & Luhnv6);
assign Azhnv6 = (Qthnv6 & Hzhnv6);
assign Zifdt6 = (~(Ozhnv6 & Zuhnv6));
assign Zuhnv6 = (Vzhnv6 & Euhnv6);
assign Vzhnv6 = (C0inv6 & J0inv6);
assign Okfdt6 = (~(Q0inv6 & Tyhnv6));
assign Q0inv6 = (Euhnv6 & Luhnv6);
assign Luhnv6 = (X0inv6 & E1inv6);
assign E1inv6 = (~(L1inv6 & S1inv6));
assign X0inv6 = (Z1inv6 & G2inv6);
assign Euhnv6 = (N2inv6 & U2inv6);
assign U2inv6 = (~(S1inv6 & B3inv6));
assign N2inv6 = (I3inv6 ? Iwhnv6 : Qthnv6);
assign Dmfdt6 = (~(Myhnv6 & Uvhnv6));
assign Snfdt6 = (~(P3inv6 & Tyhnv6));
assign P3inv6 = (Nvhnv6 & Uvhnv6);
assign Uvhnv6 = (I3inv6 ? Qthnv6 : Iwhnv6);
assign Qthnv6 = (~(W3inv6 & D4inv6));
assign W3inv6 = (K4inv6 & Yxhnv6);
assign Hpfdt6 = (~(Myhnv6 & Iwhnv6));
assign Myhnv6 = (Ozhnv6 & Dxhnv6);
assign Dxhnv6 = (R4inv6 & C0inv6);
assign R4inv6 = (J0inv6 & Hzhnv6);
assign J0inv6 = (~(Y4inv6 & Yxhnv6));
assign Ozhnv6 = (~(Pwhnv6 | F5inv6));
assign Pwhnv6 = (M5inv6 & T5inv6);
assign M5inv6 = (Yxhnv6 & I3inv6);
assign Wqfdt6 = (~(A6inv6 & Tyhnv6));
assign Tyhnv6 = (~(F5inv6 | Kxhnv6));
assign Kxhnv6 = (H6inv6 & S1inv6);
assign H6inv6 = (T5inv6 & I3inv6);
assign F5inv6 = (~(Yxhnv6 | Fyhnv6));
assign Fyhnv6 = (~(O6inv6 & V6inv6));
assign O6inv6 = (K4inv6 & T5inv6);
assign T5inv6 = (!D4inv6);
assign A6inv6 = (Nvhnv6 & Iwhnv6);
assign Iwhnv6 = (~(C7inv6 & S1inv6));
assign C7inv6 = (D4inv6 & K4inv6);
assign Nvhnv6 = (J7inv6 & C0inv6);
assign C0inv6 = (Q7inv6 & Z1inv6);
assign Z1inv6 = (~(L1inv6 & I3inv6));
assign Q7inv6 = (~(L1inv6 & Yxhnv6));
assign L1inv6 = (~(K4inv6 | D4inv6));
assign J7inv6 = (G2inv6 & Hzhnv6);
assign Hzhnv6 = (~(B3inv6 & Yxhnv6));
assign B3inv6 = (X7inv6 & D4inv6);
assign D4inv6 = (~(E8inv6 | L8inv6));
assign E8inv6 = (Z8inv6 ? Ohe7z6[6] : S8inv6);
assign S8inv6 = (G9inv6 & N9inv6);
assign N9inv6 = (~(U9inv6 & Bainv6));
assign G9inv6 = (~(Iainv6 & Painv6));
assign X7inv6 = (V6inv6 & Wainv6);
assign G2inv6 = (~(Y4inv6 & S1inv6));
assign S1inv6 = (!Yxhnv6);
assign Yxhnv6 = (~(Dbinv6 & Kbinv6));
assign Kbinv6 = (~(Rbinv6 & Ybinv6));
assign Ybinv6 = (~(U9inv6 & Fcinv6));
assign Rbinv6 = (Mcinv6 & Tcinv6);
assign Mcinv6 = (~(Iainv6 & Bainv6));
assign Dbinv6 = (~(Adinv6 & Z8inv6));
assign Adinv6 = (Hdinv6 ? N0gdt6 : Ohe7z6[4]);
assign Y4inv6 = (Wainv6 & I3inv6);
assign I3inv6 = (!V6inv6);
assign V6inv6 = (~(Odinv6 | L8inv6));
assign Odinv6 = (Z8inv6 ? Ohe7z6[5] : Vdinv6);
assign Vdinv6 = (Ceinv6 & Jeinv6);
assign Jeinv6 = (~(Iainv6 & Qeinv6));
assign Ceinv6 = (~(U9inv6 & Xeinv6));
assign Wainv6 = (!K4inv6);
assign K4inv6 = (~(Efinv6 | L8inv6));
assign L8inv6 = (~(Lfinv6 | Z8inv6));
assign Efinv6 = (Z8inv6 ? Ohe7z6[7] : Sfinv6);
assign Z8inv6 = (!Tcinv6);
assign Sfinv6 = (~(Zfinv6 & Gginv6));
assign Zfinv6 = (~(Nginv6 & Zec7z6[9]));
assign Wagdt6 = (~(Uginv6 & Bhinv6));
assign Bhinv6 = (~(O4gdt6 & Ihinv6));
assign Lcgdt6 = (~(Phinv6 & Whinv6));
assign Whinv6 = (~(D6gdt6 & Ihinv6));
assign Zei7z6[3] = (Diinv6 & Zhbdt6);
assign Diinv6 = (Kiinv6 & Riinv6);
assign Zei7z6[2] = (Yiinv6 | Fjinv6);
assign Fjinv6 = (Pkbet6 & Mjinv6);
assign Mjinv6 = (~(Riinv6 & Tjinv6));
assign Tjinv6 = (Akinv6 | K397z6);
assign Akinv6 = (!Kgbdt6);
assign Yiinv6 = (Riinv6 ? Okinv6 : Hkinv6);
assign Okinv6 = (~(Zhbdt6 & Kiinv6));
assign Zei7z6[1] = (Riinv6 ? Clinv6 : Vkinv6);
assign Riinv6 = (~(Jlinv6 & Qlinv6));
assign Jlinv6 = (Xlinv6 & Eminv6);
assign Clinv6 = (Zhbdt6 & Lminv6);
assign Lminv6 = (~(Sminv6 & Kiinv6));
assign Kiinv6 = (Pkbet6 | Kgbdt6);
assign Sminv6 = (Pkbet6 ? Zminv6 : K397z6);
assign Zminv6 = (~(K397z6 & Kgbdt6));
assign Vkinv6 = (~(Hkinv6 | Pkbet6));
assign Hkinv6 = (K7e7z6[1] & Gninv6);
assign Nj2et6 = (Yfadt6 & Nninv6);
assign Nninv6 = (~(Uninv6 & Boinv6));
assign Boinv6 = (~(Ioinv6 | Poinv6));
assign Ioinv6 = (~(Woinv6 & Dpinv6));
assign Uninv6 = (Kpinv6 & Rpinv6);
assign Rpinv6 = (Ypinv6 | Fqinv6);
assign Wqydt6 = (~(Mqinv6 & Lxydt6));
assign Mqinv6 = (~(Tqinv6 & Ot97z6));
assign Btydt6 = (~(Arinv6 & Lxydt6));
assign Arinv6 = (~(Tqinv6 & Gt97z6));
assign Gvydt6 = (~(Tqinv6 & Hrinv6));
assign Qzydt6 = (Orinv6 & Po2et6);
assign Po2et6 = (~(Vrinv6 & Csinv6));
assign Orinv6 = (~(Jsinv6 & Qsinv6));
assign Jsinv6 = (M43et6 & K73et6);
assign V1zdt6 = (Xsinv6 & Aga7z6);
assign A4zdt6 = (Etinv6 & Aga7z6);
assign F6zdt6 = (~(Vrinv6 & Ltinv6));
assign Ltinv6 = (~(O5a7z6 & Yga7z6));
assign K8zdt6 = (Y4a7z6 & Lxydt6);
assign Pazdt6 = (~(Lxydt6 & Stinv6));
assign Uczdt6 = (~(Qga7z6 & Ztinv6));
assign Ztinv6 = (~(Qs97z6 & Lxydt6));
assign Zezdt6 = (~(Qga7z6 & Guinv6));
assign Guinv6 = (~(Ot97z6 & Lxydt6));
assign Ehzdt6 = (Gt97z6 & Lxydt6);
assign Jjzdt6 = (~(Qg2nv6 & Nuinv6));
assign Nuinv6 = (~(Ys97z6 & Lxydt6));
assign Ypzdt6 = (~(Uuinv6 & Bvinv6));
assign Dszdt6 = (Uuinv6 & Is97z6);
assign Iuzdt6 = (Uuinv6 & Qs97z6);
assign Nwzdt6 = (~(Ivinv6 & Bfo7v6));
assign Ivinv6 = (~(Uuinv6 & Ot97z6));
assign Syzdt6 = (~(Pvinv6 & Wvinv6));
assign Wvinv6 = (~(Uuinv6 & Gt97z6));
assign Pvinv6 = (~(Dwinv6 & Bfo7v6));
assign X00et6 = (~(Uuinv6 & Hrinv6));
assign C30et6 = (~(Kwinv6 & Rwinv6));
assign Rwinv6 = (~(Hbo7v6 & O5a7z6));
assign H50et6 = (Cubdt6 | Gr2et6);
assign M70et6 = (O5a7z6 & Y4a7z6);
assign R90et6 = (O5a7z6 & Is97z6);
assign Wb0et6 = (O5a7z6 & Qs97z6);
assign Li0et6 = (O5a7z6 & Ys97z6);
assign Qk0et6 = (Y4a7z6 & Aga7z6);
assign Vm0et6 = (Is97z6 & Aga7z6);
assign Ap0et6 = (~(Ywinv6 & Aga7z6));
assign Fr0et6 = (~(Dpinv6 & Aga7z6));
assign Kt0et6 = (~(Fxinv6 & Aga7z6));
assign Pv0et6 = (~(Hrinv6 & Aga7z6));
assign Ux0et6 = (Ys97z6 & Aga7z6);
assign Zz0et6 = (~(Csinv6 & Mxinv6));
assign Mxinv6 = (~(Txinv6 & O5a7z6));
assign E21et6 = (Gt97z6 & Aga7z6);
assign J41et6 = (Tnzdt6 & Y4a7z6);
assign O61et6 = (Tnzdt6 & Is97z6);
assign T81et6 = (~(Tnzdt6 & Ywinv6));
assign Ya1et6 = (Tnzdt6 & Ot97z6);
assign Dd1et6 = (~(Tnzdt6 & Fxinv6));
assign If1et6 = (~(Tnzdt6 & Hrinv6));
assign Nh1et6 = (Ot97z6 & Aga7z6);
assign Sj1et6 = (Qs97z6 & Aga7z6);
assign Xl1et6 = (Be0et6 | Ayinv6);
assign Ayinv6 = (Hyinv6 & Ypinv6);
assign Hyinv6 = (!Oyinv6);
assign Be0et6 = (O5a7z6 & Ot97z6);
assign Co1et6 = (Gg0et6 | Vyinv6);
assign Vyinv6 = (Oyinv6 & Ypinv6);
assign Gg0et6 = (O5a7z6 & Gt97z6);
assign Hq1et6 = (~(O5a7z6 & Hrinv6));
assign Ms1et6 = (Czinv6 & Y4a7z6);
assign Ru1et6 = (Czinv6 & Is97z6);
assign Ww1et6 = (Czinv6 & Qs97z6);
assign Bz1et6 = (Czinv6 ? Ot97z6 : Jzinv6);
assign Jzinv6 = (~(Oyinv6 & Qzinv6));
assign G12et6 = (Czinv6 ? Gt97z6 : Xzinv6);
assign Xzinv6 = (Oyinv6 & Qzinv6);
assign Oyinv6 = (E0jnv6 & L0jnv6);
assign E0jnv6 = (B8cdt6 & S0jnv6);
assign L32et6 = (Czinv6 ? Ys97z6 : Qzinv6);
assign Czinv6 = (~(Z0jnv6 & Lxydt6));
assign Z0jnv6 = (G1jnv6 | N1jnv6);
assign G1jnv6 = (~(U1jnv6 & B2jnv6));
assign Qzinv6 = (~(L0jnv6 & I2jnv6));
assign L0jnv6 = (P2jnv6 & B2jnv6);
assign Z72et6 = (~(Csinv6 & W2jnv6));
assign Csinv6 = (!D3jnv6);
assign Ea2et6 = (~(Kwinv6 & W2jnv6));
assign W2jnv6 = (~(Txinv6 & Gr2et6));
assign Mkxdt6 = (K3jnv6 & R3jnv6);
assign R3jnv6 = (~(Qsinv6 & Qg2nv6));
assign Smxdt6 = (~(Tnzdt6 & Bvinv6));
assign Yoxdt6 = (~(Tnzdt6 & Stinv6));
assign Stinv6 = (!Is97z6);
assign Erxdt6 = (Tnzdt6 & Qs97z6);
assign Ktxdt6 = (~(Tnzdt6 & Dpinv6));
assign Qvxdt6 = (Tnzdt6 & Gt97z6);
assign Wxxdt6 = (Tnzdt6 & Ys97z6);
assign I2ydt6 = (~(Y3jnv6 & Xsinv6));
assign O4ydt6 = (~(Bvinv6 & Qg2nv6));
assign U6ydt6 = (Is97z6 & Qg2nv6);
assign A9ydt6 = (Qs97z6 & Qg2nv6);
assign Gbydt6 = (~(Dpinv6 & Qg2nv6));
assign Dpinv6 = (!Ot97z6);
assign Mdydt6 = (~(Fxinv6 & Qg2nv6));
assign Fxinv6 = (!Gt97z6);
assign Sfydt6 = (~(Hrinv6 & Qg2nv6));
assign Hrinv6 = (!Ys97z6);
assign Yhydt6 = (~(Qg2nv6 & Y3jnv6));
assign Ekydt6 = (~(Tqinv6 & Bvinv6));
assign Bvinv6 = (!Y4a7z6);
assign Kmydt6 = (Tqinv6 & Is97z6);
assign Qoydt6 = (Tqinv6 & Qs97z6);
assign Fci7z6[1] = (~(F4jnv6 | Fci7z6[0]));
assign F4jnv6 = (M4jnv6 & T4jnv6);
assign Fci7z6[0] = (A5jnv6 & H5jnv6);
assign A5jnv6 = (O5jnv6 & V5jnv6);
assign O5jnv6 = (~(C6jnv6 & J6jnv6));
assign Zkh7z6[9] = (~(Q6jnv6 & X6jnv6));
assign X6jnv6 = (~(E7jnv6 & L7jnv6));
assign Q6jnv6 = (S7jnv6 & Z7jnv6);
assign Z7jnv6 = (~(vis_pc_o[9] & G8jnv6));
assign S7jnv6 = (N8jnv6 | U8jnv6);
assign Zkh7z6[8] = (~(B9jnv6 & I9jnv6));
assign I9jnv6 = (~(E7jnv6 & P9jnv6));
assign B9jnv6 = (W9jnv6 & Dajnv6);
assign Dajnv6 = (~(vis_pc_o[8] & G8jnv6));
assign W9jnv6 = (N8jnv6 | Kajnv6);
assign Zkh7z6[7] = (~(Rajnv6 & Yajnv6));
assign Yajnv6 = (~(E7jnv6 & Fbjnv6));
assign Rajnv6 = (Mbjnv6 & Tbjnv6);
assign Tbjnv6 = (~(vis_pc_o[7] & G8jnv6));
assign Mbjnv6 = (N8jnv6 | Acjnv6);
assign Zkh7z6[6] = (~(Hcjnv6 & Ocjnv6));
assign Ocjnv6 = (~(E7jnv6 & Vcjnv6));
assign Hcjnv6 = (Cdjnv6 & Jdjnv6);
assign Jdjnv6 = (~(vis_pc_o[6] & G8jnv6));
assign Cdjnv6 = (N8jnv6 | Qdjnv6);
assign Zkh7z6[5] = (~(Xdjnv6 & Eejnv6));
assign Eejnv6 = (~(E7jnv6 & Lejnv6));
assign Xdjnv6 = (Sejnv6 & Zejnv6);
assign Zejnv6 = (~(vis_pc_o[5] & G8jnv6));
assign Sejnv6 = (N8jnv6 | Gfjnv6);
assign Zkh7z6[4] = (~(Nfjnv6 & Ufjnv6));
assign Ufjnv6 = (~(E7jnv6 & Bgjnv6));
assign Nfjnv6 = (Igjnv6 & Pgjnv6);
assign Pgjnv6 = (~(vis_pc_o[4] & G8jnv6));
assign Igjnv6 = (N8jnv6 | Wgjnv6);
assign Zkh7z6[3] = (~(Dhjnv6 & Khjnv6));
assign Khjnv6 = (~(E7jnv6 & Rhjnv6));
assign Dhjnv6 = (Yhjnv6 & Fijnv6);
assign Fijnv6 = (~(vis_pc_o[3] & G8jnv6));
assign Yhjnv6 = (N8jnv6 | Mijnv6);
assign Zkh7z6[31] = (~(Tijnv6 & Ajjnv6));
assign Ajjnv6 = (~(E7jnv6 & Hjjnv6));
assign Tijnv6 = (Ojjnv6 & Vjjnv6);
assign Vjjnv6 = (~(vis_pc_o[31] & G8jnv6));
assign Ojjnv6 = (N8jnv6 | Ckjnv6);
assign Zkh7z6[30] = (~(Jkjnv6 & Qkjnv6));
assign Qkjnv6 = (~(E7jnv6 & Xkjnv6));
assign Jkjnv6 = (Eljnv6 & Lljnv6);
assign Lljnv6 = (~(vis_pc_o[30] & G8jnv6));
assign Eljnv6 = (N8jnv6 | Sljnv6);
assign Zkh7z6[2] = (~(Zljnv6 & Gmjnv6));
assign Gmjnv6 = (~(E7jnv6 & Nmjnv6));
assign Zljnv6 = (Umjnv6 & Bnjnv6);
assign Bnjnv6 = (~(vis_pc_o[2] & G8jnv6));
assign Umjnv6 = (N8jnv6 | Injnv6);
assign Zkh7z6[29] = (~(Pnjnv6 & Wnjnv6));
assign Wnjnv6 = (~(E7jnv6 & Dojnv6));
assign Pnjnv6 = (Kojnv6 & Rojnv6);
assign Rojnv6 = (~(vis_pc_o[29] & G8jnv6));
assign Kojnv6 = (N8jnv6 | Yojnv6);
assign Zkh7z6[28] = (~(Fpjnv6 & Mpjnv6));
assign Mpjnv6 = (~(E7jnv6 & Tpjnv6));
assign Fpjnv6 = (Aqjnv6 & Hqjnv6);
assign Hqjnv6 = (~(vis_pc_o[28] & G8jnv6));
assign Aqjnv6 = (N8jnv6 | Oqjnv6);
assign Zkh7z6[27] = (~(Vqjnv6 & Crjnv6));
assign Crjnv6 = (~(E7jnv6 & Jrjnv6));
assign Vqjnv6 = (Qrjnv6 & Xrjnv6);
assign Xrjnv6 = (~(vis_pc_o[27] & G8jnv6));
assign Qrjnv6 = (N8jnv6 | Esjnv6);
assign Zkh7z6[26] = (~(Lsjnv6 & Ssjnv6));
assign Ssjnv6 = (~(E7jnv6 & Zsjnv6));
assign Lsjnv6 = (Gtjnv6 & Ntjnv6);
assign Ntjnv6 = (~(vis_pc_o[26] & G8jnv6));
assign Gtjnv6 = (N8jnv6 | Utjnv6);
assign Zkh7z6[25] = (~(Bujnv6 & Iujnv6));
assign Iujnv6 = (~(E7jnv6 & Pujnv6));
assign Bujnv6 = (Wujnv6 & Dvjnv6);
assign Dvjnv6 = (~(vis_pc_o[25] & G8jnv6));
assign Wujnv6 = (N8jnv6 | Kvjnv6);
assign Zkh7z6[24] = (~(Rvjnv6 & Yvjnv6));
assign Yvjnv6 = (~(E7jnv6 & Fwjnv6));
assign Rvjnv6 = (Mwjnv6 & Twjnv6);
assign Twjnv6 = (~(vis_pc_o[24] & G8jnv6));
assign Mwjnv6 = (N8jnv6 | Axjnv6);
assign Zkh7z6[23] = (~(Hxjnv6 & Oxjnv6));
assign Oxjnv6 = (~(E7jnv6 & Vxjnv6));
assign Hxjnv6 = (Cyjnv6 & Jyjnv6);
assign Jyjnv6 = (~(vis_pc_o[23] & G8jnv6));
assign Cyjnv6 = (N8jnv6 | Qyjnv6);
assign Zkh7z6[22] = (~(Xyjnv6 & Ezjnv6));
assign Ezjnv6 = (~(E7jnv6 & Lzjnv6));
assign Xyjnv6 = (Szjnv6 & Zzjnv6);
assign Zzjnv6 = (~(vis_pc_o[22] & G8jnv6));
assign Szjnv6 = (N8jnv6 | G0knv6);
assign Zkh7z6[21] = (~(N0knv6 & U0knv6));
assign U0knv6 = (~(E7jnv6 & B1knv6));
assign N0knv6 = (I1knv6 & P1knv6);
assign P1knv6 = (~(vis_pc_o[21] & G8jnv6));
assign I1knv6 = (N8jnv6 | W1knv6);
assign Zkh7z6[20] = (~(D2knv6 & K2knv6));
assign K2knv6 = (~(E7jnv6 & R2knv6));
assign D2knv6 = (Y2knv6 & F3knv6);
assign F3knv6 = (~(vis_pc_o[20] & G8jnv6));
assign Y2knv6 = (N8jnv6 | M3knv6);
assign Zkh7z6[1] = (~(T3knv6 & A4knv6));
assign A4knv6 = (N8jnv6 | H4knv6);
assign T3knv6 = (O4knv6 & V4knv6);
assign V4knv6 = (~(C5knv6 & E7jnv6));
assign C5knv6 = (~(J5knv6 | Q5knv6));
assign O4knv6 = (~(vis_pc_o[1] & G8jnv6));
assign Zkh7z6[19] = (~(X5knv6 & E6knv6));
assign E6knv6 = (~(E7jnv6 & L6knv6));
assign X5knv6 = (S6knv6 & Z6knv6);
assign Z6knv6 = (~(vis_pc_o[19] & G8jnv6));
assign S6knv6 = (N8jnv6 | G7knv6);
assign Zkh7z6[18] = (~(N7knv6 & U7knv6));
assign U7knv6 = (~(E7jnv6 & B8knv6));
assign N7knv6 = (I8knv6 & P8knv6);
assign P8knv6 = (~(vis_pc_o[18] & G8jnv6));
assign I8knv6 = (N8jnv6 | W8knv6);
assign Zkh7z6[17] = (~(D9knv6 & K9knv6));
assign K9knv6 = (~(E7jnv6 & R9knv6));
assign D9knv6 = (Y9knv6 & Faknv6);
assign Faknv6 = (~(vis_pc_o[17] & G8jnv6));
assign Y9knv6 = (N8jnv6 | Maknv6);
assign Zkh7z6[16] = (~(Taknv6 & Abknv6));
assign Abknv6 = (~(E7jnv6 & Hbknv6));
assign Taknv6 = (Obknv6 & Vbknv6);
assign Vbknv6 = (~(vis_pc_o[16] & G8jnv6));
assign Obknv6 = (N8jnv6 | Ccknv6);
assign Zkh7z6[15] = (~(Jcknv6 & Qcknv6));
assign Qcknv6 = (~(E7jnv6 & Xcknv6));
assign Jcknv6 = (Edknv6 & Ldknv6);
assign Ldknv6 = (~(vis_pc_o[15] & G8jnv6));
assign Edknv6 = (N8jnv6 | Sdknv6);
assign Zkh7z6[14] = (~(Zdknv6 & Geknv6));
assign Geknv6 = (~(E7jnv6 & Neknv6));
assign Zdknv6 = (Ueknv6 & Bfknv6);
assign Bfknv6 = (~(vis_pc_o[14] & G8jnv6));
assign Ueknv6 = (N8jnv6 | Ifknv6);
assign Zkh7z6[13] = (~(Pfknv6 & Wfknv6));
assign Wfknv6 = (~(E7jnv6 & Dgknv6));
assign Pfknv6 = (Kgknv6 & Rgknv6);
assign Rgknv6 = (~(vis_pc_o[13] & G8jnv6));
assign Kgknv6 = (N8jnv6 | Ygknv6);
assign Zkh7z6[12] = (~(Fhknv6 & Mhknv6));
assign Mhknv6 = (~(E7jnv6 & Thknv6));
assign Fhknv6 = (Aiknv6 & Hiknv6);
assign Hiknv6 = (~(vis_pc_o[12] & G8jnv6));
assign Aiknv6 = (N8jnv6 | Oiknv6);
assign Zkh7z6[11] = (~(Viknv6 & Cjknv6));
assign Cjknv6 = (~(E7jnv6 & Jjknv6));
assign Viknv6 = (Qjknv6 & Xjknv6);
assign Xjknv6 = (~(vis_pc_o[11] & G8jnv6));
assign Qjknv6 = (~(Ekknv6 & Lkknv6));
assign Zkh7z6[10] = (~(Skknv6 & Zkknv6));
assign Zkknv6 = (~(E7jnv6 & Glknv6));
assign Skknv6 = (Nlknv6 & Ulknv6);
assign Ulknv6 = (~(vis_pc_o[10] & G8jnv6));
assign G8jnv6 = (~(Bmknv6 | E7jnv6));
assign Nlknv6 = (~(Ekknv6 & Imknv6));
assign Ekknv6 = (!N8jnv6);
assign Zkh7z6[0] = (!Pmknv6);
assign Vvh7z6[9] = (Wmknv6 ? Fth7z6[9] : Kxb7z6[9]);
assign Vvh7z6[8] = (Wmknv6 ? Fth7z6[8] : Kxb7z6[8]);
assign Vvh7z6[7] = (Wmknv6 ? Fth7z6[7] : Kxb7z6[7]);
assign Vvh7z6[6] = (Wmknv6 ? Fth7z6[6] : Kxb7z6[6]);
assign Vvh7z6[5] = (Wmknv6 ? Fth7z6[5] : Kxb7z6[5]);
assign Vvh7z6[4] = (Wmknv6 ? Fth7z6[4] : Kxb7z6[4]);
assign Vvh7z6[3] = (Wmknv6 ? Fth7z6[3] : Kxb7z6[3]);
assign Vvh7z6[31] = (Wmknv6 ? Fth7z6[31] : Kxb7z6[31]);
assign Vvh7z6[30] = (Wmknv6 ? Fth7z6[30] : Kxb7z6[30]);
assign Vvh7z6[2] = (Wmknv6 ? Fth7z6[2] : Kxb7z6[2]);
assign Vvh7z6[29] = (Wmknv6 ? Fth7z6[29] : Kxb7z6[29]);
assign Vvh7z6[28] = (Wmknv6 ? Fth7z6[28] : Kxb7z6[28]);
assign Vvh7z6[27] = (Wmknv6 ? Fth7z6[27] : Kxb7z6[27]);
assign Vvh7z6[26] = (Wmknv6 ? Fth7z6[26] : Kxb7z6[26]);
assign Vvh7z6[25] = (Wmknv6 ? Fth7z6[25] : Kxb7z6[25]);
assign Vvh7z6[24] = (Wmknv6 ? Fth7z6[24] : Kxb7z6[24]);
assign Vvh7z6[23] = (Wmknv6 ? Fth7z6[23] : Kxb7z6[23]);
assign Vvh7z6[22] = (Wmknv6 ? Fth7z6[22] : Kxb7z6[22]);
assign Vvh7z6[21] = (Wmknv6 ? Fth7z6[21] : Kxb7z6[21]);
assign Vvh7z6[20] = (Wmknv6 ? Fth7z6[20] : Kxb7z6[20]);
assign Vvh7z6[1] = (Wmknv6 ? Fth7z6[1] : Kxb7z6[1]);
assign Vvh7z6[19] = (Wmknv6 ? Fth7z6[19] : Kxb7z6[19]);
assign Vvh7z6[18] = (Wmknv6 ? Fth7z6[18] : Kxb7z6[18]);
assign Vvh7z6[17] = (Wmknv6 ? Fth7z6[17] : Kxb7z6[17]);
assign Vvh7z6[16] = (Wmknv6 ? Fth7z6[16] : Kxb7z6[16]);
assign Vvh7z6[15] = (Wmknv6 ? Fth7z6[15] : Kxb7z6[15]);
assign Vvh7z6[14] = (Wmknv6 ? Fth7z6[14] : Kxb7z6[14]);
assign Vvh7z6[13] = (Wmknv6 ? Fth7z6[13] : Kxb7z6[13]);
assign Vvh7z6[12] = (Wmknv6 ? Fth7z6[12] : Kxb7z6[12]);
assign Vvh7z6[11] = (Wmknv6 ? Fth7z6[11] : Kxb7z6[11]);
assign Vvh7z6[10] = (Wmknv6 ? Fth7z6[10] : Kxb7z6[10]);
assign Vvh7z6[0] = (Wmknv6 ? Fth7z6[0] : Kxb7z6[0]);
assign Ed5et6 = (~(Dnknv6 ^ Ueo7v6));
assign Dnknv6 = (Knknv6 & Rnknv6);
assign Rnknv6 = (~(Ynknv6 & E3c7z6[0]));
assign Knknv6 = (~(Foknv6 & V1c7z6[0]));
assign Nf5et6 = (~(Moknv6 ^ Ueo7v6));
assign Moknv6 = (Toknv6 & Apknv6);
assign Apknv6 = (~(Foknv6 & V1c7z6[1]));
assign Toknv6 = (Hpknv6 & Opknv6);
assign Opknv6 = (~(Ynknv6 & E3c7z6[1]));
assign Hpknv6 = (~(Vpknv6 & Fth7z6[0]));
assign Wh5et6 = (~(Cqknv6 ^ Ueo7v6));
assign Cqknv6 = (Jqknv6 & Qqknv6);
assign Qqknv6 = (Xqknv6 & Erknv6);
assign Erknv6 = (~(Ynknv6 & E3c7z6[2]));
assign Xqknv6 = (Lrknv6 & Srknv6);
assign Lrknv6 = (~(Foknv6 & V1c7z6[2]));
assign Jqknv6 = (Zrknv6 & Gsknv6);
assign Gsknv6 = (~(Vpknv6 & Fth7z6[1]));
assign Fk5et6 = (~(Nsknv6 ^ Ueo7v6));
assign Nsknv6 = (Usknv6 & Btknv6);
assign Btknv6 = (Itknv6 & Ptknv6);
assign Ptknv6 = (~(Ynknv6 & E3c7z6[3]));
assign Usknv6 = (Wtknv6 & Duknv6);
assign Duknv6 = (~(Foknv6 & V1c7z6[3]));
assign Wtknv6 = (~(Vpknv6 & Fth7z6[2]));
assign Om5et6 = (~(Kuknv6 ^ Ueo7v6));
assign Kuknv6 = (Ruknv6 & Yuknv6);
assign Yuknv6 = (Fvknv6 & Mvknv6);
assign Mvknv6 = (~(Ynknv6 & E3c7z6[4]));
assign Ruknv6 = (Tvknv6 & Awknv6);
assign Awknv6 = (~(Foknv6 & V1c7z6[4]));
assign Tvknv6 = (~(Vpknv6 & Fth7z6[3]));
assign Xo5et6 = (~(Hwknv6 ^ Ueo7v6));
assign Hwknv6 = (Owknv6 & Vwknv6);
assign Vwknv6 = (Cxknv6 & Jxknv6);
assign Jxknv6 = (Qxknv6 & Xxknv6);
assign Cxknv6 = (~(Eyknv6 | Lyknv6));
assign Owknv6 = (Syknv6 & Zyknv6);
assign Zyknv6 = (Gzknv6 & Nzknv6);
assign Gzknv6 = (~(Vpknv6 & Fth7z6[4]));
assign Syknv6 = (Uzknv6 & B0lnv6);
assign B0lnv6 = (~(Foknv6 & V1c7z6[5]));
assign Uzknv6 = (~(Ynknv6 & Fhc7z6[5]));
assign Gr5et6 = (~(I0lnv6 ^ Ueo7v6));
assign I0lnv6 = (P0lnv6 & W0lnv6);
assign W0lnv6 = (D1lnv6 & K1lnv6);
assign K1lnv6 = (~(Foknv6 & V1c7z6[6]));
assign P0lnv6 = (R1lnv6 & Y1lnv6);
assign Y1lnv6 = (~(Ynknv6 & Fhc7z6[6]));
assign R1lnv6 = (~(Vpknv6 & Fth7z6[5]));
assign Pt5et6 = (~(F2lnv6 ^ Ueo7v6));
assign F2lnv6 = (M2lnv6 & T2lnv6);
assign T2lnv6 = (A3lnv6 & H3lnv6);
assign H3lnv6 = (~(Foknv6 & V1c7z6[7]));
assign M2lnv6 = (O3lnv6 & V3lnv6);
assign V3lnv6 = (~(Ynknv6 & Fhc7z6[7]));
assign O3lnv6 = (~(Vpknv6 & Fth7z6[6]));
assign Yv5et6 = (~(C4lnv6 ^ Ueo7v6));
assign C4lnv6 = (J4lnv6 & Q4lnv6);
assign Q4lnv6 = (~(Ynknv6 & Fhc7z6[8]));
assign J4lnv6 = (X4lnv6 & E5lnv6);
assign E5lnv6 = (~(Foknv6 & V1c7z6[8]));
assign X4lnv6 = (~(Vpknv6 & Fth7z6[7]));
assign Hy5et6 = (~(L5lnv6 ^ Ueo7v6));
assign L5lnv6 = (S5lnv6 & Z5lnv6);
assign Z5lnv6 = (~(Ynknv6 & Fhc7z6[9]));
assign S5lnv6 = (G6lnv6 & N6lnv6);
assign N6lnv6 = (~(Foknv6 & V1c7z6[9]));
assign G6lnv6 = (~(Vpknv6 & Fth7z6[8]));
assign Q06et6 = (~(U6lnv6 ^ Ueo7v6));
assign U6lnv6 = (B7lnv6 & I7lnv6);
assign I7lnv6 = (~(Ynknv6 & Fhc7z6[10]));
assign B7lnv6 = (P7lnv6 & W7lnv6);
assign W7lnv6 = (~(Foknv6 & V1c7z6[10]));
assign P7lnv6 = (~(Vpknv6 & Fth7z6[9]));
assign Z26et6 = (~(D8lnv6 ^ Ueo7v6));
assign D8lnv6 = (K8lnv6 & R8lnv6);
assign R8lnv6 = (~(Ynknv6 & Fhc7z6[11]));
assign K8lnv6 = (Y8lnv6 & F9lnv6);
assign F9lnv6 = (~(Foknv6 & V1c7z6[11]));
assign Y8lnv6 = (~(Vpknv6 & Fth7z6[10]));
assign I56et6 = (~(M9lnv6 ^ Ueo7v6));
assign M9lnv6 = (T9lnv6 & Aalnv6);
assign Aalnv6 = (~(Ynknv6 & Fhc7z6[12]));
assign T9lnv6 = (Halnv6 & Oalnv6);
assign Oalnv6 = (~(Foknv6 & V1c7z6[12]));
assign Halnv6 = (~(Vpknv6 & Fth7z6[11]));
assign R76et6 = (~(Valnv6 ^ Ueo7v6));
assign Valnv6 = (Cblnv6 & Jblnv6);
assign Jblnv6 = (~(Ynknv6 & Fhc7z6[13]));
assign Cblnv6 = (Qblnv6 & Xblnv6);
assign Xblnv6 = (~(Foknv6 & V1c7z6[13]));
assign Qblnv6 = (~(Vpknv6 & Fth7z6[12]));
assign Aa6et6 = (~(Eclnv6 ^ Ueo7v6));
assign Eclnv6 = (Lclnv6 & Sclnv6);
assign Sclnv6 = (~(Ynknv6 & Fhc7z6[14]));
assign Lclnv6 = (Zclnv6 & Gdlnv6);
assign Gdlnv6 = (~(Foknv6 & V1c7z6[14]));
assign Zclnv6 = (~(Vpknv6 & Fth7z6[13]));
assign Jc6et6 = (~(Ndlnv6 ^ Ueo7v6));
assign Ndlnv6 = (Udlnv6 & Belnv6);
assign Belnv6 = (~(Ynknv6 & Fhc7z6[15]));
assign Udlnv6 = (Ielnv6 & Pelnv6);
assign Pelnv6 = (~(Foknv6 & V1c7z6[15]));
assign Ielnv6 = (~(Vpknv6 & Fth7z6[14]));
assign Se6et6 = (~(Welnv6 ^ Ueo7v6));
assign Welnv6 = (Dflnv6 & Kflnv6);
assign Kflnv6 = (~(Ynknv6 & Fhc7z6[16]));
assign Dflnv6 = (Rflnv6 & Yflnv6);
assign Yflnv6 = (~(Foknv6 & V1c7z6[16]));
assign Rflnv6 = (~(Vpknv6 & Fth7z6[15]));
assign Bh6et6 = (~(Fglnv6 ^ Ueo7v6));
assign Fglnv6 = (Mglnv6 & Tglnv6);
assign Tglnv6 = (~(Foknv6 & V1c7z6[17]));
assign Mglnv6 = (~(Ynknv6 & Fhc7z6[17]));
assign Kj6et6 = (~(Ahlnv6 ^ Ueo7v6));
assign Ahlnv6 = (Hhlnv6 & Ohlnv6);
assign Ohlnv6 = (~(Foknv6 & V1c7z6[18]));
assign Hhlnv6 = (~(Ynknv6 & Fhc7z6[18]));
assign Tl6et6 = (~(Vhlnv6 ^ Ueo7v6));
assign Vhlnv6 = (Cilnv6 & Jilnv6);
assign Jilnv6 = (~(Foknv6 & V1c7z6[19]));
assign Cilnv6 = (~(Ynknv6 & Fhc7z6[19]));
assign Co6et6 = (~(Qilnv6 ^ Ueo7v6));
assign Qilnv6 = (Xilnv6 & Ejlnv6);
assign Ejlnv6 = (~(Foknv6 & V1c7z6[20]));
assign Xilnv6 = (~(Ynknv6 & Fhc7z6[20]));
assign Lq6et6 = (~(Ljlnv6 ^ Ueo7v6));
assign Ljlnv6 = (Sjlnv6 & Zjlnv6);
assign Zjlnv6 = (~(Foknv6 & V1c7z6[21]));
assign Sjlnv6 = (~(Ynknv6 & Fhc7z6[21]));
assign Us6et6 = (~(Gklnv6 ^ Ueo7v6));
assign Gklnv6 = (Nklnv6 & Uklnv6);
assign Uklnv6 = (~(Foknv6 & V1c7z6[22]));
assign Nklnv6 = (~(Ynknv6 & Fhc7z6[22]));
assign Dv6et6 = (~(Bllnv6 ^ Ueo7v6));
assign Bllnv6 = (Illnv6 & Pllnv6);
assign Pllnv6 = (~(Foknv6 & V1c7z6[23]));
assign Illnv6 = (~(Ynknv6 & Fhc7z6[23]));
assign Mx6et6 = (~(Wllnv6 ^ Ueo7v6));
assign Wllnv6 = (Dmlnv6 & Kmlnv6);
assign Kmlnv6 = (~(Foknv6 & V1c7z6[24]));
assign Dmlnv6 = (~(Ynknv6 & Fhc7z6[24]));
assign Vz6et6 = (~(Rmlnv6 ^ Ueo7v6));
assign Rmlnv6 = (Ymlnv6 & Fnlnv6);
assign Fnlnv6 = (~(Foknv6 & V1c7z6[25]));
assign Ymlnv6 = (~(Ynknv6 & Fhc7z6[25]));
assign E27et6 = (~(Mnlnv6 ^ Ueo7v6));
assign Mnlnv6 = (Tnlnv6 & Aolnv6);
assign Aolnv6 = (~(Foknv6 & V1c7z6[26]));
assign Tnlnv6 = (~(Ynknv6 & Fhc7z6[26]));
assign N47et6 = (~(Holnv6 ^ Ueo7v6));
assign Holnv6 = (Oolnv6 & Volnv6);
assign Volnv6 = (~(Foknv6 & V1c7z6[27]));
assign Oolnv6 = (~(Ynknv6 & Fhc7z6[27]));
assign W67et6 = (~(Cplnv6 ^ Ueo7v6));
assign Cplnv6 = (Jplnv6 & Qplnv6);
assign Qplnv6 = (~(Foknv6 & V1c7z6[28]));
assign Jplnv6 = (~(Ynknv6 & Fhc7z6[28]));
assign F97et6 = (Xplnv6 ^ Eqlnv6);
assign Xplnv6 = (Lqlnv6 & Sqlnv6);
assign Sqlnv6 = (~(Foknv6 & V1c7z6[29]));
assign Lqlnv6 = (~(Ynknv6 & Fhc7z6[29]));
assign Ob7et6 = (Zqlnv6 ^ Eqlnv6);
assign Zqlnv6 = (Grlnv6 & Nrlnv6);
assign Nrlnv6 = (~(Foknv6 & V1c7z6[30]));
assign Grlnv6 = (~(Ynknv6 & Fhc7z6[30]));
assign Xd7et6 = (Urlnv6 ^ Eqlnv6);
assign Urlnv6 = (Bslnv6 & Islnv6);
assign Islnv6 = (~(Foknv6 & V1c7z6[31]));
assign Foknv6 = (T3cdt6 & Pslnv6);
assign Pslnv6 = (!Wslnv6);
assign Bslnv6 = (~(Ynknv6 & Fhc7z6[31]));
assign Ynknv6 = (~(Wslnv6 | T3cdt6));
assign Wslnv6 = (Dtlnv6 & Ktlnv6);
assign Ktlnv6 = (~(Rtlnv6 & Ytlnv6));
assign Rtlnv6 = (Fulnv6 & Dwb7z6[4]);
assign Dtlnv6 = (Mulnv6 & Tulnv6);
assign Zyaet6 = (~(Avlnv6 ^ Hvlnv6));
assign Avlnv6 = (~(Zrknv6 & Ovlnv6));
assign Ovlnv6 = (~(V1c7z6[2] & Vvlnv6));
assign Zrknv6 = (~(Q1h7z6[0] & Cwlnv6));
assign I1bet6 = (~(Jwlnv6 ^ Hvlnv6));
assign Jwlnv6 = (~(Itknv6 & Qwlnv6));
assign Qwlnv6 = (~(V1c7z6[3] & Vvlnv6));
assign Itknv6 = (~(Q1h7z6[1] & Cwlnv6));
assign R3bet6 = (~(Xwlnv6 ^ Hvlnv6));
assign Xwlnv6 = (~(Fvknv6 & Exlnv6));
assign Exlnv6 = (~(V1c7z6[4] & Vvlnv6));
assign Fvknv6 = (~(Q1h7z6[2] & Cwlnv6));
assign A6bet6 = (~(Lxlnv6 ^ Hvlnv6));
assign Lxlnv6 = (~(Nzknv6 & Sxlnv6));
assign Sxlnv6 = (~(V1c7z6[5] & Vvlnv6));
assign Nzknv6 = (~(Q1h7z6[3] & Cwlnv6));
assign J8bet6 = (~(Zxlnv6 ^ Hvlnv6));
assign Hvlnv6 = (!Cfa7z6);
assign Zxlnv6 = (~(D1lnv6 & Gylnv6));
assign Gylnv6 = (~(V1c7z6[6] & Vvlnv6));
assign D1lnv6 = (~(Q1h7z6[4] & Cwlnv6));
assign Sabet6 = (Nylnv6 ^ Cfa7z6);
assign Nylnv6 = (~(A3lnv6 & Uylnv6));
assign Uylnv6 = (~(V1c7z6[7] & Vvlnv6));
assign A3lnv6 = (~(Q1h7z6[5] & Cwlnv6));
assign Bdbet6 = (Cfa7z6 ^ Bzlnv6);
assign Bzlnv6 = (V1c7z6[8] & Vvlnv6);
assign Kfbet6 = (Cfa7z6 ^ Izlnv6);
assign Izlnv6 = (V1c7z6[9] & Vvlnv6);
assign U3d7z6[5] = (~(Pzlnv6 & Wzlnv6));
assign Wzlnv6 = (~(D0mnv6 & Bfd7z6[5]));
assign Pzlnv6 = (K0mnv6 | R0mnv6);
assign U3d7z6[4] = (~(Y0mnv6 & F1mnv6));
assign F1mnv6 = (~(M1mnv6 & T1mnv6));
assign Y0mnv6 = (A2mnv6 & H2mnv6);
assign A2mnv6 = (~(Bfd7z6[4] & D0mnv6));
assign U3d7z6[3] = (~(O2mnv6 & V2mnv6));
assign V2mnv6 = (~(D0mnv6 & Bfd7z6[3]));
assign O2mnv6 = (C3mnv6 | R0mnv6);
assign U3d7z6[2] = (~(J3mnv6 & Q3mnv6));
assign Q3mnv6 = (~(Bfd7z6[2] & D0mnv6));
assign J3mnv6 = (X3mnv6 | R0mnv6);
assign U3d7z6[1] = (~(E4mnv6 & L4mnv6));
assign L4mnv6 = (R0mnv6 | S4mnv6);
assign R0mnv6 = (!T1mnv6);
assign E4mnv6 = (Z4mnv6 & G5mnv6);
assign G5mnv6 = (~(N5mnv6 & U5mnv6));
assign N5mnv6 = (B6mnv6 & H2mnv6);
assign Z4mnv6 = (~(D0mnv6 & Bfd7z6[1]));
assign U3d7z6[0] = (~(I6mnv6 & P6mnv6));
assign P6mnv6 = (~(T1mnv6 & W6mnv6));
assign T1mnv6 = (~(D7mnv6 | Mao7v6));
assign I6mnv6 = (K7mnv6 & R7mnv6);
assign R7mnv6 = (~(Y7mnv6 & F8mnv6));
assign Y7mnv6 = (U5mnv6 & H2mnv6);
assign K7mnv6 = (~(Bfd7z6[0] & D0mnv6));
assign D0mnv6 = (M8mnv6 & H2mnv6);
assign Zgddt6 = (T8mnv6 & A9mnv6);
assign T8mnv6 = (~(H9mnv6 & O9mnv6));
assign O9mnv6 = (~(V9mnv6 & Lfinv6));
assign Lfinv6 = (~(U9inv6 & Iainv6));
assign Iainv6 = (!Nginv6);
assign H9mnv6 = (~(Camnv6 & Jamnv6));
assign Yxd7z6[1] = (Yxd7z6[0] & A4a7z6);
assign S0e7z6[5] = (Yxd7z6[0] & Zec7z6[9]);
assign S0e7z6[4] = (Yxd7z6[0] & Zec7z6[7]);
assign S0e7z6[3] = (Yxd7z6[0] & Zec7z6[6]);
assign S0e7z6[2] = (Yxd7z6[0] & Zec7z6[5]);
assign S0e7z6[1] = (Yxd7z6[0] & Zec7z6[4]);
assign S0e7z6[0] = (Yxd7z6[0] & Zec7z6[3]);
assign Pcg7z6[9] = (Qamnv6 ? Ebwdt6 : Qptdt6);
assign Pcg7z6[8] = (Qamnv6 ? Bewdt6 : Ostdt6);
assign Pcg7z6[7] = (Qamnv6 ? Ygwdt6 : Mvtdt6);
assign Pcg7z6[6] = (Qamnv6 ? Vjwdt6 : Kytdt6);
assign Pcg7z6[5] = (Qamnv6 ? Smwdt6 : I1udt6);
assign Pcg7z6[4] = (Qamnv6 ? Ppwdt6 : G4udt6);
assign Pcg7z6[3] = (Qamnv6 ? Mswdt6 : E7udt6);
assign Pcg7z6[30] = (Qamnv6 ? Uludt6 : G0sdt6);
assign Pcg7z6[2] = (Qamnv6 ? Jvwdt6 : Caudt6);
assign Pcg7z6[29] = (Qamnv6 ? Soudt6 : E3sdt6);
assign Pcg7z6[28] = (Qamnv6 ? Qrudt6 : C6sdt6);
assign Pcg7z6[27] = (Qamnv6 ? Ouudt6 : A9sdt6);
assign Pcg7z6[26] = (Qamnv6 ? Mxudt6 : Ybsdt6);
assign Pcg7z6[25] = (Qamnv6 ? K0vdt6 : Wesdt6);
assign Pcg7z6[24] = (Qamnv6 ? I3vdt6 : Uhsdt6);
assign Pcg7z6[23] = (Qamnv6 ? G6vdt6 : Sksdt6);
assign Pcg7z6[22] = (Qamnv6 ? E9vdt6 : Qnsdt6);
assign Pcg7z6[21] = (Qamnv6 ? Ccvdt6 : Oqsdt6);
assign Pcg7z6[20] = (Qamnv6 ? Afvdt6 : Mtsdt6);
assign Pcg7z6[1] = (Qamnv6 ? Gywdt6 : Adudt6);
assign Pcg7z6[19] = (Qamnv6 ? Yhvdt6 : Kwsdt6);
assign Pcg7z6[18] = (Qamnv6 ? Wkvdt6 : Izsdt6);
assign Pcg7z6[17] = (Qamnv6 ? Unvdt6 : G2tdt6);
assign Pcg7z6[16] = (Qamnv6 ? Sqvdt6 : E5tdt6);
assign Pcg7z6[15] = (Qamnv6 ? Qtvdt6 : C8tdt6);
assign Pcg7z6[14] = (Qamnv6 ? Owvdt6 : Abtdt6);
assign Pcg7z6[13] = (Qamnv6 ? Mzvdt6 : Ydtdt6);
assign Pcg7z6[12] = (Qamnv6 ? K2wdt6 : Wgtdt6);
assign Pcg7z6[11] = (Qamnv6 ? I5wdt6 : Ujtdt6);
assign Pcg7z6[10] = (Qamnv6 ? G8wdt6 : Smtdt6);
assign Pcg7z6[0] = (Qamnv6 ? D1xdt6 : Yfudt6);
assign Jjg7z6[9] = (~(Xamnv6 ^ Alf7z6[9]));
assign Jjg7z6[8] = (~(Xamnv6 ^ Alf7z6[8]));
assign Jjg7z6[7] = (~(Xamnv6 ^ Alf7z6[7]));
assign Jjg7z6[6] = (~(Xamnv6 ^ Alf7z6[6]));
assign Jjg7z6[5] = (~(Xamnv6 ^ Alf7z6[5]));
assign Jjg7z6[4] = (~(Xamnv6 ^ Alf7z6[4]));
assign Jjg7z6[3] = (~(Xamnv6 ^ Alf7z6[3]));
assign Jjg7z6[32] = (~(Xamnv6 ^ A4xdt6));
assign A4xdt6 = (Elgdt6 & Alf7z6[31]);
assign Jjg7z6[31] = (Xamnv6 ^ Ebmnv6);
assign Jjg7z6[30] = (Wvl8v6 ^ Alf7z6[30]);
assign Jjg7z6[2] = (~(Xamnv6 ^ Alf7z6[2]));
assign Jjg7z6[29] = (~(Xamnv6 ^ Alf7z6[29]));
assign Jjg7z6[28] = (~(Xamnv6 ^ Alf7z6[28]));
assign Jjg7z6[27] = (~(Xamnv6 ^ Alf7z6[27]));
assign Jjg7z6[26] = (~(Xamnv6 ^ Alf7z6[26]));
assign Jjg7z6[25] = (~(Xamnv6 ^ Alf7z6[25]));
assign Jjg7z6[24] = (~(Xamnv6 ^ Alf7z6[24]));
assign Jjg7z6[23] = (~(Xamnv6 ^ Alf7z6[23]));
assign Jjg7z6[22] = (~(Xamnv6 ^ Alf7z6[22]));
assign Jjg7z6[21] = (~(Xamnv6 ^ Alf7z6[21]));
assign Jjg7z6[20] = (~(Xamnv6 ^ Alf7z6[20]));
assign Jjg7z6[1] = (~(Xamnv6 ^ Alf7z6[1]));
assign Jjg7z6[19] = (~(Xamnv6 ^ Alf7z6[19]));
assign Jjg7z6[18] = (~(Xamnv6 ^ Alf7z6[18]));
assign Jjg7z6[17] = (~(Xamnv6 ^ Alf7z6[17]));
assign Jjg7z6[16] = (Wvl8v6 ^ Alf7z6[16]);
assign Jjg7z6[15] = (~(Xamnv6 ^ Alf7z6[15]));
assign Jjg7z6[14] = (Wvl8v6 ^ Alf7z6[14]);
assign Jjg7z6[13] = (Wvl8v6 ^ Alf7z6[13]);
assign Jjg7z6[12] = (~(Xamnv6 ^ Alf7z6[12]));
assign Jjg7z6[11] = (~(Xamnv6 ^ Alf7z6[11]));
assign Xamnv6 = (!Wvl8v6);
assign Jjg7z6[10] = (Wvl8v6 ^ Alf7z6[10]);
assign Dqg7z6[9] = (~(Alf7z6[8] ^ Lbmnv6));
assign Dqg7z6[8] = (~(Alf7z6[7] ^ Lbmnv6));
assign Dqg7z6[7] = (~(Alf7z6[6] ^ Lbmnv6));
assign Dqg7z6[6] = (~(Alf7z6[5] ^ Lbmnv6));
assign Dqg7z6[5] = (~(Alf7z6[4] ^ Lbmnv6));
assign Dqg7z6[4] = (~(Alf7z6[3] ^ Lbmnv6));
assign Dqg7z6[3] = (~(Alf7z6[2] ^ Lbmnv6));
assign Dqg7z6[32] = (Ebmnv6 ^ Lbmnv6);
assign Dqg7z6[31] = (Alf7z6[30] ^ Geo7v6);
assign Dqg7z6[30] = (~(Alf7z6[29] ^ Lbmnv6));
assign Dqg7z6[2] = (~(Alf7z6[1] ^ Lbmnv6));
assign Dqg7z6[29] = (~(Alf7z6[28] ^ Lbmnv6));
assign Dqg7z6[28] = (~(Alf7z6[27] ^ Lbmnv6));
assign Dqg7z6[27] = (~(Alf7z6[26] ^ Lbmnv6));
assign Dqg7z6[26] = (~(Alf7z6[25] ^ Lbmnv6));
assign Dqg7z6[25] = (~(Alf7z6[24] ^ Lbmnv6));
assign Dqg7z6[24] = (~(Alf7z6[23] ^ Lbmnv6));
assign Dqg7z6[23] = (~(Alf7z6[22] ^ Lbmnv6));
assign Dqg7z6[22] = (~(Alf7z6[21] ^ Lbmnv6));
assign Dqg7z6[21] = (~(Alf7z6[20] ^ Lbmnv6));
assign Dqg7z6[20] = (~(Alf7z6[19] ^ Lbmnv6));
assign Dqg7z6[1] = (Alf7z6[0] ^ Geo7v6);
assign Dqg7z6[19] = (~(Alf7z6[18] ^ Lbmnv6));
assign Dqg7z6[18] = (~(Alf7z6[17] ^ Lbmnv6));
assign Dqg7z6[17] = (Alf7z6[16] ^ Geo7v6);
assign Dqg7z6[16] = (~(Alf7z6[15] ^ Lbmnv6));
assign Dqg7z6[15] = (Alf7z6[14] ^ Geo7v6);
assign Dqg7z6[14] = (Alf7z6[13] ^ Geo7v6);
assign Dqg7z6[13] = (~(Alf7z6[12] ^ Lbmnv6));
assign Lbmnv6 = (!Geo7v6);
assign Dqg7z6[12] = (Alf7z6[11] ^ Geo7v6);
assign Dqg7z6[11] = (Alf7z6[10] ^ Geo7v6);
assign Dqg7z6[10] = (Alf7z6[9] ^ Geo7v6);
assign Ssf7z6[9] = (Alf7z6[25] & Sbmnv6);
assign Ssf7z6[8] = (Alf7z6[24] & Sbmnv6);
assign Ssf7z6[7] = (Alf7z6[23] & Sbmnv6);
assign Ssf7z6[6] = (Alf7z6[22] & Sbmnv6);
assign Ssf7z6[5] = (Alf7z6[21] & Sbmnv6);
assign Ssf7z6[4] = (Alf7z6[20] & Sbmnv6);
assign Ssf7z6[3] = (Alf7z6[19] & Sbmnv6);
assign Ssf7z6[2] = (Alf7z6[18] & Sbmnv6);
assign Ssf7z6[1] = (Alf7z6[17] & Sbmnv6);
assign Ssf7z6[15] = (Alf7z6[31] & Sbmnv6);
assign Ssf7z6[14] = (Alf7z6[30] & Sbmnv6);
assign Ssf7z6[13] = (Alf7z6[29] & Sbmnv6);
assign Ssf7z6[12] = (Alf7z6[28] & Sbmnv6);
assign Ssf7z6[11] = (Alf7z6[27] & Sbmnv6);
assign Ssf7z6[10] = (Alf7z6[26] & Sbmnv6);
assign Ssf7z6[0] = (Alf7z6[16] & Sbmnv6);
assign Ivf7z6[9] = (Yxf7z6[25] & Zbmnv6);
assign Ivf7z6[8] = (Yxf7z6[24] & Zbmnv6);
assign Ivf7z6[7] = (Yxf7z6[23] & Zbmnv6);
assign Ivf7z6[6] = (Yxf7z6[22] & Zbmnv6);
assign Ivf7z6[5] = (Yxf7z6[21] & Zbmnv6);
assign Ivf7z6[4] = (Yxf7z6[20] & Zbmnv6);
assign Ivf7z6[3] = (Yxf7z6[19] & Zbmnv6);
assign Ivf7z6[2] = (Yxf7z6[18] & Zbmnv6);
assign Ivf7z6[1] = (Yxf7z6[17] & Zbmnv6);
assign Ivf7z6[15] = (Yxf7z6[31] & Zbmnv6);
assign Ivf7z6[14] = (Yxf7z6[30] & Zbmnv6);
assign Ivf7z6[13] = (Yxf7z6[29] & Zbmnv6);
assign Ivf7z6[12] = (Yxf7z6[28] & Zbmnv6);
assign Ivf7z6[11] = (Yxf7z6[27] & Zbmnv6);
assign Ivf7z6[10] = (Yxf7z6[26] & Zbmnv6);
assign Ivf7z6[0] = (Yxf7z6[16] & Zbmnv6);
assign Hqidt6 = (L0g7z6[32] & Sbmnv6);
assign Sbmnv6 = (Zbmnv6 | Gcmnv6);
assign V7g7z6[9] = (~(Ncmnv6 & Ucmnv6));
assign Ucmnv6 = (~(S7f7z6[4] & Fhc7z6[25]));
assign Ncmnv6 = (~(S7f7z6[3] & Fhc7z6[9]));
assign V7g7z6[8] = (~(Bdmnv6 & Idmnv6));
assign Idmnv6 = (~(S7f7z6[4] & Fhc7z6[24]));
assign Bdmnv6 = (~(S7f7z6[3] & Fhc7z6[8]));
assign V7g7z6[7] = (~(Pdmnv6 & Wdmnv6));
assign Wdmnv6 = (~(S7f7z6[4] & Fhc7z6[23]));
assign Pdmnv6 = (~(S7f7z6[3] & Fhc7z6[7]));
assign V7g7z6[6] = (~(Demnv6 & Kemnv6));
assign Kemnv6 = (~(S7f7z6[4] & Fhc7z6[22]));
assign Demnv6 = (~(S7f7z6[3] & Fhc7z6[6]));
assign V7g7z6[5] = (~(Remnv6 & Yemnv6));
assign Yemnv6 = (~(S7f7z6[4] & Fhc7z6[21]));
assign Remnv6 = (~(S7f7z6[3] & Fhc7z6[5]));
assign V7g7z6[4] = (~(Ffmnv6 & Mfmnv6));
assign Mfmnv6 = (~(S7f7z6[3] & E3c7z6[4]));
assign Ffmnv6 = (~(S7f7z6[4] & Fhc7z6[20]));
assign V7g7z6[3] = (~(Tfmnv6 & Agmnv6));
assign Agmnv6 = (~(S7f7z6[3] & E3c7z6[3]));
assign Tfmnv6 = (~(S7f7z6[4] & Fhc7z6[19]));
assign V7g7z6[31] = (S7f7z6[5] & Fhc7z6[31]);
assign V7g7z6[30] = (S7f7z6[5] & Fhc7z6[30]);
assign V7g7z6[2] = (~(Hgmnv6 & Ogmnv6));
assign Ogmnv6 = (~(S7f7z6[3] & E3c7z6[2]));
assign Hgmnv6 = (~(S7f7z6[4] & Fhc7z6[18]));
assign V7g7z6[29] = (S7f7z6[5] & Fhc7z6[29]);
assign V7g7z6[28] = (S7f7z6[5] & Fhc7z6[28]);
assign V7g7z6[27] = (S7f7z6[5] & Fhc7z6[27]);
assign V7g7z6[26] = (S7f7z6[5] & Fhc7z6[26]);
assign V7g7z6[25] = (S7f7z6[5] & Fhc7z6[25]);
assign V7g7z6[24] = (S7f7z6[5] & Fhc7z6[24]);
assign V7g7z6[23] = (S7f7z6[5] & Fhc7z6[23]);
assign V7g7z6[22] = (S7f7z6[5] & Fhc7z6[22]);
assign V7g7z6[21] = (S7f7z6[5] & Fhc7z6[21]);
assign V7g7z6[20] = (S7f7z6[5] & Fhc7z6[20]);
assign V7g7z6[1] = (~(Vgmnv6 & Chmnv6));
assign Chmnv6 = (~(S7f7z6[3] & E3c7z6[1]));
assign Vgmnv6 = (~(S7f7z6[4] & Fhc7z6[17]));
assign V7g7z6[19] = (S7f7z6[5] & Fhc7z6[19]);
assign V7g7z6[18] = (S7f7z6[5] & Fhc7z6[18]);
assign V7g7z6[17] = (S7f7z6[5] & Fhc7z6[17]);
assign V7g7z6[16] = (S7f7z6[5] & Fhc7z6[16]);
assign V7g7z6[15] = (~(Jhmnv6 & Qhmnv6));
assign Qhmnv6 = (~(S7f7z6[3] & Fhc7z6[15]));
assign Jhmnv6 = (~(S7f7z6[4] & Fhc7z6[31]));
assign V7g7z6[14] = (~(Xhmnv6 & Eimnv6));
assign Eimnv6 = (~(S7f7z6[3] & Fhc7z6[14]));
assign Xhmnv6 = (~(S7f7z6[4] & Fhc7z6[30]));
assign V7g7z6[13] = (~(Limnv6 & Simnv6));
assign Simnv6 = (~(S7f7z6[3] & Fhc7z6[13]));
assign Limnv6 = (~(S7f7z6[4] & Fhc7z6[29]));
assign V7g7z6[12] = (~(Zimnv6 & Gjmnv6));
assign Gjmnv6 = (~(S7f7z6[3] & Fhc7z6[12]));
assign Zimnv6 = (~(S7f7z6[4] & Fhc7z6[28]));
assign V7g7z6[11] = (~(Njmnv6 & Ujmnv6));
assign Ujmnv6 = (~(S7f7z6[3] & Fhc7z6[11]));
assign Njmnv6 = (~(S7f7z6[4] & Fhc7z6[27]));
assign V7g7z6[10] = (~(Bkmnv6 & Ikmnv6));
assign Ikmnv6 = (~(S7f7z6[3] & Fhc7z6[10]));
assign Bkmnv6 = (~(S7f7z6[4] & Fhc7z6[26]));
assign V7g7z6[0] = (~(Pkmnv6 & Wkmnv6));
assign Wkmnv6 = (~(S7f7z6[3] & E3c7z6[0]));
assign Pkmnv6 = (~(S7f7z6[4] & Fhc7z6[16]));
assign Fag7z6[9] = (~(Dlmnv6 & Klmnv6));
assign Klmnv6 = (~(S7f7z6[1] & Kxb7z6[25]));
assign Dlmnv6 = (~(S7f7z6[0] & Kxb7z6[9]));
assign Fag7z6[8] = (~(Rlmnv6 & Ylmnv6));
assign Ylmnv6 = (~(S7f7z6[1] & Kxb7z6[24]));
assign Rlmnv6 = (~(S7f7z6[0] & Kxb7z6[8]));
assign Fag7z6[7] = (~(Fmmnv6 & Mmmnv6));
assign Mmmnv6 = (~(S7f7z6[1] & Kxb7z6[23]));
assign Fmmnv6 = (~(S7f7z6[0] & Kxb7z6[7]));
assign Fag7z6[6] = (~(Tmmnv6 & Anmnv6));
assign Anmnv6 = (~(S7f7z6[1] & Kxb7z6[22]));
assign Tmmnv6 = (~(S7f7z6[0] & Kxb7z6[6]));
assign Fag7z6[5] = (~(Hnmnv6 & Onmnv6));
assign Onmnv6 = (~(S7f7z6[1] & Kxb7z6[21]));
assign Hnmnv6 = (~(S7f7z6[0] & Kxb7z6[5]));
assign Fag7z6[4] = (~(Vnmnv6 & Comnv6));
assign Comnv6 = (~(S7f7z6[1] & Kxb7z6[20]));
assign Vnmnv6 = (~(S7f7z6[0] & Kxb7z6[4]));
assign Fag7z6[3] = (~(Jomnv6 & Qomnv6));
assign Qomnv6 = (~(S7f7z6[1] & Kxb7z6[19]));
assign Jomnv6 = (~(S7f7z6[0] & Kxb7z6[3]));
assign Fag7z6[31] = (S7f7z6[2] & Kxb7z6[31]);
assign Fag7z6[30] = (S7f7z6[2] & Kxb7z6[30]);
assign Fag7z6[2] = (~(Xomnv6 & Epmnv6));
assign Epmnv6 = (~(S7f7z6[1] & Kxb7z6[18]));
assign Xomnv6 = (~(S7f7z6[0] & Kxb7z6[2]));
assign Fag7z6[29] = (S7f7z6[2] & Kxb7z6[29]);
assign Fag7z6[28] = (S7f7z6[2] & Kxb7z6[28]);
assign Fag7z6[27] = (S7f7z6[2] & Kxb7z6[27]);
assign Fag7z6[26] = (S7f7z6[2] & Kxb7z6[26]);
assign Fag7z6[25] = (S7f7z6[2] & Kxb7z6[25]);
assign Fag7z6[24] = (S7f7z6[2] & Kxb7z6[24]);
assign Fag7z6[23] = (S7f7z6[2] & Kxb7z6[23]);
assign Fag7z6[22] = (S7f7z6[2] & Kxb7z6[22]);
assign Fag7z6[21] = (S7f7z6[2] & Kxb7z6[21]);
assign Fag7z6[20] = (S7f7z6[2] & Kxb7z6[20]);
assign Fag7z6[1] = (~(Lpmnv6 & Spmnv6));
assign Spmnv6 = (~(S7f7z6[1] & Kxb7z6[17]));
assign Lpmnv6 = (~(S7f7z6[0] & Kxb7z6[1]));
assign Fag7z6[19] = (S7f7z6[2] & Kxb7z6[19]);
assign Fag7z6[18] = (S7f7z6[2] & Kxb7z6[18]);
assign Fag7z6[17] = (S7f7z6[2] & Kxb7z6[17]);
assign Fag7z6[16] = (S7f7z6[2] & Kxb7z6[16]);
assign Fag7z6[15] = (~(Zpmnv6 & Gqmnv6));
assign Gqmnv6 = (~(S7f7z6[0] & Kxb7z6[15]));
assign Zpmnv6 = (~(S7f7z6[1] & Kxb7z6[31]));
assign Fag7z6[14] = (~(Nqmnv6 & Uqmnv6));
assign Uqmnv6 = (~(S7f7z6[0] & Kxb7z6[14]));
assign Nqmnv6 = (~(S7f7z6[1] & Kxb7z6[30]));
assign Fag7z6[13] = (~(Brmnv6 & Irmnv6));
assign Irmnv6 = (~(S7f7z6[0] & Kxb7z6[13]));
assign Brmnv6 = (~(S7f7z6[1] & Kxb7z6[29]));
assign Fag7z6[12] = (~(Prmnv6 & Wrmnv6));
assign Wrmnv6 = (~(S7f7z6[0] & Kxb7z6[12]));
assign Prmnv6 = (~(S7f7z6[1] & Kxb7z6[28]));
assign Fag7z6[11] = (~(Dsmnv6 & Ksmnv6));
assign Ksmnv6 = (~(S7f7z6[0] & Kxb7z6[11]));
assign Dsmnv6 = (~(S7f7z6[1] & Kxb7z6[27]));
assign Fag7z6[10] = (~(Rsmnv6 & Ysmnv6));
assign Ysmnv6 = (~(S7f7z6[0] & Kxb7z6[10]));
assign Rsmnv6 = (~(S7f7z6[1] & Kxb7z6[26]));
assign Fag7z6[0] = (~(Ftmnv6 & Mtmnv6));
assign Mtmnv6 = (~(S7f7z6[0] & Kxb7z6[0]));
assign Ftmnv6 = (~(S7f7z6[1] & Kxb7z6[16]));
assign Kif7z6[9] = (X2g7z6[9] ^ J5g7z6[9]);
assign Kif7z6[8] = (X2g7z6[8] ^ J5g7z6[8]);
assign Kif7z6[7] = (X2g7z6[7] ^ J5g7z6[7]);
assign Kif7z6[6] = (X2g7z6[6] ^ J5g7z6[6]);
assign Kif7z6[5] = (X2g7z6[5] ^ J5g7z6[5]);
assign Kif7z6[4] = (X2g7z6[4] ^ J5g7z6[4]);
assign Kif7z6[3] = (X2g7z6[3] ^ J5g7z6[3]);
assign Kif7z6[31] = (X2g7z6[31] ^ J5g7z6[31]);
assign Kif7z6[30] = (X2g7z6[30] ^ J5g7z6[30]);
assign Kif7z6[2] = (X2g7z6[2] ^ J5g7z6[2]);
assign Kif7z6[29] = (X2g7z6[29] ^ J5g7z6[29]);
assign Kif7z6[28] = (X2g7z6[28] ^ J5g7z6[28]);
assign Kif7z6[27] = (X2g7z6[27] ^ J5g7z6[27]);
assign Kif7z6[26] = (X2g7z6[26] ^ J5g7z6[26]);
assign Kif7z6[25] = (X2g7z6[25] ^ J5g7z6[25]);
assign Kif7z6[24] = (X2g7z6[24] ^ J5g7z6[24]);
assign Kif7z6[23] = (X2g7z6[23] ^ J5g7z6[23]);
assign Kif7z6[22] = (X2g7z6[22] ^ J5g7z6[22]);
assign Kif7z6[21] = (X2g7z6[21] ^ J5g7z6[21]);
assign Kif7z6[20] = (X2g7z6[20] ^ J5g7z6[20]);
assign Kif7z6[1] = (X2g7z6[1] ^ J5g7z6[1]);
assign Kif7z6[19] = (X2g7z6[19] ^ J5g7z6[19]);
assign Kif7z6[18] = (X2g7z6[18] ^ J5g7z6[18]);
assign Kif7z6[17] = (X2g7z6[17] ^ J5g7z6[17]);
assign Kif7z6[16] = (X2g7z6[16] ^ J5g7z6[16]);
assign Kif7z6[15] = (X2g7z6[15] ^ J5g7z6[15]);
assign Kif7z6[14] = (X2g7z6[14] ^ J5g7z6[14]);
assign Kif7z6[13] = (X2g7z6[13] ^ J5g7z6[13]);
assign Kif7z6[12] = (X2g7z6[12] ^ J5g7z6[12]);
assign Kif7z6[11] = (X2g7z6[11] ^ J5g7z6[11]);
assign Kif7z6[10] = (X2g7z6[10] ^ J5g7z6[10]);
assign Kif7z6[0] = (X2g7z6[0] ^ J5g7z6[0]);
assign Uff7z6[9] = (X2g7z6[9] | J5g7z6[9]);
assign J5g7z6[9] = (Ttmnv6 & Aumnv6);
assign X2g7z6[9] = (~(Humnv6 | Oumnv6));
assign Uff7z6[8] = (X2g7z6[8] | J5g7z6[8]);
assign J5g7z6[8] = (Vumnv6 & Aumnv6);
assign X2g7z6[8] = (~(Cvmnv6 | Oumnv6));
assign Uff7z6[7] = (X2g7z6[7] | J5g7z6[7]);
assign J5g7z6[7] = (Jvmnv6 & Aumnv6);
assign X2g7z6[7] = (~(Qvmnv6 | Oumnv6));
assign Uff7z6[6] = (X2g7z6[6] | J5g7z6[6]);
assign J5g7z6[6] = (Xvmnv6 & Aumnv6);
assign X2g7z6[6] = (~(Ewmnv6 | Oumnv6));
assign Uff7z6[5] = (X2g7z6[5] | J5g7z6[5]);
assign J5g7z6[5] = (Lwmnv6 & Aumnv6);
assign X2g7z6[5] = (~(Swmnv6 | Oumnv6));
assign Uff7z6[4] = (X2g7z6[4] | J5g7z6[4]);
assign J5g7z6[4] = (Zwmnv6 & Aumnv6);
assign X2g7z6[4] = (~(Gxmnv6 | Oumnv6));
assign Uff7z6[3] = (X2g7z6[3] | J5g7z6[3]);
assign J5g7z6[3] = (Nxmnv6 & Aumnv6);
assign X2g7z6[3] = (~(Uxmnv6 | Oumnv6));
assign Uff7z6[30] = (X2g7z6[30] | J5g7z6[30]);
assign J5g7z6[30] = (Bymnv6 & Aumnv6);
assign X2g7z6[30] = (~(Iymnv6 | Oumnv6));
assign Uff7z6[2] = (X2g7z6[2] | J5g7z6[2]);
assign J5g7z6[2] = (Pymnv6 & Aumnv6);
assign X2g7z6[2] = (~(Wymnv6 | Oumnv6));
assign Uff7z6[29] = (X2g7z6[29] | J5g7z6[29]);
assign J5g7z6[29] = (Dzmnv6 & Aumnv6);
assign X2g7z6[29] = (~(Kzmnv6 | Oumnv6));
assign Uff7z6[28] = (X2g7z6[28] | J5g7z6[28]);
assign J5g7z6[28] = (Rzmnv6 & Aumnv6);
assign X2g7z6[28] = (~(Yzmnv6 | Oumnv6));
assign Uff7z6[27] = (X2g7z6[27] | J5g7z6[27]);
assign J5g7z6[27] = (F0nnv6 & Aumnv6);
assign X2g7z6[27] = (~(M0nnv6 | Oumnv6));
assign Uff7z6[26] = (X2g7z6[26] | J5g7z6[26]);
assign J5g7z6[26] = (T0nnv6 & Aumnv6);
assign X2g7z6[26] = (~(A1nnv6 | Oumnv6));
assign Uff7z6[25] = (X2g7z6[25] | J5g7z6[25]);
assign J5g7z6[25] = (H1nnv6 & Aumnv6);
assign X2g7z6[25] = (~(O1nnv6 | Oumnv6));
assign Uff7z6[24] = (X2g7z6[24] | J5g7z6[24]);
assign J5g7z6[24] = (V1nnv6 & Aumnv6);
assign X2g7z6[24] = (~(C2nnv6 | Oumnv6));
assign Uff7z6[23] = (X2g7z6[23] | J5g7z6[23]);
assign J5g7z6[23] = (J2nnv6 & Aumnv6);
assign X2g7z6[23] = (~(Q2nnv6 | Oumnv6));
assign Uff7z6[22] = (X2g7z6[22] | J5g7z6[22]);
assign J5g7z6[22] = (X2nnv6 & Aumnv6);
assign X2g7z6[22] = (~(E3nnv6 | Oumnv6));
assign Uff7z6[21] = (X2g7z6[21] | J5g7z6[21]);
assign J5g7z6[21] = (L3nnv6 & Aumnv6);
assign X2g7z6[21] = (~(S3nnv6 | Oumnv6));
assign Uff7z6[20] = (X2g7z6[20] | J5g7z6[20]);
assign J5g7z6[20] = (Z3nnv6 & Aumnv6);
assign X2g7z6[20] = (~(G4nnv6 | Oumnv6));
assign Uff7z6[1] = (X2g7z6[1] | J5g7z6[1]);
assign J5g7z6[1] = (N4nnv6 & Aumnv6);
assign X2g7z6[1] = (~(U4nnv6 | Oumnv6));
assign Uff7z6[19] = (X2g7z6[19] | J5g7z6[19]);
assign J5g7z6[19] = (B5nnv6 & Aumnv6);
assign X2g7z6[19] = (~(I5nnv6 | Oumnv6));
assign Uff7z6[18] = (X2g7z6[18] | J5g7z6[18]);
assign J5g7z6[18] = (P5nnv6 & Aumnv6);
assign X2g7z6[18] = (~(W5nnv6 | Oumnv6));
assign Uff7z6[17] = (X2g7z6[17] | J5g7z6[17]);
assign J5g7z6[17] = (D6nnv6 & Aumnv6);
assign X2g7z6[17] = (~(K6nnv6 | Oumnv6));
assign Uff7z6[16] = (X2g7z6[16] | J5g7z6[16]);
assign J5g7z6[16] = (R6nnv6 & Aumnv6);
assign X2g7z6[16] = (~(Y6nnv6 | Oumnv6));
assign Uff7z6[15] = (X2g7z6[15] | J5g7z6[15]);
assign J5g7z6[15] = (F7nnv6 & Aumnv6);
assign X2g7z6[15] = (~(M7nnv6 | Oumnv6));
assign Uff7z6[14] = (X2g7z6[14] | J5g7z6[14]);
assign J5g7z6[14] = (T7nnv6 & Aumnv6);
assign X2g7z6[14] = (~(A8nnv6 | Oumnv6));
assign Uff7z6[13] = (X2g7z6[13] | J5g7z6[13]);
assign J5g7z6[13] = (H8nnv6 & Aumnv6);
assign X2g7z6[13] = (~(O8nnv6 | Oumnv6));
assign Uff7z6[12] = (X2g7z6[12] | J5g7z6[12]);
assign J5g7z6[12] = (V8nnv6 & Aumnv6);
assign X2g7z6[12] = (~(C9nnv6 | Oumnv6));
assign Uff7z6[11] = (X2g7z6[11] | J5g7z6[11]);
assign J5g7z6[11] = (J9nnv6 & Aumnv6);
assign X2g7z6[11] = (~(Q9nnv6 | Oumnv6));
assign Uff7z6[10] = (X2g7z6[10] | J5g7z6[10]);
assign J5g7z6[10] = (X9nnv6 & Aumnv6);
assign X2g7z6[10] = (~(Eannv6 | Oumnv6));
assign Uff7z6[0] = (X2g7z6[0] | J5g7z6[0]);
assign J5g7z6[0] = (~(Lannv6 | Sannv6));
assign X2g7z6[0] = (Zannv6 & Gbnnv6);
assign Arkdt6 = (~(Nbnnv6 & Ubnnv6));
assign Ubnnv6 = (~(Bcnnv6 & Gbnnv6));
assign Bcnnv6 = (~(Icnnv6 & Pcnnv6));
assign Pcnnv6 = (~(D7hdt6 & Wcnnv6));
assign Icnnv6 = (~(Dte7z6[20] & S7gdt6));
assign Nbnnv6 = (~(Ddnnv6 & Kdnnv6));
assign Kdnnv6 = (~(Dte7z6[20] & Rdnnv6));
assign Ddnnv6 = (~(Ydnnv6 | Fennv6));
assign Ydnnv6 = (Mennv6 & Tennv6);
assign Jaf7z6[5] = (~(Afnnv6 & Hfnnv6));
assign Afnnv6 = (~(Ofnnv6 & Vfnnv6));
assign Vfnnv6 = (~(Q9hdt6 & Mrbdt6));
assign Jaf7z6[4] = (Cgnnv6 & Jgnnv6);
assign Jaf7z6[3] = (Qgnnv6 & Jgnnv6);
assign Jaf7z6[2] = (Xgnnv6 & Jgnnv6);
assign Jaf7z6[1] = (Ehnnv6 & Jgnnv6);
assign Jaf7z6[0] = (Lhnnv6 & Jgnnv6);
assign Jgnnv6 = (~(Shnnv6 & Zhnnv6));
assign Zhnnv6 = (~(Ginnv6 & Ofnnv6));
assign Ginnv6 = (Q9hdt6 & Mrbdt6);
assign Shnnv6 = (Ninnv6 & Uinnv6);
assign Rze7z6[5] = (Bjnnv6 & Ijnnv6);
assign Rze7z6[4] = (Ijnnv6 & Pjnnv6);
assign Rze7z6[3] = (Ijnnv6 & Wjnnv6);
assign Rze7z6[2] = (Ijnnv6 & Dknnv6);
assign Rze7z6[1] = (Ijnnv6 & Kknnv6);
assign Rze7z6[0] = (Ijnnv6 & Rknnv6);
assign K2f7z6[5] = (D5f7z6[5] & Ijnnv6);
assign K2f7z6[4] = (D5f7z6[4] & Ijnnv6);
assign K2f7z6[3] = (D5f7z6[3] & Ijnnv6);
assign K2f7z6[2] = (D5f7z6[2] & Ijnnv6);
assign K2f7z6[1] = (D5f7z6[1] & Ijnnv6);
assign K2f7z6[0] = (D5f7z6[0] & Ijnnv6);
assign Flc7z6[9] = (~(Yknnv6 & Flnnv6));
assign Yknnv6 = (Mlnnv6 & Tlnnv6);
assign Tlnnv6 = (~(Zec7z6[24] & Amnnv6));
assign Flc7z6[8] = (~(Hmnnv6 & Omnnv6));
assign Omnnv6 = (~(Zec7z6[23] & Amnnv6));
assign Hmnnv6 = (~(Zec7z6[7] & Vmnnv6));
assign Flc7z6[7] = (~(Cnnnv6 & Jnnnv6));
assign Jnnnv6 = (~(Zec7z6[22] & Amnnv6));
assign Cnnnv6 = (~(Zec7z6[6] & Vmnnv6));
assign Flc7z6[6] = (~(Qnnnv6 & Xnnnv6));
assign Xnnnv6 = (~(Zec7z6[21] & Amnnv6));
assign Qnnnv6 = (~(Zec7z6[5] & Vmnnv6));
assign Flc7z6[5] = (~(Eonnv6 & Lonnv6));
assign Lonnv6 = (~(Zec7z6[20] & Amnnv6));
assign Eonnv6 = (~(Zec7z6[4] & Vmnnv6));
assign Flc7z6[4] = (~(Sonnv6 & Zonnv6));
assign Zonnv6 = (~(Zec7z6[19] & Amnnv6));
assign Sonnv6 = (~(Zec7z6[3] & Vmnnv6));
assign Flc7z6[3] = (~(Gpnnv6 & Npnnv6));
assign Npnnv6 = (~(Zec7z6[18] & Amnnv6));
assign Gpnnv6 = (~(Zec7z6[2] & Vmnnv6));
assign Flc7z6[31] = (~(Upnnv6 & Bqnnv6));
assign Bqnnv6 = (~(Zec7z6[10] & Amnnv6));
assign Flc7z6[2] = (~(Iqnnv6 & Pqnnv6));
assign Pqnnv6 = (~(Zec7z6[17] & Amnnv6));
assign Iqnnv6 = (~(Zec7z6[1] & Vmnnv6));
assign Flc7z6[23] = (~(Wqnnv6 & Drnnv6));
assign Drnnv6 = (~(Krnnv6 & Rrnnv6));
assign Krnnv6 = (Zec7z6[10] ^ Yrnnv6);
assign Yrnnv6 = (!Zec7z6[29]);
assign Flc7z6[22] = (~(Wqnnv6 & Fsnnv6));
assign Fsnnv6 = (~(Msnnv6 & Rrnnv6));
assign Flc7z6[21] = (~(Wqnnv6 & Tsnnv6));
assign Tsnnv6 = (~(Rrnnv6 & Zec7z6[9]));
assign Flc7z6[20] = (~(Wqnnv6 & Atnnv6));
assign Atnnv6 = (~(Rrnnv6 & Zec7z6[8]));
assign Wqnnv6 = (Upnnv6 & Htnnv6);
assign Flc7z6[1] = (~(Otnnv6 & Vtnnv6));
assign Vtnnv6 = (~(Zec7z6[16] & Amnnv6));
assign Otnnv6 = (~(Zec7z6[0] & Vmnnv6));
assign Flc7z6[19] = (~(Cunnv6 & Upnnv6));
assign Cunnv6 = (Junnv6 & Qunnv6);
assign Qunnv6 = (~(Rrnnv6 & Zec7z6[7]));
assign Junnv6 = (~(Nginv6 & Zec7z6[27]));
assign Flc7z6[18] = (~(Xunnv6 & Upnnv6));
assign Xunnv6 = (Evnnv6 & Lvnnv6);
assign Lvnnv6 = (~(Rrnnv6 & Zec7z6[6]));
assign Evnnv6 = (~(Nginv6 & Zec7z6[29]));
assign Flc7z6[17] = (~(Upnnv6 & Svnnv6));
assign Svnnv6 = (~(Zec7z6[5] & Amnnv6));
assign Flc7z6[16] = (~(Upnnv6 & Zvnnv6));
assign Zvnnv6 = (~(Zec7z6[4] & Amnnv6));
assign Flc7z6[15] = (~(Upnnv6 & Gwnnv6));
assign Gwnnv6 = (~(Zec7z6[3] & Amnnv6));
assign Flc7z6[14] = (~(Upnnv6 & Nwnnv6));
assign Nwnnv6 = (~(Zec7z6[2] & Amnnv6));
assign Flc7z6[13] = (~(Upnnv6 & Uwnnv6));
assign Uwnnv6 = (~(Zec7z6[1] & Amnnv6));
assign Flc7z6[12] = (~(Upnnv6 & Bxnnv6));
assign Bxnnv6 = (~(Zec7z6[0] & Amnnv6));
assign Flc7z6[11] = (~(Upnnv6 & Ixnnv6));
assign Ixnnv6 = (~(Zec7z6[26] & Amnnv6));
assign Upnnv6 = (Flnnv6 & Pxnnv6);
assign Flc7z6[10] = (~(Wxnnv6 & Flnnv6));
assign Wxnnv6 = (Dynnv6 & Kynnv6);
assign Kynnv6 = (~(Zec7z6[25] & Amnnv6));
assign Axbdt6 = (Rynnv6 & Yynnv6);
assign Yynnv6 = (Fznnv6 & Mznnv6);
assign Mznnv6 = (~(Icy7v6 | Bdi8v6));
assign Fznnv6 = (~(Tznnv6 | A0onv6));
assign Rynnv6 = (H0onv6 & O0onv6);
assign O0onv6 = (~(V0onv6 | C1onv6));
assign H0onv6 = (Oaadt6 & J1onv6);
assign J1onv6 = (~(Q1onv6 & X1onv6));
assign X1onv6 = (~(E2onv6 & L2onv6));
assign L2onv6 = (Lybdt6 & S2onv6);
assign E2onv6 = (Z2onv6 & G3onv6);
assign Q1onv6 = (~(N3onv6 & U3onv6));
assign U3onv6 = (~(B4onv6 & I4onv6));
assign I4onv6 = (P4onv6 & W4onv6);
assign P4onv6 = (~(D5onv6 & K5onv6));
assign D5onv6 = (~(R5onv6 & Y5onv6));
assign Y5onv6 = (F6onv6 & M6onv6);
assign F6onv6 = (T6onv6 & A7onv6);
assign R5onv6 = (H7onv6 & O7onv6);
assign H7onv6 = (V7onv6 & C8onv6);
assign V7onv6 = (~(J8onv6 & Q8onv6));
assign J8onv6 = (X8onv6 & E9onv6);
assign B4onv6 = (L9onv6 & S9onv6);
assign S9onv6 = (~(Z9onv6 & Gaonv6));
assign O7o7z6[1] = (Pl0ft6 & Naonv6);
assign HMASTERS[1] = (~(Uaonv6 | Bbonv6));
assign HMASTERD[1] = (~(Ibonv6 | Bbonv6));
assign Bbonv6 = (~(Pbonv6 & Xnnet6));
assign L3oet6 = (Wbonv6 & Dconv6);
assign Wbonv6 = (Kconv6 & Rconv6);
assign Pvnet6 = (Iynet6 ? Fdonv6 : Yconv6);
assign Fdonv6 = (~(Mdonv6 & Tdonv6));
assign Tdonv6 = (Aeonv6 | Qteet6);
assign Yconv6 = (Heonv6 & Oeonv6);
assign Oeonv6 = (!Veonv6);
assign Heonv6 = (Cfonv6 & Jfonv6);
assign Spnet6 = (Qfonv6 & Xfonv6);
assign Xfonv6 = (Egonv6 & Lgonv6);
assign Egonv6 = (Sgonv6 & Zgonv6);
assign Qfonv6 = (Ghonv6 & B2jnv6);
assign Ssnet6 = (Nhonv6 & Uhonv6);
assign Uhonv6 = (~(Xjh7v6 & Bionv6));
assign M7yet6 = (~(Iionv6 & Pionv6));
assign Pionv6 = (~(Wionv6 & Djonv6));
assign Wionv6 = (Znn7z6[1] & Kjonv6);
assign Iionv6 = (~(Rjonv6 & Yjonv6));
assign Rjonv6 = (~(Fkonv6 ^ Mkonv6));
assign Fkonv6 = (Tkonv6 | Alonv6);
assign Dhyet6 = (~(Hlonv6 & Olonv6));
assign Olonv6 = (~(Sjyet6 & Vlonv6));
assign Vlonv6 = (Cmonv6 | Jmonv6);
assign Hlonv6 = (!Qmonv6);
assign Dmyet6 = (Xmonv6 & Enonv6);
assign Xmonv6 = (~(Cmonv6 | Jmonv6));
assign Jmonv6 = (!Yjonv6);
assign S4yet6 = (~(Lnonv6 & Snonv6));
assign Snonv6 = (~(Znonv6 & Dkm7z6[0]));
assign Znonv6 = (HRESPD[0] & Goonv6);
assign Lnonv6 = (~(Noonv6 & HRESPS[0]));
assign Kvxet6 = (~(Uoonv6 & Bponv6));
assign Bponv6 = (~(Styet6 & Iponv6));
assign Iponv6 = (~(Pponv6 & Wponv6));
assign Wponv6 = (~(Dqonv6 & Kqonv6));
assign Pponv6 = (~(Rqonv6 & Yqonv6));
assign Uoonv6 = (Fronv6 & Mronv6);
assign Mronv6 = (~(Tronv6 & Asonv6));
assign Fronv6 = (~(Ewyet6 & Hsonv6));
assign Hsonv6 = (~(Osonv6 & Vsonv6));
assign Vsonv6 = (~(Dqonv6 & Itb7z6[8]));
assign Dqonv6 = (Ctonv6 & S7n7z6[0]);
assign Ctonv6 = (Evadt6 & Jtonv6);
assign Osonv6 = (~(Rqonv6 & Itb7z6[24]));
assign Ean7z6[4] = (Qtonv6 | Qvm7z6[1]);
assign Qvm7z6[1] = (Hjn7z6[6] & Xtonv6);
assign Xtonv6 = (Jtonv6 | S7n7z6[0]);
assign Qtonv6 = (Hjn7z6[6] ? Euonv6 : Rqonv6);
assign Rqonv6 = (Luonv6 & S7n7z6[1]);
assign Luonv6 = (~(Euonv6 | S7n7z6[0]));
assign Ean7z6[3] = (Suonv6 | Qvm7z6[0]);
assign Qvm7z6[0] = (Hjn7z6[5] & Zuonv6);
assign Suonv6 = (Evadt6 ? Gvonv6 : Hjn7z6[5]);
assign Gvonv6 = (~(Zuonv6 | Hjn7z6[5]));
assign Chn7z6[9] = (~(Nvonv6 & Uvonv6));
assign Uvonv6 = (Bwonv6 & Iwonv6);
assign Iwonv6 = (~(Pwonv6 & Cmm7z6[9]));
assign Bwonv6 = (~(Wwonv6 & HADDRI[9]));
assign Nvonv6 = (Dxonv6 & Kxonv6);
assign Kxonv6 = (~(Fvb7z6[9] & Rxonv6));
assign Dxonv6 = (~(Hjn7z6[9] & Djonv6));
assign Chn7z6[8] = (~(Yxonv6 & Fyonv6));
assign Fyonv6 = (Myonv6 & Tyonv6);
assign Tyonv6 = (~(Pwonv6 & Cmm7z6[8]));
assign Myonv6 = (~(Wwonv6 & HADDRI[8]));
assign Yxonv6 = (Azonv6 & Hzonv6);
assign Hzonv6 = (~(Fvb7z6[8] & Rxonv6));
assign Azonv6 = (~(Hjn7z6[8] & Djonv6));
assign Chn7z6[7] = (~(Ozonv6 & Vzonv6));
assign Vzonv6 = (C0pnv6 & J0pnv6);
assign J0pnv6 = (~(Pwonv6 & Cmm7z6[7]));
assign C0pnv6 = (~(Wwonv6 & HADDRI[7]));
assign Ozonv6 = (Q0pnv6 & X0pnv6);
assign X0pnv6 = (~(Fvb7z6[7] & Rxonv6));
assign Q0pnv6 = (~(Hjn7z6[7] & Djonv6));
assign Chn7z6[6] = (~(E1pnv6 & L1pnv6));
assign L1pnv6 = (S1pnv6 & Z1pnv6);
assign Z1pnv6 = (~(Pwonv6 & Cmm7z6[6]));
assign S1pnv6 = (~(Wwonv6 & HADDRI[6]));
assign E1pnv6 = (G2pnv6 & N2pnv6);
assign N2pnv6 = (~(Fvb7z6[6] & Rxonv6));
assign G2pnv6 = (~(Hjn7z6[6] & Djonv6));
assign Chn7z6[5] = (~(U2pnv6 & B3pnv6));
assign B3pnv6 = (I3pnv6 & P3pnv6);
assign P3pnv6 = (~(Pwonv6 & Cmm7z6[5]));
assign I3pnv6 = (~(Wwonv6 & HADDRI[5]));
assign U2pnv6 = (W3pnv6 & D4pnv6);
assign D4pnv6 = (~(Fvb7z6[5] & Rxonv6));
assign W3pnv6 = (~(Hjn7z6[5] & Djonv6));
assign Chn7z6[4] = (~(K4pnv6 & R4pnv6));
assign R4pnv6 = (Y4pnv6 & F5pnv6);
assign F5pnv6 = (~(Pwonv6 & Cmm7z6[4]));
assign Y4pnv6 = (~(Wwonv6 & HADDRI[4]));
assign K4pnv6 = (M5pnv6 & T5pnv6);
assign T5pnv6 = (~(Fvb7z6[4] & Rxonv6));
assign M5pnv6 = (~(Ryyet6 & Djonv6));
assign Chn7z6[3] = (~(A6pnv6 & H6pnv6));
assign H6pnv6 = (O6pnv6 & V6pnv6);
assign V6pnv6 = (~(Pwonv6 & Cmm7z6[3]));
assign O6pnv6 = (~(Wwonv6 & HADDRI[3]));
assign A6pnv6 = (C7pnv6 & J7pnv6);
assign J7pnv6 = (~(Fvb7z6[3] & Rxonv6));
assign C7pnv6 = (~(S0zet6 & Djonv6));
assign Chn7z6[31] = (~(Q7pnv6 & X7pnv6));
assign X7pnv6 = (E8pnv6 & L8pnv6);
assign L8pnv6 = (~(Pwonv6 & Cmm7z6[31]));
assign E8pnv6 = (~(Wwonv6 & Njfnv6));
assign Q7pnv6 = (S8pnv6 & Z8pnv6);
assign Z8pnv6 = (~(Rxonv6 & Fvb7z6[31]));
assign S8pnv6 = (~(Hjn7z6[31] & Djonv6));
assign Chn7z6[30] = (~(G9pnv6 & N9pnv6));
assign N9pnv6 = (U9pnv6 & Bapnv6);
assign Bapnv6 = (~(Pwonv6 & Cmm7z6[30]));
assign U9pnv6 = (~(Wwonv6 & Ujfnv6));
assign G9pnv6 = (Iapnv6 & Papnv6);
assign Papnv6 = (~(Rxonv6 & Fvb7z6[30]));
assign Iapnv6 = (~(Hjn7z6[30] & Djonv6));
assign Chn7z6[2] = (~(Wapnv6 & Dbpnv6));
assign Dbpnv6 = (Kbpnv6 & Rbpnv6);
assign Rbpnv6 = (~(Pwonv6 & Yefnv6));
assign Kbpnv6 = (~(Wwonv6 & HADDRI[2]));
assign Wapnv6 = (Ybpnv6 & Fcpnv6);
assign Fcpnv6 = (~(Fvb7z6[2] & Rxonv6));
assign Ybpnv6 = (~(T2zet6 & Djonv6));
assign Chn7z6[29] = (~(Mcpnv6 & Tcpnv6));
assign Tcpnv6 = (Adpnv6 & Hdpnv6);
assign Hdpnv6 = (~(Pwonv6 & Cmm7z6[29]));
assign Adpnv6 = (~(Wwonv6 & Bkfnv6));
assign Mcpnv6 = (Odpnv6 & Vdpnv6);
assign Vdpnv6 = (~(Rxonv6 & Fvb7z6[29]));
assign Odpnv6 = (~(Hjn7z6[29] & Djonv6));
assign Chn7z6[28] = (~(Cepnv6 & Jepnv6));
assign Jepnv6 = (Qepnv6 & Xepnv6);
assign Xepnv6 = (~(Pwonv6 & Cmm7z6[28]));
assign Qepnv6 = (~(Wwonv6 & HADDRI[28]));
assign Cepnv6 = (Efpnv6 & Lfpnv6);
assign Lfpnv6 = (~(Fvb7z6[28] & Rxonv6));
assign Efpnv6 = (~(Hjn7z6[28] & Djonv6));
assign Chn7z6[27] = (~(Sfpnv6 & Zfpnv6));
assign Zfpnv6 = (Ggpnv6 & Ngpnv6);
assign Ngpnv6 = (~(Pwonv6 & Cmm7z6[27]));
assign Ggpnv6 = (~(Wwonv6 & HADDRI[27]));
assign Sfpnv6 = (Ugpnv6 & Bhpnv6);
assign Bhpnv6 = (~(Fvb7z6[27] & Rxonv6));
assign Ugpnv6 = (~(Hjn7z6[27] & Djonv6));
assign Chn7z6[26] = (~(Ihpnv6 & Phpnv6));
assign Phpnv6 = (Whpnv6 & Dipnv6);
assign Dipnv6 = (~(Pwonv6 & Cmm7z6[26]));
assign Whpnv6 = (~(Wwonv6 & HADDRI[26]));
assign Ihpnv6 = (Kipnv6 & Ripnv6);
assign Ripnv6 = (~(Fvb7z6[26] & Rxonv6));
assign Kipnv6 = (~(Hjn7z6[26] & Djonv6));
assign Chn7z6[25] = (~(Yipnv6 & Fjpnv6));
assign Fjpnv6 = (Mjpnv6 & Tjpnv6);
assign Tjpnv6 = (~(Pwonv6 & Cmm7z6[25]));
assign Mjpnv6 = (~(Wwonv6 & HADDRI[25]));
assign Yipnv6 = (Akpnv6 & Hkpnv6);
assign Hkpnv6 = (~(Rxonv6 & Fvb7z6[25]));
assign Akpnv6 = (~(Hjn7z6[25] & Djonv6));
assign Chn7z6[24] = (~(Okpnv6 & Vkpnv6));
assign Vkpnv6 = (Clpnv6 & Jlpnv6);
assign Jlpnv6 = (~(Pwonv6 & Cmm7z6[24]));
assign Clpnv6 = (~(Wwonv6 & HADDRI[24]));
assign Okpnv6 = (Qlpnv6 & Xlpnv6);
assign Xlpnv6 = (~(Fvb7z6[24] & Rxonv6));
assign Qlpnv6 = (~(Hjn7z6[24] & Djonv6));
assign Chn7z6[23] = (~(Empnv6 & Lmpnv6));
assign Lmpnv6 = (Smpnv6 & Zmpnv6);
assign Zmpnv6 = (~(Pwonv6 & Cmm7z6[23]));
assign Smpnv6 = (~(Wwonv6 & HADDRI[23]));
assign Empnv6 = (Gnpnv6 & Nnpnv6);
assign Nnpnv6 = (~(Fvb7z6[23] & Rxonv6));
assign Gnpnv6 = (~(Hjn7z6[23] & Djonv6));
assign Chn7z6[22] = (~(Unpnv6 & Bopnv6));
assign Bopnv6 = (Iopnv6 & Popnv6);
assign Popnv6 = (~(Pwonv6 & Cmm7z6[22]));
assign Iopnv6 = (~(Wwonv6 & HADDRI[22]));
assign Unpnv6 = (Wopnv6 & Dppnv6);
assign Dppnv6 = (~(Fvb7z6[22] & Rxonv6));
assign Wopnv6 = (~(Hjn7z6[22] & Djonv6));
assign Chn7z6[21] = (~(Kppnv6 & Rppnv6));
assign Rppnv6 = (Yppnv6 & Fqpnv6);
assign Fqpnv6 = (~(Pwonv6 & Cmm7z6[21]));
assign Yppnv6 = (~(Wwonv6 & HADDRI[21]));
assign Kppnv6 = (Mqpnv6 & Tqpnv6);
assign Tqpnv6 = (~(Fvb7z6[21] & Rxonv6));
assign Mqpnv6 = (~(Hjn7z6[21] & Djonv6));
assign Chn7z6[20] = (~(Arpnv6 & Hrpnv6));
assign Hrpnv6 = (Orpnv6 & Vrpnv6);
assign Vrpnv6 = (~(Pwonv6 & Cmm7z6[20]));
assign Orpnv6 = (~(Wwonv6 & HADDRI[20]));
assign Arpnv6 = (Cspnv6 & Jspnv6);
assign Jspnv6 = (~(Fvb7z6[20] & Rxonv6));
assign Cspnv6 = (~(Hjn7z6[20] & Djonv6));
assign Chn7z6[1] = (~(Qspnv6 & Xspnv6));
assign Xspnv6 = (~(Icyet6 & Djonv6));
assign Qspnv6 = (Etpnv6 & Ltpnv6);
assign Ltpnv6 = (~(Pwonv6 & Cmm7z6[1]));
assign Etpnv6 = (~(Rxonv6 & Stpnv6));
assign Chn7z6[19] = (~(Ztpnv6 & Gupnv6));
assign Gupnv6 = (Nupnv6 & Uupnv6);
assign Uupnv6 = (~(Pwonv6 & Cmm7z6[19]));
assign Nupnv6 = (~(Wwonv6 & HADDRI[19]));
assign Ztpnv6 = (Bvpnv6 & Ivpnv6);
assign Ivpnv6 = (~(Fvb7z6[19] & Rxonv6));
assign Bvpnv6 = (~(Hjn7z6[19] & Djonv6));
assign Chn7z6[18] = (~(Pvpnv6 & Wvpnv6));
assign Wvpnv6 = (Dwpnv6 & Kwpnv6);
assign Kwpnv6 = (~(Pwonv6 & Cmm7z6[18]));
assign Dwpnv6 = (~(Wwonv6 & HADDRI[18]));
assign Pvpnv6 = (Rwpnv6 & Ywpnv6);
assign Ywpnv6 = (~(Fvb7z6[18] & Rxonv6));
assign Rwpnv6 = (~(Hjn7z6[18] & Djonv6));
assign Chn7z6[17] = (~(Fxpnv6 & Mxpnv6));
assign Mxpnv6 = (Txpnv6 & Aypnv6);
assign Aypnv6 = (~(Pwonv6 & Cmm7z6[17]));
assign Txpnv6 = (~(Wwonv6 & HADDRI[17]));
assign Fxpnv6 = (Hypnv6 & Oypnv6);
assign Oypnv6 = (~(Fvb7z6[17] & Rxonv6));
assign Hypnv6 = (~(Hjn7z6[17] & Djonv6));
assign Chn7z6[16] = (~(Vypnv6 & Czpnv6));
assign Czpnv6 = (Jzpnv6 & Qzpnv6);
assign Qzpnv6 = (~(Pwonv6 & Cmm7z6[16]));
assign Jzpnv6 = (~(Wwonv6 & HADDRI[16]));
assign Vypnv6 = (Xzpnv6 & E0qnv6);
assign E0qnv6 = (~(Fvb7z6[16] & Rxonv6));
assign Xzpnv6 = (~(Hjn7z6[16] & Djonv6));
assign Chn7z6[15] = (~(L0qnv6 & S0qnv6));
assign S0qnv6 = (Z0qnv6 & G1qnv6);
assign G1qnv6 = (~(Pwonv6 & Cmm7z6[15]));
assign Z0qnv6 = (~(Wwonv6 & HADDRI[15]));
assign L0qnv6 = (N1qnv6 & U1qnv6);
assign U1qnv6 = (~(Fvb7z6[15] & Rxonv6));
assign N1qnv6 = (~(Hjn7z6[15] & Djonv6));
assign Chn7z6[14] = (~(B2qnv6 & I2qnv6));
assign I2qnv6 = (P2qnv6 & W2qnv6);
assign W2qnv6 = (~(Pwonv6 & Cmm7z6[14]));
assign P2qnv6 = (~(Wwonv6 & HADDRI[14]));
assign B2qnv6 = (D3qnv6 & K3qnv6);
assign K3qnv6 = (~(Fvb7z6[14] & Rxonv6));
assign D3qnv6 = (~(Hjn7z6[14] & Djonv6));
assign Chn7z6[13] = (~(R3qnv6 & Y3qnv6));
assign Y3qnv6 = (F4qnv6 & M4qnv6);
assign M4qnv6 = (~(Pwonv6 & Cmm7z6[13]));
assign F4qnv6 = (~(Wwonv6 & HADDRI[13]));
assign R3qnv6 = (T4qnv6 & A5qnv6);
assign A5qnv6 = (~(Fvb7z6[13] & Rxonv6));
assign T4qnv6 = (~(Hjn7z6[13] & Djonv6));
assign Chn7z6[12] = (~(H5qnv6 & O5qnv6));
assign O5qnv6 = (V5qnv6 & C6qnv6);
assign C6qnv6 = (~(Pwonv6 & Cmm7z6[12]));
assign V5qnv6 = (~(Wwonv6 & HADDRI[12]));
assign H5qnv6 = (J6qnv6 & Q6qnv6);
assign Q6qnv6 = (~(Fvb7z6[12] & Rxonv6));
assign J6qnv6 = (~(Hjn7z6[12] & Djonv6));
assign Chn7z6[11] = (~(X6qnv6 & E7qnv6));
assign E7qnv6 = (L7qnv6 & S7qnv6);
assign S7qnv6 = (~(Pwonv6 & Cmm7z6[11]));
assign L7qnv6 = (~(Wwonv6 & HADDRI[11]));
assign X6qnv6 = (Z7qnv6 & G8qnv6);
assign G8qnv6 = (~(Fvb7z6[11] & Rxonv6));
assign Z7qnv6 = (~(Hjn7z6[11] & Djonv6));
assign Chn7z6[10] = (~(N8qnv6 & U8qnv6));
assign U8qnv6 = (B9qnv6 & I9qnv6);
assign I9qnv6 = (~(Pwonv6 & Cmm7z6[10]));
assign B9qnv6 = (~(Wwonv6 & HADDRI[10]));
assign N8qnv6 = (P9qnv6 & W9qnv6);
assign W9qnv6 = (~(Fvb7z6[10] & Rxonv6));
assign P9qnv6 = (~(Hjn7z6[10] & Djonv6));
assign Chn7z6[0] = (~(Daqnv6 & Kaqnv6));
assign Kaqnv6 = (~(X9yet6 & Djonv6));
assign Daqnv6 = (Raqnv6 & Yaqnv6);
assign Yaqnv6 = (~(Pwonv6 & Cmm7z6[0]));
assign Pwonv6 = (Fbqnv6 & Yjonv6);
assign Raqnv6 = (~(Rxonv6 & Mbqnv6));
assign Gqpet6 = (Tbqnv6 ? W2n7z6[1] : J0n7z6[1]);
assign Hspet6 = (Tbqnv6 ? W2n7z6[0] : J0n7z6[0]);
assign Iupet6 = (Tbqnv6 ? J5n7z6[3] : Aym7z6[3]);
assign Jwpet6 = (Tbqnv6 ? J5n7z6[2] : Aym7z6[2]);
assign Kypet6 = (Tbqnv6 ? J5n7z6[1] : Aym7z6[1]);
assign L0qet6 = (Styet6 | J5n7z6[0]);
assign M2qet6 = (~(Acqnv6 & Hcqnv6));
assign Hcqnv6 = (~(W2n7z6[1] & Ocqnv6));
assign Acqnv6 = (Vcqnv6 & Cdqnv6);
assign Cdqnv6 = (~(Jdqnv6 & Qdqnv6));
assign Vcqnv6 = (~(Xdqnv6 & J0n7z6[1]));
assign N4qet6 = (~(Eeqnv6 & Leqnv6));
assign Leqnv6 = (~(W2n7z6[0] & Ocqnv6));
assign Eeqnv6 = (Seqnv6 & Zeqnv6);
assign Zeqnv6 = (~(Jdqnv6 & Gfqnv6));
assign Seqnv6 = (~(Xdqnv6 & J0n7z6[0]));
assign O6qet6 = (~(Nfqnv6 & Ufqnv6));
assign Ufqnv6 = (~(J5n7z6[3] & Ocqnv6));
assign Nfqnv6 = (Bgqnv6 & Igqnv6);
assign Igqnv6 = (~(Jdqnv6 & Pgqnv6));
assign Bgqnv6 = (~(Xdqnv6 & Aym7z6[3]));
assign P8qet6 = (~(Wgqnv6 & Dhqnv6));
assign Dhqnv6 = (~(J5n7z6[2] & Ocqnv6));
assign Wgqnv6 = (Khqnv6 & Rhqnv6);
assign Rhqnv6 = (~(Jdqnv6 & Yhqnv6));
assign Khqnv6 = (~(Xdqnv6 & Aym7z6[2]));
assign Qaqet6 = (~(Fiqnv6 & Miqnv6));
assign Miqnv6 = (~(J5n7z6[1] & Ocqnv6));
assign Fiqnv6 = (Tiqnv6 & Ajqnv6);
assign Ajqnv6 = (~(Jdqnv6 & Hjqnv6));
assign Tiqnv6 = (~(Xdqnv6 & Aym7z6[1]));
assign Rcqet6 = (Ojqnv6 | Jdqnv6);
assign Jdqnv6 = (~(Ocqnv6 | Vjqnv6));
assign Ojqnv6 = (Xdqnv6 | J5n7z6[0]);
assign Xdqnv6 = (~(Ocqnv6 | Gmnet6));
assign Ocqnv6 = (~(Ckqnv6 & Styet6));
assign Ckqnv6 = (~(Jkqnv6 | Kjonv6));
assign H8bdt6 = (Qkqnv6 & Ox9dt6);
assign Qkqnv6 = (~(Xkqnv6 & Elqnv6));
assign Elqnv6 = (~(G7bdt6 & Ez9dt6));
assign Us77v6 = (Drymz6[0] | Drymz6[1]);
assign Drymz6[1] = (~(Llqnv6 & Slqnv6));
assign Slqnv6 = (Zlqnv6 & Gmqnv6);
assign Gmqnv6 = (~(Nmqnv6 & Umqnv6));
assign Nmqnv6 = (W177v6 & Bnqnv6);
assign Zlqnv6 = (~(Inqnv6 & Pnqnv6));
assign Pnqnv6 = (Wnqnv6 | Doqnv6);
assign Llqnv6 = (Koqnv6 & Roqnv6);
assign Roqnv6 = (~(Yoqnv6 & Fpqnv6));
assign Drymz6[0] = (~(Mpqnv6 & Tpqnv6));
assign Tpqnv6 = (Aqqnv6 & Hqqnv6);
assign Hqqnv6 = (~(Oqqnv6 & Vqqnv6));
assign Vqqnv6 = (Crqnv6 & Jrqnv6);
assign Crqnv6 = (Bnqnv6 & Fpqnv6);
assign Oqqnv6 = (~(Qrqnv6 | Xrqnv6));
assign Xrqnv6 = (Unymz6[8] ? Lsqnv6 : Esqnv6);
assign Lsqnv6 = (Ssqnv6 & Zsqnv6);
assign Ssqnv6 = (~(Unymz6[10] & Gtqnv6));
assign Gtqnv6 = (Ntqnv6 | Utqnv6);
assign Ntqnv6 = (!Unymz6[9]);
assign Esqnv6 = (Unymz6[10] ? Iuqnv6 : Buqnv6);
assign Iuqnv6 = (Utqnv6 & Zsqnv6);
assign Zsqnv6 = (!Buqnv6);
assign Qrqnv6 = (~(Puqnv6 & Fy67v6));
assign Puqnv6 = (Unymz6[10] ? Dvqnv6 : Wuqnv6);
assign Dvqnv6 = (Kvqnv6 | Unymz6[9]);
assign Kvqnv6 = (Unymz6[8] ? Rvqnv6 : Utqnv6);
assign Rvqnv6 = (~(Buqnv6 & Utqnv6));
assign Buqnv6 = (Yvqnv6 & Fwqnv6);
assign Fwqnv6 = (Unymz6[1] ? Twqnv6 : Mwqnv6);
assign Twqnv6 = (~(Axqnv6 & Hxqnv6));
assign Hxqnv6 = (~(Unymz6[0] | Unymz6[3]));
assign Axqnv6 = (Lfp7z6[2] & Unymz6[2]);
assign Mwqnv6 = (~(Oxqnv6 & Vxqnv6));
assign Oxqnv6 = (Unymz6[3] ? Jyqnv6 : Cyqnv6);
assign Jyqnv6 = (Uh77v6 & Qyqnv6);
assign Cyqnv6 = (Lfp7z6[0] & Unymz6[2]);
assign Yvqnv6 = (Xyqnv6 & Ezqnv6);
assign Ezqnv6 = (~(Tn77v6 & Lzqnv6));
assign Xyqnv6 = (~(Unymz6[2] & Szqnv6));
assign Szqnv6 = (Zzqnv6 | Lzqnv6);
assign Zzqnv6 = (~(G0rnv6 | Vxqnv6));
assign Vxqnv6 = (!Unymz6[0]);
assign G0rnv6 = (Unymz6[1] ? U0rnv6 : N0rnv6);
assign N0rnv6 = (B1rnv6 | Unymz6[3]);
assign Wuqnv6 = (~(Utqnv6 & Unymz6[9]));
assign Utqnv6 = (I1rnv6 & P1rnv6);
assign P1rnv6 = (Unymz6[4] ? D2rnv6 : W1rnv6);
assign D2rnv6 = (~(Unymz6[6] & K2rnv6));
assign K2rnv6 = (Unymz6[5] ? Y2rnv6 : R2rnv6);
assign Y2rnv6 = (Unymz6[7] | Lfp7z6[3]);
assign R2rnv6 = (~(B1rnv6 | Unymz6[7]));
assign W1rnv6 = (~(F3rnv6 & M3rnv6));
assign F3rnv6 = (Unymz6[7] ? A4rnv6 : T3rnv6);
assign A4rnv6 = (Uh77v6 & H4rnv6);
assign H4rnv6 = (!Unymz6[6]);
assign T3rnv6 = (Lfp7z6[0] & Unymz6[6]);
assign I1rnv6 = (Unymz6[4] ? V4rnv6 : O4rnv6);
assign V4rnv6 = (~(Tn77v6 & C5rnv6));
assign O4rnv6 = (~(J5rnv6 & Q5rnv6));
assign Q5rnv6 = (~(M3rnv6 | Unymz6[7]));
assign M3rnv6 = (!Unymz6[5]);
assign J5rnv6 = (Lfp7z6[2] & Unymz6[6]);
assign Aqqnv6 = (~(Umqnv6 & Doqnv6));
assign Umqnv6 = (Inqnv6 & Ipymz6[1]);
assign Inqnv6 = (X5rnv6 & E6rnv6);
assign Mpqnv6 = (Koqnv6 & L6rnv6);
assign L6rnv6 = (~(Yoqnv6 & Wnqnv6));
assign Yoqnv6 = (S6rnv6 & Z6rnv6);
assign S6rnv6 = (P52nv6 & E6rnv6);
assign Koqnv6 = (G7rnv6 & N7rnv6);
assign N7rnv6 = (~(U7rnv6 & E6rnv6));
assign U7rnv6 = (~(B8rnv6 & I8rnv6));
assign I8rnv6 = (~(Wnqnv6 & P8rnv6));
assign P8rnv6 = (~(W177v6 & Ldo7v6));
assign B8rnv6 = (~(Ipymz6[1] & W8rnv6));
assign W8rnv6 = (~(D9rnv6 & K9rnv6));
assign K9rnv6 = (~(Doqnv6 & P52nv6));
assign Doqnv6 = (Ipymz6[0] & R9rnv6);
assign R9rnv6 = (Y9rnv6 | Uw77v6);
assign D9rnv6 = (~(F02nv6 & Bnqnv6));
assign G7rnv6 = (~(Farnv6 & Marnv6));
assign Marnv6 = (P52nv6 & Bnqnv6);
assign Farnv6 = (Z6rnv6 & Tarnv6);
assign Tarnv6 = (~(X477v6 & Ipymz6[1]));
assign Z6rnv6 = (!X5rnv6);
assign Ru77v6 = (~(Abrnv6 & Hbrnv6));
assign Hbrnv6 = (X5rnv6 | Jrqnv6);
assign Abrnv6 = (~(Uw77v6 & Y9rnv6));
assign Br77v6 = (Obrnv6 & Vbrnv6);
assign Vbrnv6 = (E6rnv6 & Jrqnv6);
assign Obrnv6 = (Ldo7v6 & Ccrnv6);
assign Ccrnv6 = (~(Jcrnv6 & Qcrnv6));
assign Qcrnv6 = (~(Wnqnv6 & W177v6));
assign Jcrnv6 = (~(Ipymz6[1] & Bnqnv6));
assign Bnqnv6 = (!Ipymz6[0]);
assign Ty77v6 = (~(Xcrnv6 & Edrnv6));
assign Edrnv6 = (~(Tn77v6 & Ldrnv6));
assign Ldrnv6 = (~(Sdrnv6 & Zdrnv6));
assign Zdrnv6 = (~(Bj77v6 & Gernv6));
assign Sdrnv6 = (Jrqnv6 ? Uernv6 : Nernv6);
assign Uernv6 = (~(Bfrnv6 & Ifrnv6));
assign Ifrnv6 = (Pfrnv6 & Wfrnv6);
assign Wfrnv6 = (~(Lfp7z6[1] & Blymz6[1]));
assign Pfrnv6 = (Dgrnv6 & Y9rnv6);
assign Dgrnv6 = (~(Lfp7z6[0] & Blymz6[0]));
assign Bfrnv6 = (Kgrnv6 & Rgrnv6);
assign Rgrnv6 = (~(Lfp7z6[2] & Blymz6[2]));
assign Kgrnv6 = (~(Lfp7z6[3] & Blymz6[3]));
assign Xcrnv6 = (Nernv6 ? Fhrnv6 : Ygrnv6);
assign Ygrnv6 = (~(Mhrnv6 & Jrqnv6));
assign Mhrnv6 = (~(Thrnv6 & Airnv6));
assign Airnv6 = (Hirnv6 & Oirnv6);
assign Oirnv6 = (~(Lfp7z6[0] & Kmymz6[0]));
assign Hirnv6 = (~(Lfp7z6[1] & Kmymz6[1]));
assign Thrnv6 = (Virnv6 & Cjrnv6);
assign Cjrnv6 = (~(Lfp7z6[2] & Kmymz6[2]));
assign Virnv6 = (~(Lfp7z6[3] & Kmymz6[3]));
assign Frc7v6 = (~(Jjrnv6 | Qjrnv6));
assign Phd7v6 = (Xjrnv6 & Vv67v6);
assign Xjrnv6 = (Ekrnv6 & Jrqnv6);
assign Ekrnv6 = (~(Lkrnv6 & Skrnv6));
assign Skrnv6 = (~(Zkrnv6 & Glrnv6));
assign Glrnv6 = (~(Hcymz6[4] ^ Nlrnv6));
assign Lkrnv6 = (~(Ulrnv6 & Bmrnv6));
assign Bmrnv6 = (~(Imrnv6 & Pmrnv6));
assign Pmrnv6 = (~(Nlrnv6 & Wmrnv6));
assign Wmrnv6 = (Dnrnv6 | Hcymz6[3]);
assign Ulrnv6 = (Knrnv6 & Rnrnv6);
assign Rnrnv6 = (~(Ynrnv6 & Fornv6));
assign Fornv6 = (Mornv6 | Tornv6);
assign Mornv6 = (Aprnv6 & Hprnv6);
assign Hprnv6 = (~(Hcymz6[1] & Oprnv6));
assign Oprnv6 = (~(Vprnv6 & Cqrnv6));
assign Cqrnv6 = (~(Fjd7v6 & Jqrnv6));
assign Jqrnv6 = (~(Qqrnv6 & Xqrnv6));
assign Xqrnv6 = (!Hcymz6[2]);
assign Vprnv6 = (~(Hcymz6[2] & Errnv6));
assign Aprnv6 = (Lrrnv6 & Dnrnv6);
assign Lrrnv6 = (~(Srrnv6 & Zrrnv6));
assign Srrnv6 = (~(Gsrnv6 | Fjd7v6));
assign Ynrnv6 = (Nsrnv6 & Usrnv6);
assign Usrnv6 = (~(Zrrnv6 & Btrnv6));
assign Btrnv6 = (~(Dnrnv6 & Itrnv6));
assign Itrnv6 = (~(Hcymz6[2] & Ptrnv6));
assign Ptrnv6 = (~(Wtrnv6 & Tornv6));
assign Tornv6 = (Durnv6 & Kurnv6);
assign Kurnv6 = (~(Errnv6 & Rurnv6));
assign Wtrnv6 = (~(Hcymz6[1] | Fjd7v6));
assign Nsrnv6 = (~(Yurnv6 & Fvrnv6));
assign Yurnv6 = (Dnrnv6 ^ Hcymz6[3]);
assign Knrnv6 = (~(Mvrnv6 & Tvrnv6));
assign Mvrnv6 = (Nlrnv6 ^ Hcymz6[4]);
assign Nlrnv6 = (~(Hcymz6[3] & Dnrnv6));
assign Dnrnv6 = (~(Awrnv6 & Rurnv6));
assign Rurnv6 = (!Hcymz6[1]);
assign Awrnv6 = (~(Hcymz6[2] | Fjd7v6));
assign G0d7v6 = (~(Hwrnv6 ^ Owrnv6));
assign Hwrnv6 = (~(Rr0nz6[0] & Vwrnv6));
assign M1d7v6 = (Cxrnv6 ^ Vwrnv6);
assign Vwrnv6 = (Jxrnv6 | E5d7v6);
assign S2d7v6 = (~(Qxrnv6 & Xxrnv6));
assign Qxrnv6 = (Lyrnv6 ? Eyrnv6 : Hw0nz6[2]);
assign G287v6 = (Syrnv6 & Zyrnv6);
assign Zyrnv6 = (Gzrnv6 & Nzrnv6);
assign Nzrnv6 = (E6rnv6 & Uzrnv6);
assign Gzrnv6 = (B0snv6 & I0snv6);
assign Syrnv6 = (P0snv6 & Xz67v6);
assign P0snv6 = (W0snv6 & D1snv6);
assign W0snv6 = (~(K1snv6 & R1snv6));
assign W387v6 = (Xz67v6 & Y1snv6);
assign Y1snv6 = (~(F2snv6 & M2snv6));
assign M2snv6 = (~(T2snv6 & I0snv6));
assign T2snv6 = (~(A3snv6 & H3snv6));
assign H3snv6 = (O3snv6 & V3snv6);
assign V3snv6 = (~(L587v6 | Tf87v6));
assign O3snv6 = (C4snv6 & J4snv6);
assign C4snv6 = (~(Q4snv6 & Qmbet6));
assign Q4snv6 = (~(X4snv6 | Wfo7v6));
assign A3snv6 = (E5snv6 & L5snv6);
assign L5snv6 = (Sgymz6[8] ? Z5snv6 : S5snv6);
assign Z5snv6 = (~(G6snv6 & N6snv6));
assign N6snv6 = (~(U6snv6 & B7snv6));
assign B7snv6 = (Sgymz6[10] | Sgymz6[9]);
assign S5snv6 = (I7snv6 | G6snv6);
assign I7snv6 = (Sgymz6[9] ? U6snv6 : Sgymz6[10]);
assign E5snv6 = (P7snv6 & W7snv6);
assign W7snv6 = (~(D8snv6 & Sgymz6[10]));
assign D8snv6 = (G6snv6 ? R8snv6 : K8snv6);
assign G6snv6 = (Y8snv6 & F9snv6);
assign F9snv6 = (Sgymz6[0] ? T9snv6 : M9snv6);
assign T9snv6 = (~(Aasnv6 & Hasnv6));
assign Hasnv6 = (~(Sgymz6[1] | Sgymz6[3]));
assign Aasnv6 = (Sgymz6[2] & Oasnv6);
assign M9snv6 = (~(Vasnv6 & Cbsnv6));
assign Vasnv6 = (Sgymz6[3] ? Qbsnv6 : Jbsnv6);
assign Qbsnv6 = (Uh77v6 & Xbsnv6);
assign Jbsnv6 = (Sgymz6[2] & Ecsnv6);
assign Y8snv6 = (Lcsnv6 & Scsnv6);
assign Scsnv6 = (~(Tn77v6 & Zcsnv6));
assign Lcsnv6 = (~(Sgymz6[2] & Gdsnv6));
assign Gdsnv6 = (Ndsnv6 | Zcsnv6);
assign Ndsnv6 = (~(Udsnv6 | Cbsnv6));
assign Cbsnv6 = (!Sgymz6[1]);
assign Udsnv6 = (Sgymz6[0] ? Iesnv6 : Besnv6);
assign Besnv6 = (Sgymz6[3] | Pesnv6);
assign R8snv6 = (~(Wesnv6 & Dfsnv6));
assign Wesnv6 = (~(U6snv6 & Kfsnv6));
assign K8snv6 = (Sgymz6[8] & Rfsnv6);
assign Rfsnv6 = (Dfsnv6 | U6snv6);
assign U6snv6 = (Yfsnv6 & Fgsnv6);
assign Fgsnv6 = (Sgymz6[4] ? Tgsnv6 : Mgsnv6);
assign Tgsnv6 = (Ahsnv6 | Hhsnv6);
assign Mgsnv6 = (Ohsnv6 & Vhsnv6);
assign Vhsnv6 = (~(Cisnv6 & Jisnv6));
assign Jisnv6 = (~(Sgymz6[5] | Sgymz6[6]));
assign Cisnv6 = (Uh77v6 & Sgymz6[7]);
assign Ohsnv6 = (Ahsnv6 | Qisnv6);
assign Ahsnv6 = (~(Xisnv6 & Sgymz6[6]));
assign Xisnv6 = (~(Sgymz6[5] | Sgymz6[7]));
assign Yfsnv6 = (Ejsnv6 & Ljsnv6);
assign Ljsnv6 = (~(Sjsnv6 & Zjsnv6));
assign Zjsnv6 = (Sgymz6[4] ? Nksnv6 : Gksnv6);
assign Nksnv6 = (Uksnv6 | Sgymz6[7]);
assign Gksnv6 = (~(Sgymz6[7] | Pesnv6));
assign Sjsnv6 = (Sgymz6[6] & Sgymz6[5]);
assign Ejsnv6 = (~(Tn77v6 & Blsnv6));
assign Dfsnv6 = (!Sgymz6[9]);
assign W8zmz6[1] = (~(Ilsnv6 & Plsnv6));
assign Plsnv6 = (~(Wlsnv6 & Hbb7v6));
assign Wlsnv6 = (Dmsnv6 & Uzrnv6);
assign Dmsnv6 = (~(Fgzmz6[0] & X477v6));
assign Ilsnv6 = (~(Kmsnv6 & Rmsnv6));
assign Rmsnv6 = (~(Ymsnv6 & Fnsnv6));
assign Xm87v6 = (~(Mnsnv6 & Tnsnv6));
assign Tnsnv6 = (~(Aosnv6 & Hosnv6));
assign Hosnv6 = (~(Wha7z6 | U7a7v6));
assign Aosnv6 = (N6c7v6 & Oosnv6);
assign Mnsnv6 = (~(Vosnv6 & Cpsnv6));
assign Oga7v6 = (~(J4snv6 & Jpsnv6));
assign Jpsnv6 = (~(Fgzmz6[0] & Qpsnv6));
assign Qpsnv6 = (~(Xpsnv6 & Eqsnv6));
assign Eqsnv6 = (~(Xco7v6 | Cdb7v6));
assign Xpsnv6 = (Lqsnv6 & Sqsnv6);
assign T5b7v6 = (~(Wfo7v6 & Zqsnv6));
assign Zqsnv6 = (~(Grsnv6 & Gdc7v6));
assign Grsnv6 = (Pfo7v6 & Nrsnv6);
assign L5zmz6[6] = (Ursnv6 ? Slzmz6[6] : Rjzmz6[6]);
assign L5zmz6[5] = (Ursnv6 ? Slzmz6[5] : Rjzmz6[5]);
assign L5zmz6[4] = (Ursnv6 ? Slzmz6[4] : Rjzmz6[4]);
assign L5zmz6[3] = (Ursnv6 ? Slzmz6[3] : Rjzmz6[3]);
assign L5zmz6[2] = (Ursnv6 ? Slzmz6[2] : Rjzmz6[2]);
assign L5zmz6[1] = (Ursnv6 ? Slzmz6[1] : Rjzmz6[1]);
assign Vzymz6[3] = (~(Bssnv6 & Issnv6));
assign Issnv6 = (~(Pssnv6 & Lczmz6[3]));
assign Bssnv6 = (Wssnv6 & Dtsnv6);
assign Dtsnv6 = (~(Ktsnv6 & Lczmz6[2]));
assign Wssnv6 = (Rtsnv6 | Ytsnv6);
assign Vzymz6[2] = (Rtsnv6 ^ Ytsnv6);
assign Ytsnv6 = (~(Ktsnv6 ^ Fusnv6));
assign Fusnv6 = (Pssnv6 & Lczmz6[2]);
assign Ktsnv6 = (~(Musnv6 | Tusnv6));
assign Rtsnv6 = (Avsnv6 | Hvsnv6);
assign Avsnv6 = (Ovsnv6 | Vvsnv6);
assign Vzymz6[1] = (~(Cwsnv6 ^ Vvsnv6));
assign Vvsnv6 = (~(Jwsnv6 ^ Musnv6));
assign Jwsnv6 = (~(Pssnv6 & Lczmz6[1]));
assign Cwsnv6 = (~(Hvsnv6 | Ovsnv6));
assign Vzymz6[0] = (Hvsnv6 ^ Ovsnv6);
assign Ovsnv6 = (~(Qwsnv6 & W9c7v6));
assign Qwsnv6 = (W8zmz6[0] & Cpsnv6);
assign Hvsnv6 = (~(Musnv6 & Xwsnv6));
assign Xwsnv6 = (~(Exsnv6 & Lxsnv6));
assign Lxsnv6 = (~(Lczmz6[0] & Pssnv6));
assign Musnv6 = (~(Sxsnv6 & Lczmz6[0]));
assign Sxsnv6 = (~(B0snv6 | Exsnv6));
assign Exsnv6 = (Wha7z6 ? Gysnv6 : Zxsnv6);
assign Gysnv6 = (Nysnv6 | H8c7v6);
assign Nysnv6 = (!W8zmz6[0]);
assign Zxsnv6 = (~(Uysnv6 & Oosnv6));
assign Uysnv6 = (~(U7a7v6 | N6c7v6));
assign U7a7v6 = (Bzsnv6 | K9a7v6);
assign K9a7v6 = (~(Izsnv6 & Pzsnv6));
assign Pzsnv6 = (~(Wzsnv6 & D0tnv6));
assign D0tnv6 = (K0tnv6 & R0tnv6);
assign K0tnv6 = (X4snv6 & Uzrnv6);
assign Wzsnv6 = (Y0tnv6 & Ztb7v6);
assign Y0tnv6 = (~(Xco7v6 | W577v6));
assign Bzsnv6 = (F1tnv6 & Jsb7v6);
assign F1tnv6 = (~(M1tnv6 | Wha7z6));
assign F787v6 = (~(T1tnv6 & A2tnv6));
assign A2tnv6 = (~(H2tnv6 | Oob7v6));
assign T1tnv6 = (Tvrnv6 & O2tnv6);
assign O2tnv6 = (~(Fgzmz6[0] & V2tnv6));
assign V2tnv6 = (~(C3tnv6 & J3tnv6));
assign J3tnv6 = (Q3tnv6 & X3tnv6);
assign Q3tnv6 = (~(S677v6 | Bba7v6));
assign C3tnv6 = (~(E4tnv6 | Edo7v6));
assign E4tnv6 = (W577v6 & L4tnv6);
assign L4tnv6 = (Nw97v6 | H8c7v6);
assign P0b7v6 = (~(S4tnv6 & Z4tnv6));
assign Z4tnv6 = (~(G5tnv6 & N5tnv6));
assign N5tnv6 = (U5tnv6 & B6tnv6);
assign B6tnv6 = (~(I6tnv6 | ETMINTNUM[6]));
assign I6tnv6 = (ETMINTNUM[7] | ETMINTNUM[8]);
assign U5tnv6 = (~(ETMINTNUM[4] | ETMINTNUM[5]));
assign G5tnv6 = (P6tnv6 & W6tnv6);
assign W6tnv6 = (~(D7tnv6 | ETMINTNUM[1]));
assign D7tnv6 = (ETMINTNUM[2] | ETMINTNUM[3]);
assign P6tnv6 = (~(ETMINTNUM[0] | K7tnv6));
assign S4tnv6 = (~(R7tnv6 & Y7tnv6));
assign Y7tnv6 = (Sqsnv6 & F8tnv6);
assign R7tnv6 = (D4b7v6 & Ldo7v6);
assign Qea7v6 = (~(Uzrnv6 & M8tnv6));
assign M8tnv6 = (~(T8tnv6 & Zt67v6));
assign Pma7v6 = (A9tnv6 & H9tnv6);
assign H9tnv6 = (Gsa7v6 & O9tnv6);
assign Ih87v6 = (Bhb7v6 & Fgzmz6[0]);
assign W3a7v6 = (~(V9tnv6 & Qjh7v6));
assign V9tnv6 = (W1a7v6 ? Rmb7v6 : Catnv6);
assign Catnv6 = (~(Soa7v6 & Mqa7v6));
assign P7b7v6 = (~(D1snv6 & Jatnv6));
assign Jatnv6 = (~(Qatnv6 & W8zmz6[0]));
assign D1snv6 = (!Oosnv6);
assign Vca7v6 = (!X3tnv6);
assign Yk87v6 = (Vosnv6 & W9c7v6);
assign Fj87v6 = (Xatnv6 & Ebtnv6);
assign Ebtnv6 = (Lbtnv6 & Sbtnv6);
assign Sbtnv6 = (~(Zbtnv6 & Gctnv6));
assign Gctnv6 = (~(Nctnv6 & Uctnv6));
assign Nctnv6 = (Bdtnv6 & Idtnv6);
assign Zbtnv6 = (!Pdtnv6);
assign Lbtnv6 = (Wdtnv6 & Detnv6);
assign Xatnv6 = (Ketnv6 & Vosnv6);
assign Vosnv6 = (Retnv6 & Wha7z6);
assign Retnv6 = (H8c7v6 & W8zmz6[0]);
assign Rwa7v6 = (~(Yetnv6 & Fftnv6));
assign Yetnv6 = (~(Mftnv6 & Tftnv6));
assign Gsa7v6 = (I9b7v6 | Agtnv6);
assign Zxymz6[4] = (~(Hgtnv6 & Ogtnv6));
assign Ogtnv6 = (~(Vgtnv6 & Chtnv6));
assign Chtnv6 = (~(Jhtnv6 & Qhtnv6));
assign Jhtnv6 = (Xhtnv6 & Eitnv6);
assign Xhtnv6 = (~(Litnv6 & Sitnv6));
assign Sitnv6 = (~(Zitnv6 & Gjtnv6));
assign Gjtnv6 = (Yhzmz6[0] | Yhzmz6[4]);
assign Litnv6 = (Njtnv6 & Ujtnv6);
assign Hgtnv6 = (Bktnv6 & Iktnv6);
assign Iktnv6 = (~(Pktnv6 & Wktnv6));
assign Pktnv6 = (Dltnv6 & Ujtnv6);
assign Bktnv6 = (~(Yhzmz6[4] & Kltnv6));
assign Kltnv6 = (Rltnv6 | Yhzmz6[3]);
assign Zxymz6[3] = (~(Yltnv6 & Fmtnv6));
assign Fmtnv6 = (Mmtnv6 & Tmtnv6);
assign Yltnv6 = (Antnv6 & Hntnv6);
assign Hntnv6 = (~(Dltnv6 & Ontnv6));
assign Ontnv6 = (Vntnv6 | Cotnv6);
assign Cotnv6 = (~(Njtnv6 | Jotnv6));
assign Vntnv6 = (Yhzmz6[2] ? Wktnv6 : Qotnv6);
assign Qotnv6 = (Yhzmz6[4] & Njtnv6);
assign Antnv6 = (Xotnv6 | Eptnv6);
assign Zxymz6[2] = (~(Lptnv6 & Sptnv6));
assign Sptnv6 = (Mmtnv6 & Eitnv6);
assign Eitnv6 = (Ujtnv6 | Zptnv6);
assign Mmtnv6 = (~(Gqtnv6 & Nqtnv6));
assign Nqtnv6 = (Uqtnv6 & Vgtnv6);
assign Uqtnv6 = (Brtnv6 & Njtnv6);
assign Gqtnv6 = (~(Ujtnv6 | Jotnv6));
assign Lptnv6 = (Irtnv6 & Prtnv6);
assign Prtnv6 = (~(Vgtnv6 & Wrtnv6));
assign Wrtnv6 = (~(Dstnv6 & Kstnv6));
assign Kstnv6 = (~(Rstnv6 & Yhzmz6[0]));
assign Rstnv6 = (Wktnv6 & Njtnv6);
assign Irtnv6 = (~(Yhzmz6[2] & Ystnv6));
assign Zxymz6[1] = (~(Fttnv6 & Mttnv6));
assign Mttnv6 = (Tttnv6 & Zptnv6);
assign Zptnv6 = (~(Autnv6 & Yhzmz6[1]));
assign Fttnv6 = (Hutnv6 & Outnv6);
assign Outnv6 = (~(Yhzmz6[1] & Ystnv6));
assign Ystnv6 = (~(Eptnv6 & Zitnv6));
assign Hutnv6 = (Rltnv6 | Vutnv6);
assign Zxymz6[0] = (~(Cvtnv6 & Jvtnv6));
assign Jvtnv6 = (Qvtnv6 & Tmtnv6);
assign Tmtnv6 = (~(Xvtnv6 & Yhzmz6[1]));
assign Xvtnv6 = (Yhzmz6[0] & Wktnv6);
assign Wktnv6 = (!Zitnv6);
assign Qvtnv6 = (Ewtnv6 | Jotnv6);
assign Ewtnv6 = (~(Dltnv6 & Tttnv6));
assign Tttnv6 = (!Lwtnv6);
assign Dltnv6 = (~(Rltnv6 | Yhzmz6[0]));
assign Cvtnv6 = (Qhtnv6 & Swtnv6);
assign Swtnv6 = (Brtnv6 | Eptnv6);
assign Eptnv6 = (~(Rltnv6 | Yhzmz6[4]));
assign Rltnv6 = (!Vgtnv6);
assign Vgtnv6 = (Zwtnv6 & Gxtnv6);
assign Gxtnv6 = (~(Zxymz6[7] | Zxymz6[8]));
assign Zwtnv6 = (~(Zxymz6[5] | Zxymz6[6]));
assign Qhtnv6 = (Vutnv6 & Dstnv6);
assign Dstnv6 = (Nxtnv6 | Jotnv6);
assign Vutnv6 = (Uxtnv6 & Bytnv6);
assign Bytnv6 = (Nxtnv6 | Zitnv6);
assign Zitnv6 = (Xotnv6 | Yhzmz6[4]);
assign Xotnv6 = (!Yhzmz6[3]);
assign Nxtnv6 = (~(Iytnv6 & Yhzmz6[2]));
assign Iytnv6 = (Yhzmz6[0] & Njtnv6);
assign Njtnv6 = (!Yhzmz6[1]);
assign Uxtnv6 = (~(Autnv6 & Lwtnv6));
assign Lwtnv6 = (Yhzmz6[1] & Ujtnv6);
assign Ujtnv6 = (!Yhzmz6[2]);
assign Autnv6 = (~(Brtnv6 | Jotnv6));
assign Jotnv6 = (Yhzmz6[3] | Yhzmz6[4]);
assign Brtnv6 = (!Yhzmz6[0]);
assign Rka7v6 = (~(Pytnv6 & Nrsnv6));
assign Pytnv6 = (Jjh7v6 & Wytnv6);
assign Wytnv6 = (!Mbc7v6);
assign I7zmz6[9] = (~(Dztnv6 & Kztnv6));
assign Kztnv6 = (~(Ot77z6 & Rztnv6));
assign Dztnv6 = (Yztnv6 & F0unv6);
assign F0unv6 = (~(Kk97v6 & M0unv6));
assign Yztnv6 = (~(T0unv6 & Rjzmz6[9]));
assign I7zmz6[8] = (~(A1unv6 & H1unv6));
assign H1unv6 = (~(Wt77z6 & Rztnv6));
assign A1unv6 = (O1unv6 & V1unv6);
assign V1unv6 = (~(Tl97v6 & M0unv6));
assign O1unv6 = (~(T0unv6 & Rjzmz6[8]));
assign I7zmz6[7] = (~(C2unv6 & J2unv6));
assign J2unv6 = (~(Eu77z6 & Rztnv6));
assign C2unv6 = (Q2unv6 & X2unv6);
assign X2unv6 = (~(Cn97v6 & M0unv6));
assign Q2unv6 = (~(T0unv6 & Rjzmz6[7]));
assign I7zmz6[6] = (~(E3unv6 & L3unv6));
assign L3unv6 = (~(Mu77z6 & Rztnv6));
assign E3unv6 = (S3unv6 & Z3unv6);
assign Z3unv6 = (~(Lo97v6 & M0unv6));
assign S3unv6 = (~(T0unv6 & Rjzmz6[6]));
assign I7zmz6[5] = (~(G4unv6 & N4unv6));
assign N4unv6 = (~(Uu77z6 & Rztnv6));
assign G4unv6 = (U4unv6 & B5unv6);
assign B5unv6 = (~(Up97v6 & M0unv6));
assign U4unv6 = (~(T0unv6 & Rjzmz6[5]));
assign I7zmz6[4] = (~(I5unv6 & P5unv6));
assign P5unv6 = (~(Cv77z6 & Rztnv6));
assign I5unv6 = (W5unv6 & D6unv6);
assign D6unv6 = (~(Dr97v6 & M0unv6));
assign W5unv6 = (~(T0unv6 & Rjzmz6[4]));
assign I7zmz6[3] = (~(K6unv6 & R6unv6));
assign R6unv6 = (~(Kv77z6 & Rztnv6));
assign K6unv6 = (Y6unv6 & F7unv6);
assign F7unv6 = (~(Ms97v6 & M0unv6));
assign Y6unv6 = (~(T0unv6 & Rjzmz6[3]));
assign I7zmz6[31] = (~(M7unv6 & T7unv6));
assign T7unv6 = (~(Um77z6 & Rztnv6));
assign M7unv6 = (A8unv6 & H8unv6);
assign H8unv6 = (~(Uq87v6 & M0unv6));
assign A8unv6 = (~(T0unv6 & Rjzmz6[31]));
assign I7zmz6[30] = (~(O8unv6 & V8unv6));
assign V8unv6 = (~(Cn77z6 & Rztnv6));
assign O8unv6 = (C9unv6 & J9unv6);
assign J9unv6 = (~(Ds87v6 & M0unv6));
assign C9unv6 = (~(T0unv6 & Rjzmz6[30]));
assign I7zmz6[2] = (~(Q9unv6 & X9unv6));
assign X9unv6 = (~(Sv77z6 & Rztnv6));
assign Q9unv6 = (Eaunv6 & Launv6);
assign Launv6 = (~(Vt97v6 & M0unv6));
assign Eaunv6 = (~(T0unv6 & Rjzmz6[2]));
assign I7zmz6[29] = (~(Saunv6 & Zaunv6));
assign Zaunv6 = (~(Kn77z6 & Rztnv6));
assign Saunv6 = (Gbunv6 & Nbunv6);
assign Nbunv6 = (~(Mt87v6 & M0unv6));
assign Gbunv6 = (~(T0unv6 & Rjzmz6[29]));
assign I7zmz6[28] = (~(Ubunv6 & Bcunv6));
assign Bcunv6 = (~(Sn77z6 & Rztnv6));
assign Ubunv6 = (Icunv6 & Pcunv6);
assign Pcunv6 = (~(Vu87v6 & M0unv6));
assign Icunv6 = (~(T0unv6 & Rjzmz6[28]));
assign I7zmz6[27] = (~(Wcunv6 & Ddunv6));
assign Ddunv6 = (~(Ao77z6 & Rztnv6));
assign Wcunv6 = (Kdunv6 & Rdunv6);
assign Rdunv6 = (~(Ew87v6 & M0unv6));
assign Kdunv6 = (~(T0unv6 & Rjzmz6[27]));
assign I7zmz6[26] = (~(Ydunv6 & Feunv6));
assign Feunv6 = (~(Io77z6 & Rztnv6));
assign Ydunv6 = (Meunv6 & Teunv6);
assign Teunv6 = (~(Nx87v6 & M0unv6));
assign Meunv6 = (~(T0unv6 & Rjzmz6[26]));
assign I7zmz6[25] = (~(Afunv6 & Hfunv6));
assign Hfunv6 = (~(Qo77z6 & Rztnv6));
assign Afunv6 = (Ofunv6 & Vfunv6);
assign Vfunv6 = (~(Wy87v6 & M0unv6));
assign Ofunv6 = (~(T0unv6 & Rjzmz6[25]));
assign I7zmz6[24] = (~(Cgunv6 & Jgunv6));
assign Jgunv6 = (~(Yo77z6 & Rztnv6));
assign Cgunv6 = (Qgunv6 & Xgunv6);
assign Xgunv6 = (~(F097v6 & M0unv6));
assign Qgunv6 = (~(T0unv6 & Rjzmz6[24]));
assign I7zmz6[23] = (~(Ehunv6 & Lhunv6));
assign Lhunv6 = (~(Gp77z6 & Rztnv6));
assign Ehunv6 = (Shunv6 & Zhunv6);
assign Zhunv6 = (~(O197v6 & M0unv6));
assign Shunv6 = (~(T0unv6 & Rjzmz6[23]));
assign I7zmz6[22] = (~(Giunv6 & Niunv6));
assign Niunv6 = (~(Op77z6 & Rztnv6));
assign Giunv6 = (Uiunv6 & Bjunv6);
assign Bjunv6 = (~(X297v6 & M0unv6));
assign Uiunv6 = (~(T0unv6 & Rjzmz6[22]));
assign I7zmz6[21] = (~(Ijunv6 & Pjunv6));
assign Pjunv6 = (~(Wp77z6 & Rztnv6));
assign Ijunv6 = (Wjunv6 & Dkunv6);
assign Dkunv6 = (~(G497v6 & M0unv6));
assign Wjunv6 = (~(T0unv6 & Rjzmz6[21]));
assign I7zmz6[20] = (~(Kkunv6 & Rkunv6));
assign Rkunv6 = (~(Eq77z6 & Rztnv6));
assign Kkunv6 = (Ykunv6 & Flunv6);
assign Flunv6 = (~(P597v6 & M0unv6));
assign Ykunv6 = (~(Rjzmz6[20] & T0unv6));
assign I7zmz6[1] = (~(Mlunv6 & Tlunv6));
assign Tlunv6 = (~(Aw77z6 & Rztnv6));
assign Mlunv6 = (Amunv6 & Hmunv6);
assign Hmunv6 = (~(Ev97v6 & M0unv6));
assign Amunv6 = (~(T0unv6 & Rjzmz6[1]));
assign I7zmz6[19] = (~(Omunv6 & Vmunv6));
assign Vmunv6 = (~(Mq77z6 & Rztnv6));
assign Omunv6 = (Cnunv6 & Jnunv6);
assign Jnunv6 = (~(Y697v6 & M0unv6));
assign Cnunv6 = (~(T0unv6 & Rjzmz6[19]));
assign I7zmz6[18] = (~(Qnunv6 & Xnunv6));
assign Xnunv6 = (~(Uq77z6 & Rztnv6));
assign Qnunv6 = (Eounv6 & Lounv6);
assign Lounv6 = (~(H897v6 & M0unv6));
assign Eounv6 = (~(T0unv6 & Rjzmz6[18]));
assign I7zmz6[17] = (~(Sounv6 & Zounv6));
assign Zounv6 = (~(Cr77z6 & Rztnv6));
assign Sounv6 = (Gpunv6 & Npunv6);
assign Npunv6 = (~(Q997v6 & M0unv6));
assign Gpunv6 = (~(T0unv6 & Rjzmz6[17]));
assign I7zmz6[16] = (~(Upunv6 & Bqunv6));
assign Bqunv6 = (~(Kr77z6 & Rztnv6));
assign Upunv6 = (Iqunv6 & Pqunv6);
assign Pqunv6 = (~(Za97v6 & M0unv6));
assign Iqunv6 = (~(T0unv6 & Rjzmz6[16]));
assign I7zmz6[15] = (~(Wqunv6 & Drunv6));
assign Drunv6 = (~(Sr77z6 & Rztnv6));
assign Wqunv6 = (Krunv6 & Rrunv6);
assign Rrunv6 = (~(Ic97v6 & M0unv6));
assign Krunv6 = (~(T0unv6 & Rjzmz6[15]));
assign I7zmz6[14] = (~(Yrunv6 & Fsunv6));
assign Fsunv6 = (~(As77z6 & Rztnv6));
assign Yrunv6 = (Msunv6 & Tsunv6);
assign Tsunv6 = (~(Rd97v6 & M0unv6));
assign Msunv6 = (~(T0unv6 & Rjzmz6[14]));
assign I7zmz6[13] = (~(Atunv6 & Htunv6));
assign Htunv6 = (~(Is77z6 & Rztnv6));
assign Atunv6 = (Otunv6 & Vtunv6);
assign Vtunv6 = (~(Af97v6 & M0unv6));
assign Otunv6 = (~(T0unv6 & Rjzmz6[13]));
assign I7zmz6[12] = (~(Cuunv6 & Juunv6));
assign Juunv6 = (~(Qs77z6 & Rztnv6));
assign Cuunv6 = (Quunv6 & Xuunv6);
assign Xuunv6 = (~(Jg97v6 & M0unv6));
assign Quunv6 = (~(T0unv6 & Rjzmz6[12]));
assign I7zmz6[11] = (~(Evunv6 & Lvunv6));
assign Lvunv6 = (~(Ys77z6 & Rztnv6));
assign Evunv6 = (Svunv6 & Zvunv6);
assign Zvunv6 = (~(Sh97v6 & M0unv6));
assign Svunv6 = (~(T0unv6 & Rjzmz6[11]));
assign I7zmz6[10] = (~(Gwunv6 & Nwunv6));
assign Nwunv6 = (~(Gt77z6 & Rztnv6));
assign Gwunv6 = (Uwunv6 & Bxunv6);
assign Bxunv6 = (~(Bj97v6 & M0unv6));
assign Uwunv6 = (~(T0unv6 & Rjzmz6[10]));
assign Lua7v6 = (Ixunv6 & Agtnv6);
assign Agtnv6 = (!K7tnv6);
assign Ixunv6 = (F02nv6 & R0tnv6);
assign Mqa7v6 = (!Pxunv6);
assign Nw97v6 = (~(Wxunv6 & Dyunv6));
assign Dyunv6 = (~(Kyunv6 & Detnv6));
assign Kyunv6 = (~(Ryunv6 & Yyunv6));
assign Yyunv6 = (~(M0unv6 & H8c7v6));
assign M0unv6 = (~(Rztnv6 | Fzunv6));
assign Ryunv6 = (~(T0unv6 & N6c7v6));
assign T0unv6 = (~(Mzunv6 | Rztnv6));
assign Rztnv6 = (Wdtnv6 | Xco7v6);
assign Mzunv6 = (!Fzunv6);
assign Wxunv6 = (~(Ketnv6 & Wdtnv6));
assign Cy97v6 = (Tzunv6 & Wdtnv6);
assign Tzunv6 = (T077v6 ? Qobet6 : A0vnv6);
assign T1zmz6[9] = (H0vnv6 ? L5zmz6[9] : L5zmz6[8]);
assign T1zmz6[8] = (H0vnv6 ? L5zmz6[8] : L5zmz6[7]);
assign T1zmz6[7] = (~(O0vnv6 & V0vnv6));
assign V0vnv6 = (~(C1vnv6 & J1vnv6));
assign J1vnv6 = (~(Q1vnv6 & X1vnv6));
assign X1vnv6 = (E2vnv6 & L2vnv6);
assign L2vnv6 = (S2vnv6 & Z2vnv6);
assign S2vnv6 = (~(P3zmz6[7] & G3vnv6));
assign E2vnv6 = (N3vnv6 & U3vnv6);
assign U3vnv6 = (~(L5zmz6[10] ^ P3zmz6[10]));
assign N3vnv6 = (~(L5zmz6[11] ^ P3zmz6[11]));
assign Q1vnv6 = (B4vnv6 & I4vnv6);
assign I4vnv6 = (~(L5zmz6[9] ^ P3zmz6[9]));
assign B4vnv6 = (P4vnv6 & W4vnv6);
assign W4vnv6 = (~(L5zmz6[12] ^ P3zmz6[12]));
assign P4vnv6 = (~(L5zmz6[8] ^ P3zmz6[8]));
assign O0vnv6 = (D5vnv6 & K5vnv6);
assign D5vnv6 = (~(L5zmz6[7] & R5vnv6));
assign R5vnv6 = (~(P3zmz6[7] & C1vnv6));
assign T1zmz6[35] = (C1vnv6 & L5zmz6[31]);
assign T1zmz6[34] = (C1vnv6 & L5zmz6[30]);
assign T1zmz6[33] = (~(Y5vnv6 & F6vnv6));
assign F6vnv6 = (~(Oosnv6 & M6vnv6));
assign M6vnv6 = (Y5a7v6 | Fgzmz6[1]);
assign Y5vnv6 = (~(C1vnv6 & L5zmz6[29]));
assign T1zmz6[32] = (~(T6vnv6 & A7vnv6));
assign A7vnv6 = (~(Oosnv6 & H7vnv6));
assign H7vnv6 = (Uzrnv6 | Y5a7v6);
assign Y5a7v6 = (I1c7v6 ? R0tnv6 : O7vnv6);
assign O7vnv6 = (Qvb7v6 & V7vnv6);
assign V7vnv6 = (~(Xw67v6 & C8vnv6));
assign C8vnv6 = (J2b7v6 | Hqb7v6);
assign T6vnv6 = (~(C1vnv6 & L5zmz6[28]));
assign T1zmz6[31] = (H0vnv6 ? L5zmz6[31] : J8vnv6);
assign T1zmz6[30] = (!Q8vnv6);
assign Q8vnv6 = (C1vnv6 ? E9vnv6 : X8vnv6);
assign E9vnv6 = (J8vnv6 ? L9vnv6 : Z2vnv6);
assign T1zmz6[29] = (H0vnv6 ? L5zmz6[29] : L5zmz6[26]);
assign T1zmz6[28] = (H0vnv6 ? L5zmz6[28] : L5zmz6[25]);
assign T1zmz6[27] = (H0vnv6 ? L5zmz6[27] : L5zmz6[24]);
assign T1zmz6[26] = (H0vnv6 ? L5zmz6[26] : L5zmz6[23]);
assign T1zmz6[25] = (H0vnv6 ? L5zmz6[25] : L5zmz6[22]);
assign T1zmz6[24] = (H0vnv6 ? L5zmz6[24] : L5zmz6[21]);
assign T1zmz6[23] = (H0vnv6 ? L5zmz6[23] : S9vnv6);
assign T1zmz6[22] = (H0vnv6 ? L5zmz6[22] : Z9vnv6);
assign Z9vnv6 = (S9vnv6 ? Tct8v6 : Zz97v6);
assign T1zmz6[21] = (H0vnv6 ? L5zmz6[21] : L5zmz6[19]);
assign T1zmz6[20] = (H0vnv6 ? Tct8v6 : L5zmz6[18]);
assign T1zmz6[19] = (H0vnv6 ? L5zmz6[19] : L5zmz6[17]);
assign T1zmz6[18] = (H0vnv6 ? L5zmz6[18] : L5zmz6[16]);
assign T1zmz6[17] = (H0vnv6 ? L5zmz6[17] : L5zmz6[15]);
assign T1zmz6[16] = (H0vnv6 ? L5zmz6[16] : L5zmz6[14]);
assign T1zmz6[15] = (~(K5vnv6 & Gavnv6));
assign Gavnv6 = (~(L5zmz6[15] & H0vnv6));
assign K5vnv6 = (!Navnv6);
assign T1zmz6[14] = (Uavnv6 | Bbvnv6);
assign Bbvnv6 = (Navnv6 & L5zmz6[13]);
assign Navnv6 = (~(H0vnv6 | Ibvnv6));
assign Uavnv6 = (C1vnv6 ? Pbvnv6 : L5zmz6[14]);
assign C1vnv6 = (!H0vnv6);
assign Pbvnv6 = (Ibvnv6 & Zz97v6);
assign Ibvnv6 = (Wbvnv6 & Dcvnv6);
assign Dcvnv6 = (Kcvnv6 & Rcvnv6);
assign Rcvnv6 = (Ycvnv6 & Fdvnv6);
assign Fdvnv6 = (!S9vnv6);
assign S9vnv6 = (~(Mdvnv6 & Tdvnv6));
assign Tdvnv6 = (Aevnv6 & Hevnv6);
assign Hevnv6 = (Oevnv6 & Vevnv6);
assign Vevnv6 = (!J8vnv6);
assign J8vnv6 = (~(Cfvnv6 & Jfvnv6));
assign Jfvnv6 = (Qfvnv6 & Xfvnv6);
assign Xfvnv6 = (~(L5zmz6[29] ^ P3zmz6[29]));
assign Qfvnv6 = (Egvnv6 & Lgvnv6);
assign Lgvnv6 = (~(L5zmz6[31] ^ P3zmz6[31]));
assign Egvnv6 = (X8vnv6 ^ P3zmz6[30]);
assign Cfvnv6 = (Sgvnv6 & Zgvnv6);
assign Zgvnv6 = (L9vnv6 ^ P3zmz6[27]);
assign Sgvnv6 = (~(L5zmz6[28] ^ P3zmz6[28]));
assign Oevnv6 = (~(P3zmz6[20] ^ Tct8v6));
assign Aevnv6 = (Ghvnv6 & Nhvnv6);
assign Nhvnv6 = (~(L5zmz6[21] ^ P3zmz6[21]));
assign Ghvnv6 = (~(L5zmz6[22] ^ P3zmz6[22]));
assign Mdvnv6 = (Uhvnv6 & Bivnv6);
assign Bivnv6 = (Iivnv6 & Pivnv6);
assign Pivnv6 = (~(L5zmz6[23] ^ P3zmz6[23]));
assign Iivnv6 = (~(L5zmz6[24] ^ P3zmz6[24]));
assign Uhvnv6 = (Wivnv6 & Djvnv6);
assign Djvnv6 = (~(L5zmz6[25] ^ P3zmz6[25]));
assign Wivnv6 = (~(L5zmz6[26] ^ P3zmz6[26]));
assign Ycvnv6 = (~(L5zmz6[13] ^ P3zmz6[13]));
assign Kcvnv6 = (Kjvnv6 & Rjvnv6);
assign Rjvnv6 = (~(L5zmz6[14] ^ P3zmz6[14]));
assign Kjvnv6 = (~(L5zmz6[15] ^ P3zmz6[15]));
assign Wbvnv6 = (Yjvnv6 & Fkvnv6);
assign Fkvnv6 = (Mkvnv6 & Tkvnv6);
assign Tkvnv6 = (~(L5zmz6[16] ^ P3zmz6[16]));
assign Mkvnv6 = (~(L5zmz6[17] ^ P3zmz6[17]));
assign Yjvnv6 = (Alvnv6 & Hlvnv6);
assign Hlvnv6 = (~(L5zmz6[18] ^ P3zmz6[18]));
assign Alvnv6 = (~(L5zmz6[19] ^ P3zmz6[19]));
assign T1zmz6[13] = (H0vnv6 ? L5zmz6[13] : L5zmz6[12]);
assign T1zmz6[12] = (H0vnv6 ? L5zmz6[12] : L5zmz6[11]);
assign T1zmz6[11] = (H0vnv6 ? L5zmz6[11] : L5zmz6[10]);
assign T1zmz6[10] = (H0vnv6 ? L5zmz6[10] : L5zmz6[9]);
assign Sa77v6 = (Ue77z6 & Jrqnv6);
assign T0adt6 = (~(Olvnv6 & Vlvnv6));
assign Vlvnv6 = (~(D1adt6 & Xkqnv6));
assign Is97z6 = (~(Cmvnv6 & Jmvnv6));
assign Jmvnv6 = (Qmvnv6 & Xmvnv6);
assign Cmvnv6 = (Envnv6 & Woinv6);
assign Woinv6 = (~(Lnvnv6 & Snvnv6));
assign Lnvnv6 = (Znvnv6 & Bfo7v6);
assign Ys97z6 = (~(Govnv6 & Envnv6));
assign Govnv6 = (Xmvnv6 & Ywinv6);
assign Ywinv6 = (!Qs97z6);
assign Qs97z6 = (~(Novnv6 & Uovnv6));
assign Uovnv6 = (Bpvnv6 & Ipvnv6);
assign Novnv6 = (~(Poinv6 | Ppvnv6));
assign Ppvnv6 = (!Wpvnv6);
assign Gt97z6 = (~(Dqvnv6 & Kpinv6));
assign Kpinv6 = (Kqvnv6 & Rqvnv6);
assign Rqvnv6 = (~(Yqvnv6 & Frvnv6));
assign Dqvnv6 = (Mrvnv6 & Trvnv6);
assign Mrvnv6 = (~(Poinv6 & Asvnv6));
assign Asvnv6 = (~(Hsvnv6 & Osvnv6));
assign Osvnv6 = (Vsvnv6 & Ctvnv6);
assign Ctvnv6 = (~(Jtvnv6 & Qtvnv6));
assign Jtvnv6 = (~(Xtvnv6 & Dwb7z6[2]));
assign Vsvnv6 = (~(Euvnv6 & Luvnv6));
assign Hsvnv6 = (Suvnv6 & Zuvnv6);
assign Zuvnv6 = (~(Dwb7z6[2] & Gvvnv6));
assign Suvnv6 = (Bwvnv6 ? Uvvnv6 : Nvvnv6);
assign Poinv6 = (Iwvnv6 & Bfo7v6);
assign Ot97z6 = (~(Pwvnv6 & Trvnv6));
assign Trvnv6 = (~(Wwvnv6 & Frvnv6));
assign Pwvnv6 = (Ipvnv6 & Dxvnv6);
assign Ipvnv6 = (~(Kxvnv6 & Frvnv6));
assign Frvnv6 = (~(Gaonv6 | Iga7z6));
assign C3a7z6 = (!SWCLKTCK);
assign Y4a7z6 = (~(Rxvnv6 & Kqvnv6));
assign Kqvnv6 = (Yxvnv6 & Envnv6);
assign Envnv6 = (Fyvnv6 & Myvnv6);
assign Myvnv6 = (~(Tyvnv6 & Azvnv6));
assign Azvnv6 = (Hzvnv6 & Ozvnv6);
assign Hzvnv6 = (Vzvnv6 & C0wnv6);
assign Tyvnv6 = (J0wnv6 & Q0wnv6);
assign J0wnv6 = (X0wnv6 & E1wnv6);
assign Fyvnv6 = (~(L1wnv6 & S1wnv6));
assign L1wnv6 = (Ldo7v6 & Qg2nv6);
assign Yxvnv6 = (Qmvnv6 & Bpvnv6);
assign Qmvnv6 = (~(Z1wnv6 & G2wnv6));
assign G2wnv6 = (Dxvnv6 & Iga7z6);
assign Z1wnv6 = (Fqinv6 & Bpvnv6);
assign Fqinv6 = (Wpvnv6 & Xmvnv6);
assign Rxvnv6 = (Wpvnv6 & Dxvnv6);
assign W5a7z6 = (!Bj2nv6);
assign Cfa7z6 = (V5jnv6 & N2wnv6);
assign N2wnv6 = (~(M4jnv6 & T4jnv6));
assign M4jnv6 = (!Vvlnv6);
assign Vvlnv6 = (H5jnv6 | U2wnv6);
assign H5jnv6 = (~(B3wnv6 & I3wnv6));
assign Qga7z6 = (!Olzdt6);
assign Yga7z6 = (!Rgo7v6);
assign Kja7z6 = (!Hsi7z6[1]);
assign Sja7z6 = (!Hsi7z6[0]);
assign Dwl8v6 = (P3wnv6 & Glh7v6);
assign P3wnv6 = (~(W3wnv6 | Zkh7v6));
assign Wvl8v6 = (D4wnv6 ^ Tmg7z6[32]);
assign Pvl8v6 = (Bt0ft6 & K4wnv6);
assign K4wnv6 = (!G5a7z6);
assign G5a7z6 = (~(R4wnv6 & Y4wnv6));
assign Y4wnv6 = (~(F5wnv6 & Ejo7z6[0]));
assign F5wnv6 = (M5wnv6 & Ejo7z6[1]);
assign R4wnv6 = (T5wnv6 | A6wnv6);
assign Bt0ft6 = (~(H6wnv6 & O6wnv6));
assign O6wnv6 = (~(V6wnv6 & C7wnv6));
assign H6wnv6 = (J7wnv6 & A6wnv6);
assign J7wnv6 = (~(M5wnv6 & Ejo7z6[1]));
assign M5wnv6 = (!Q7wnv6);
assign Ivl8v6 = (~(X7wnv6 & E8wnv6));
assign E8wnv6 = (~(L8wnv6 & Itb7z6[31]));
assign X7wnv6 = (S8wnv6 & Z8wnv6);
assign Z8wnv6 = (~(G9wnv6 & N9wnv6));
assign N9wnv6 = (~(U9wnv6 & Bawnv6));
assign Bawnv6 = (Iawnv6 & Pawnv6);
assign Pawnv6 = (Wawnv6 | Dbwnv6);
assign Iawnv6 = (~(Dtm7z6[3] & Kbwnv6));
assign U9wnv6 = (Rbwnv6 & Ybwnv6);
assign Ybwnv6 = (~(Dtm7z6[0] & HRDATAD[31]));
assign Rbwnv6 = (~(Dtm7z6[1] & HRDATAS[31]));
assign S8wnv6 = (~(Fcwnv6 & Mcwnv6));
assign Bvl8v6 = (Adwnv6 ? Tcwnv6 : Dbymz6[1]);
assign Tcwnv6 = (Dbymz6[0] & Hdwnv6);
assign Hdwnv6 = (~(Odwnv6 & Vdwnv6));
assign Vdwnv6 = (Dbymz6[1] & Cewnv6);
assign Odwnv6 = (Jewnv6 & Qewnv6);
assign Uul8v6 = (~(Xewnv6 & Efwnv6));
assign Efwnv6 = (Lfwnv6 & Sfwnv6);
assign Sfwnv6 = (~(Tfxmz6[11] & Zfwnv6));
assign Lfwnv6 = (~(Njxmz6[11] & Ggwnv6));
assign Xewnv6 = (Ngwnv6 & Ugwnv6);
assign Ugwnv6 = (~(Ub67v6 & Bhwnv6));
assign Ngwnv6 = (~(Hnxmz6[11] & Ihwnv6));
assign Nul8v6 = (~(Phwnv6 & Whwnv6));
assign Whwnv6 = (~(Diwnv6 & Tfxmz6[11]));
assign Phwnv6 = (Kiwnv6 & Riwnv6);
assign Riwnv6 = (~(Yiwnv6 & Hnxmz6[11]));
assign Kiwnv6 = (~(L5ymz6[26] & Fjwnv6));
assign Gul8v6 = (~(Mjwnv6 & Tjwnv6));
assign Tjwnv6 = (Akwnv6 & Hkwnv6);
assign Hkwnv6 = (~(Ii47v6 & Okwnv6));
assign Akwnv6 = (Vkwnv6 & Clwnv6);
assign Clwnv6 = (~(Uixmz6[31] & Jlwnv6));
assign Vkwnv6 = (~(Coxmz6[31] & Qlwnv6));
assign Mjwnv6 = (Xlwnv6 & Emwnv6);
assign Emwnv6 = (~(L5ymz6[34] & Lmwnv6));
assign Xlwnv6 = (~(TDI & Smwnv6));
assign Ztl8v6 = (Zmwnv6 ? U3o7z6[31] : Mcwnv6);
assign Stl8v6 = (~(Gnwnv6 & Nnwnv6));
assign Nnwnv6 = (~(Unwnv6 & Bownv6));
assign Gnwnv6 = (~(Iownv6 & Dtm7z6[2]));
assign Ltl8v6 = (~(Pownv6 & Wownv6));
assign Wownv6 = (~(Dpwnv6 & Itb7z6[0]));
assign Pownv6 = (Kpwnv6 & Rpwnv6);
assign Rpwnv6 = (~(Ypwnv6 & Fqwnv6));
assign Ypwnv6 = (~(Mqwnv6 & Tqwnv6));
assign Tqwnv6 = (Arwnv6 & Hrwnv6);
assign Hrwnv6 = (~(Dtm7z6[3] & Orwnv6));
assign Arwnv6 = (Wawnv6 | Vrwnv6);
assign Mqwnv6 = (Cswnv6 & Jswnv6);
assign Jswnv6 = (~(Dtm7z6[0] & HRDATAD[0]));
assign Cswnv6 = (~(Dtm7z6[1] & HRDATAS[0]));
assign Kpwnv6 = (~(Fcwnv6 & Qswnv6));
assign Etl8v6 = (~(Xswnv6 & Etwnv6));
assign Etwnv6 = (Ltwnv6 & Stwnv6);
assign Stwnv6 = (~(Ztwnv6 & Kxb7z6[31]));
assign Ltwnv6 = (Guwnv6 & Nuwnv6);
assign Nuwnv6 = (~(Uuwnv6 & Bvwnv6));
assign Guwnv6 = (~(Ivwnv6 & Fhc7z6[31]));
assign Xswnv6 = (Pvwnv6 & Wvwnv6);
assign Wvwnv6 = (~(Dwwnv6 & Nqh7z6[31]));
assign Pvwnv6 = (~(Kwwnv6 & Fth7z6[31]));
assign Xsl8v6 = (~(Rwwnv6 & Ywwnv6));
assign Ywwnv6 = (Fxwnv6 & Mxwnv6);
assign Mxwnv6 = (Txwnv6 & Aywnv6);
assign Txwnv6 = (~(Hywnv6 & Bvwnv6));
assign Fxwnv6 = (Oywnv6 & Vywnv6);
assign Vywnv6 = (~(Czwnv6 & Fhc7z6[31]));
assign Oywnv6 = (~(Jzwnv6 & Pic7z6[31]));
assign Rwwnv6 = (Qzwnv6 & Xzwnv6);
assign Xzwnv6 = (E0xnv6 & L0xnv6);
assign L0xnv6 = (S0xnv6 | Z0xnv6);
assign E0xnv6 = (~(G1xnv6 & N1xnv6));
assign Qzwnv6 = (U1xnv6 & B2xnv6);
assign B2xnv6 = (~(I2xnv6 & P2xnv6));
assign U1xnv6 = (~(W2xnv6 & Pdc7z6[31]));
assign Qsl8v6 = (~(D3xnv6 & Dconv6));
assign Jsl8v6 = (~(K3xnv6 & R3xnv6));
assign R3xnv6 = (~(D3xnv6 & Y3xnv6));
assign D3xnv6 = (!F4xnv6);
assign K3xnv6 = (~(Ujnet6 & M4xnv6));
assign Csl8v6 = (~(T4xnv6 & A5xnv6));
assign A5xnv6 = (~(H5xnv6 & Ujnet6));
assign T4xnv6 = (~(O5xnv6 & L9d7z6[5]));
assign Vrl8v6 = (~(V5xnv6 & C6xnv6));
assign C6xnv6 = (~(J6xnv6 & Q6xnv6));
assign Q6xnv6 = (Dxvnv6 & X6xnv6);
assign J6xnv6 = (Geddt6 & E7xnv6);
assign E7xnv6 = (~(L7xnv6 & K3jnv6));
assign V5xnv6 = (~(S7xnv6 & Q0wnv6));
assign S7xnv6 = (Z7xnv6 & G8xnv6);
assign Z7xnv6 = (!N8xnv6);
assign Orl8v6 = (~(U8xnv6 & B9xnv6));
assign B9xnv6 = (I9xnv6 & Aywnv6);
assign I9xnv6 = (~(G1xnv6 & P9xnv6));
assign U8xnv6 = (W9xnv6 & Daxnv6);
assign Daxnv6 = (~(I2xnv6 & Kaxnv6));
assign W9xnv6 = (~(Pdc7z6[0] & W2xnv6));
assign Hrl8v6 = (~(Raxnv6 & Yaxnv6));
assign Yaxnv6 = (Fbxnv6 & Mbxnv6);
assign Mbxnv6 = (Tbxnv6 & Aywnv6);
assign Tbxnv6 = (~(Hywnv6 & Acxnv6));
assign Fbxnv6 = (Hcxnv6 & Ocxnv6);
assign Ocxnv6 = (~(Czwnv6 & Fhc7z6[30]));
assign Hcxnv6 = (~(Jzwnv6 & Pic7z6[30]));
assign Raxnv6 = (Vcxnv6 & Cdxnv6);
assign Cdxnv6 = (Jdxnv6 & Qdxnv6);
assign Qdxnv6 = (S0xnv6 | Xdxnv6);
assign Jdxnv6 = (~(G1xnv6 & Eexnv6));
assign Vcxnv6 = (Lexnv6 & Sexnv6);
assign Sexnv6 = (~(I2xnv6 & Zexnv6));
assign Lexnv6 = (~(W2xnv6 & Pdc7z6[30]));
assign Arl8v6 = (~(Gfxnv6 & Nfxnv6));
assign Nfxnv6 = (Ufxnv6 & Bgxnv6);
assign Bgxnv6 = (Igxnv6 & Aywnv6);
assign Igxnv6 = (~(Hywnv6 & Pgxnv6));
assign Ufxnv6 = (Wgxnv6 & Dhxnv6);
assign Dhxnv6 = (~(Czwnv6 & Fhc7z6[29]));
assign Wgxnv6 = (~(Jzwnv6 & Pic7z6[29]));
assign Gfxnv6 = (Khxnv6 & Rhxnv6);
assign Rhxnv6 = (Yhxnv6 & Fixnv6);
assign Fixnv6 = (S0xnv6 | Mixnv6);
assign Yhxnv6 = (~(G1xnv6 & Tixnv6));
assign Khxnv6 = (Ajxnv6 & Hjxnv6);
assign Hjxnv6 = (~(I2xnv6 & Ojxnv6));
assign Ajxnv6 = (~(W2xnv6 & Pdc7z6[29]));
assign Tql8v6 = (~(Vjxnv6 & Ckxnv6));
assign Ckxnv6 = (Jkxnv6 & Qkxnv6);
assign Qkxnv6 = (Xkxnv6 & Aywnv6);
assign Xkxnv6 = (~(Hywnv6 & Elxnv6));
assign Jkxnv6 = (Llxnv6 & Slxnv6);
assign Slxnv6 = (~(Czwnv6 & Fhc7z6[28]));
assign Llxnv6 = (~(Jzwnv6 & Pic7z6[28]));
assign Vjxnv6 = (Zlxnv6 & Gmxnv6);
assign Gmxnv6 = (Nmxnv6 & Umxnv6);
assign Umxnv6 = (S0xnv6 | Bnxnv6);
assign Nmxnv6 = (~(G1xnv6 & Inxnv6));
assign Zlxnv6 = (Pnxnv6 & Wnxnv6);
assign Wnxnv6 = (~(I2xnv6 & Doxnv6));
assign Pnxnv6 = (~(W2xnv6 & Pdc7z6[28]));
assign Mql8v6 = (~(Koxnv6 & Roxnv6));
assign Roxnv6 = (Yoxnv6 & Fpxnv6);
assign Fpxnv6 = (Mpxnv6 & Aywnv6);
assign Mpxnv6 = (~(Hywnv6 & Tpxnv6));
assign Yoxnv6 = (Aqxnv6 & Hqxnv6);
assign Hqxnv6 = (~(Czwnv6 & Fhc7z6[27]));
assign Aqxnv6 = (~(Jzwnv6 & Pic7z6[27]));
assign Koxnv6 = (Oqxnv6 & Vqxnv6);
assign Vqxnv6 = (Crxnv6 & Jrxnv6);
assign Jrxnv6 = (S0xnv6 | Qrxnv6);
assign Crxnv6 = (~(G1xnv6 & Xrxnv6));
assign Oqxnv6 = (Esxnv6 & Lsxnv6);
assign Lsxnv6 = (~(I2xnv6 & Ssxnv6));
assign Esxnv6 = (~(W2xnv6 & Pdc7z6[27]));
assign Fql8v6 = (~(Zsxnv6 & Gtxnv6));
assign Gtxnv6 = (Ntxnv6 & Utxnv6);
assign Utxnv6 = (Buxnv6 & Aywnv6);
assign Buxnv6 = (~(Hywnv6 & Iuxnv6));
assign Ntxnv6 = (Puxnv6 & Wuxnv6);
assign Wuxnv6 = (~(Czwnv6 & Fhc7z6[26]));
assign Puxnv6 = (~(Jzwnv6 & Pic7z6[26]));
assign Zsxnv6 = (Dvxnv6 & Kvxnv6);
assign Kvxnv6 = (Rvxnv6 & Yvxnv6);
assign Yvxnv6 = (S0xnv6 | Fwxnv6);
assign Rvxnv6 = (~(G1xnv6 & Mwxnv6));
assign Dvxnv6 = (Twxnv6 & Axxnv6);
assign Axxnv6 = (~(I2xnv6 & Hxxnv6));
assign Twxnv6 = (~(W2xnv6 & Pdc7z6[26]));
assign Ypl8v6 = (~(Oxxnv6 & Vxxnv6));
assign Vxxnv6 = (Cyxnv6 & Jyxnv6);
assign Jyxnv6 = (Qyxnv6 & Aywnv6);
assign Qyxnv6 = (~(Hywnv6 & Xyxnv6));
assign Cyxnv6 = (Ezxnv6 & Lzxnv6);
assign Lzxnv6 = (~(Czwnv6 & Fhc7z6[25]));
assign Ezxnv6 = (~(Jzwnv6 & Pic7z6[25]));
assign Oxxnv6 = (Szxnv6 & Zzxnv6);
assign Zzxnv6 = (G0ynv6 & N0ynv6);
assign N0ynv6 = (S0xnv6 | U0ynv6);
assign G0ynv6 = (~(G1xnv6 & B1ynv6));
assign Szxnv6 = (I1ynv6 & P1ynv6);
assign P1ynv6 = (~(I2xnv6 & W1ynv6));
assign I1ynv6 = (~(W2xnv6 & Pdc7z6[25]));
assign Rpl8v6 = (~(D2ynv6 & K2ynv6));
assign K2ynv6 = (R2ynv6 & Y2ynv6);
assign Y2ynv6 = (F3ynv6 & Aywnv6);
assign F3ynv6 = (~(Hywnv6 & M3ynv6));
assign R2ynv6 = (T3ynv6 & A4ynv6);
assign A4ynv6 = (~(Czwnv6 & Fhc7z6[24]));
assign T3ynv6 = (~(Jzwnv6 & Pic7z6[24]));
assign D2ynv6 = (H4ynv6 & O4ynv6);
assign O4ynv6 = (V4ynv6 & C5ynv6);
assign C5ynv6 = (S0xnv6 | J5ynv6);
assign V4ynv6 = (~(G1xnv6 & Kaxnv6));
assign H4ynv6 = (Q5ynv6 & X5ynv6);
assign X5ynv6 = (~(I2xnv6 & P9xnv6));
assign Q5ynv6 = (~(W2xnv6 & Pdc7z6[24]));
assign Kpl8v6 = (~(E6ynv6 & L6ynv6));
assign L6ynv6 = (S6ynv6 & Z6ynv6);
assign Z6ynv6 = (G7ynv6 & Aywnv6);
assign G7ynv6 = (~(Hywnv6 & N7ynv6));
assign S6ynv6 = (U7ynv6 & B8ynv6);
assign B8ynv6 = (~(Czwnv6 & Fhc7z6[23]));
assign U7ynv6 = (~(Jzwnv6 & Pic7z6[23]));
assign E6ynv6 = (I8ynv6 & P8ynv6);
assign P8ynv6 = (W8ynv6 & D9ynv6);
assign D9ynv6 = (S0xnv6 | K9ynv6);
assign W8ynv6 = (~(G1xnv6 & R9ynv6));
assign I8ynv6 = (Y9ynv6 & Faynv6);
assign Faynv6 = (~(I2xnv6 & Maynv6));
assign Y9ynv6 = (~(W2xnv6 & Pdc7z6[23]));
assign Dpl8v6 = (~(Taynv6 & Abynv6));
assign Abynv6 = (Hbynv6 & Obynv6);
assign Obynv6 = (Vbynv6 & Aywnv6);
assign Vbynv6 = (~(Hywnv6 & Ccynv6));
assign Hbynv6 = (Jcynv6 & Qcynv6);
assign Qcynv6 = (~(Czwnv6 & Fhc7z6[22]));
assign Jcynv6 = (~(Jzwnv6 & Pic7z6[22]));
assign Taynv6 = (Xcynv6 & Edynv6);
assign Edynv6 = (Ldynv6 & Sdynv6);
assign Sdynv6 = (S0xnv6 | Zdynv6);
assign Ldynv6 = (~(G1xnv6 & Geynv6));
assign Xcynv6 = (Neynv6 & Ueynv6);
assign Ueynv6 = (~(I2xnv6 & Bfynv6));
assign Neynv6 = (~(W2xnv6 & Pdc7z6[22]));
assign Wol8v6 = (~(Ifynv6 & Pfynv6));
assign Pfynv6 = (Wfynv6 & Dgynv6);
assign Dgynv6 = (Kgynv6 & Aywnv6);
assign Kgynv6 = (~(Hywnv6 & Rgynv6));
assign Wfynv6 = (Ygynv6 & Fhynv6);
assign Fhynv6 = (~(Czwnv6 & Fhc7z6[21]));
assign Ygynv6 = (~(Jzwnv6 & Pic7z6[21]));
assign Ifynv6 = (Mhynv6 & Thynv6);
assign Thynv6 = (Aiynv6 & Hiynv6);
assign Hiynv6 = (S0xnv6 | Oiynv6);
assign Aiynv6 = (~(G1xnv6 & Viynv6));
assign Mhynv6 = (Cjynv6 & Jjynv6);
assign Jjynv6 = (~(I2xnv6 & Qjynv6));
assign Cjynv6 = (~(W2xnv6 & Pdc7z6[21]));
assign Pol8v6 = (~(Xjynv6 & Ekynv6));
assign Ekynv6 = (Lkynv6 & Skynv6);
assign Skynv6 = (Zkynv6 & Aywnv6);
assign Zkynv6 = (~(Hywnv6 & Glynv6));
assign Lkynv6 = (Nlynv6 & Ulynv6);
assign Ulynv6 = (~(Czwnv6 & Fhc7z6[20]));
assign Nlynv6 = (~(Jzwnv6 & Pic7z6[20]));
assign Xjynv6 = (Bmynv6 & Imynv6);
assign Imynv6 = (Pmynv6 & Wmynv6);
assign Wmynv6 = (S0xnv6 | Dnynv6);
assign Pmynv6 = (~(G1xnv6 & Knynv6));
assign Bmynv6 = (Rnynv6 & Ynynv6);
assign Ynynv6 = (~(I2xnv6 & Foynv6));
assign Rnynv6 = (~(W2xnv6 & Pdc7z6[20]));
assign Iol8v6 = (~(Moynv6 & Toynv6));
assign Toynv6 = (Apynv6 & Hpynv6);
assign Hpynv6 = (Opynv6 & Aywnv6);
assign Opynv6 = (~(Hywnv6 & Vpynv6));
assign Apynv6 = (Cqynv6 & Jqynv6);
assign Jqynv6 = (~(Czwnv6 & Fhc7z6[19]));
assign Cqynv6 = (~(Jzwnv6 & Pic7z6[19]));
assign Moynv6 = (Qqynv6 & Xqynv6);
assign Xqynv6 = (Erynv6 & Lrynv6);
assign Lrynv6 = (S0xnv6 | Srynv6);
assign Erynv6 = (~(G1xnv6 & Zrynv6));
assign Qqynv6 = (Gsynv6 & Nsynv6);
assign Nsynv6 = (~(I2xnv6 & Usynv6));
assign Gsynv6 = (~(W2xnv6 & Pdc7z6[19]));
assign Bol8v6 = (~(Btynv6 & Itynv6));
assign Itynv6 = (Ptynv6 & Wtynv6);
assign Wtynv6 = (Duynv6 & Aywnv6);
assign Duynv6 = (~(Hywnv6 & Kuynv6));
assign Ptynv6 = (Ruynv6 & Yuynv6);
assign Yuynv6 = (~(Czwnv6 & Fhc7z6[18]));
assign Ruynv6 = (~(Jzwnv6 & Pic7z6[18]));
assign Btynv6 = (Fvynv6 & Mvynv6);
assign Mvynv6 = (Tvynv6 & Awynv6);
assign Awynv6 = (S0xnv6 | Hwynv6);
assign Tvynv6 = (~(G1xnv6 & Owynv6));
assign Fvynv6 = (Vwynv6 & Cxynv6);
assign Cxynv6 = (~(I2xnv6 & Jxynv6));
assign Vwynv6 = (~(W2xnv6 & Pdc7z6[18]));
assign Unl8v6 = (~(Qxynv6 & Xxynv6));
assign Xxynv6 = (Eyynv6 & Lyynv6);
assign Lyynv6 = (Syynv6 & Aywnv6);
assign Syynv6 = (~(Hywnv6 & Zyynv6));
assign Eyynv6 = (Gzynv6 & Nzynv6);
assign Nzynv6 = (~(Czwnv6 & Fhc7z6[17]));
assign Gzynv6 = (~(Jzwnv6 & Pic7z6[17]));
assign Qxynv6 = (Uzynv6 & B0znv6);
assign B0znv6 = (I0znv6 & P0znv6);
assign P0znv6 = (S0xnv6 | W0znv6);
assign I0znv6 = (~(G1xnv6 & D1znv6));
assign Uzynv6 = (K1znv6 & R1znv6);
assign R1znv6 = (~(I2xnv6 & Y1znv6));
assign K1znv6 = (~(W2xnv6 & Pdc7z6[17]));
assign Nnl8v6 = (~(F2znv6 & M2znv6));
assign M2znv6 = (T2znv6 & A3znv6);
assign A3znv6 = (H3znv6 & Aywnv6);
assign H3znv6 = (~(Hywnv6 & O3znv6));
assign T2znv6 = (V3znv6 & C4znv6);
assign C4znv6 = (~(Czwnv6 & Fhc7z6[16]));
assign V3znv6 = (~(Jzwnv6 & Pic7z6[16]));
assign F2znv6 = (J4znv6 & Q4znv6);
assign Q4znv6 = (X4znv6 & E5znv6);
assign E5znv6 = (S0xnv6 | L5znv6);
assign X4znv6 = (~(G1xnv6 & S5znv6));
assign J4znv6 = (Z5znv6 & G6znv6);
assign G6znv6 = (~(I2xnv6 & N6znv6));
assign Z5znv6 = (~(W2xnv6 & Pdc7z6[16]));
assign Gnl8v6 = (~(U6znv6 & B7znv6));
assign B7znv6 = (I7znv6 & P7znv6);
assign P7znv6 = (W7znv6 & Aywnv6);
assign W7znv6 = (~(Hywnv6 & D8znv6));
assign I7znv6 = (K8znv6 & R8znv6);
assign R8znv6 = (~(Czwnv6 & Fhc7z6[15]));
assign K8znv6 = (~(Jzwnv6 & Pic7z6[15]));
assign U6znv6 = (Y8znv6 & F9znv6);
assign F9znv6 = (M9znv6 & T9znv6);
assign T9znv6 = (S0xnv6 | Aaznv6);
assign M9znv6 = (~(G1xnv6 & Maynv6));
assign Y8znv6 = (Haznv6 & Oaznv6);
assign Oaznv6 = (~(I2xnv6 & R9ynv6));
assign Haznv6 = (~(W2xnv6 & Pdc7z6[15]));
assign Zml8v6 = (~(Vaznv6 & Cbznv6));
assign Cbznv6 = (Jbznv6 & Qbznv6);
assign Qbznv6 = (Xbznv6 & Aywnv6);
assign Xbznv6 = (~(Hywnv6 & Ecznv6));
assign Jbznv6 = (Lcznv6 & Scznv6);
assign Scznv6 = (~(Czwnv6 & Fhc7z6[14]));
assign Lcznv6 = (~(Jzwnv6 & Pic7z6[14]));
assign Vaznv6 = (Zcznv6 & Gdznv6);
assign Gdznv6 = (Ndznv6 & Udznv6);
assign Udznv6 = (S0xnv6 | Beznv6);
assign Ndznv6 = (~(G1xnv6 & Bfynv6));
assign Zcznv6 = (Ieznv6 & Peznv6);
assign Peznv6 = (~(I2xnv6 & Geynv6));
assign Ieznv6 = (~(W2xnv6 & Pdc7z6[14]));
assign Sml8v6 = (~(Weznv6 & Dfznv6));
assign Dfznv6 = (Kfznv6 & Rfznv6);
assign Rfznv6 = (Yfznv6 & Aywnv6);
assign Yfznv6 = (~(Hywnv6 & Fgznv6));
assign Kfznv6 = (Mgznv6 & Tgznv6);
assign Tgznv6 = (~(Czwnv6 & Fhc7z6[13]));
assign Mgznv6 = (~(Jzwnv6 & Pic7z6[13]));
assign Weznv6 = (Ahznv6 & Hhznv6);
assign Hhznv6 = (Ohznv6 & Vhznv6);
assign Vhznv6 = (S0xnv6 | Ciznv6);
assign Ohznv6 = (~(G1xnv6 & Qjynv6));
assign Ahznv6 = (Jiznv6 & Qiznv6);
assign Qiznv6 = (~(I2xnv6 & Viynv6));
assign Jiznv6 = (~(W2xnv6 & Pdc7z6[13]));
assign Lml8v6 = (~(Xiznv6 & Ejznv6));
assign Ejznv6 = (Ljznv6 & Sjznv6);
assign Sjznv6 = (Zjznv6 & Aywnv6);
assign Zjznv6 = (~(Hywnv6 & Gkznv6));
assign Ljznv6 = (Nkznv6 & Ukznv6);
assign Ukznv6 = (~(Czwnv6 & Fhc7z6[12]));
assign Nkznv6 = (~(Jzwnv6 & Pic7z6[12]));
assign Xiznv6 = (Blznv6 & Ilznv6);
assign Ilznv6 = (Plznv6 & Wlznv6);
assign Wlznv6 = (S0xnv6 | Dmznv6);
assign Plznv6 = (~(G1xnv6 & Foynv6));
assign Blznv6 = (Kmznv6 & Rmznv6);
assign Rmznv6 = (~(I2xnv6 & Knynv6));
assign Kmznv6 = (~(W2xnv6 & Pdc7z6[12]));
assign Eml8v6 = (~(Ymznv6 & Fnznv6));
assign Fnznv6 = (Mnznv6 & Tnznv6);
assign Tnznv6 = (Aoznv6 & Aywnv6);
assign Aoznv6 = (~(Hywnv6 & Hoznv6));
assign Mnznv6 = (Ooznv6 & Voznv6);
assign Voznv6 = (~(Czwnv6 & Fhc7z6[11]));
assign Ooznv6 = (~(Jzwnv6 & Pic7z6[11]));
assign Ymznv6 = (Cpznv6 & Jpznv6);
assign Jpznv6 = (Qpznv6 & Xpznv6);
assign Xpznv6 = (S0xnv6 | Eqznv6);
assign Qpznv6 = (~(G1xnv6 & Usynv6));
assign Cpznv6 = (Lqznv6 & Sqznv6);
assign Sqznv6 = (~(I2xnv6 & Zrynv6));
assign Lqznv6 = (~(W2xnv6 & Pdc7z6[11]));
assign Xll8v6 = (~(Zqznv6 & Grznv6));
assign Grznv6 = (Nrznv6 & Urznv6);
assign Urznv6 = (Bsznv6 & Aywnv6);
assign Bsznv6 = (~(Hywnv6 & Isznv6));
assign Nrznv6 = (Psznv6 & Wsznv6);
assign Wsznv6 = (~(Czwnv6 & Fhc7z6[10]));
assign Psznv6 = (~(Jzwnv6 & Pic7z6[10]));
assign Zqznv6 = (Dtznv6 & Ktznv6);
assign Ktznv6 = (Rtznv6 & Ytznv6);
assign Ytznv6 = (S0xnv6 | Fuznv6);
assign Rtznv6 = (~(G1xnv6 & Jxynv6));
assign Dtznv6 = (Muznv6 & Tuznv6);
assign Tuznv6 = (~(I2xnv6 & Owynv6));
assign Muznv6 = (~(W2xnv6 & Pdc7z6[10]));
assign Qll8v6 = (~(Avznv6 & Hvznv6));
assign Hvznv6 = (Ovznv6 & Vvznv6);
assign Vvznv6 = (Cwznv6 & Aywnv6);
assign Cwznv6 = (~(Hywnv6 & Jwznv6));
assign Ovznv6 = (Qwznv6 & Xwznv6);
assign Xwznv6 = (~(Czwnv6 & Fhc7z6[9]));
assign Qwznv6 = (~(Jzwnv6 & Pic7z6[9]));
assign Avznv6 = (Exznv6 & Lxznv6);
assign Lxznv6 = (Sxznv6 & Zxznv6);
assign Zxznv6 = (S0xnv6 | Gyznv6);
assign Sxznv6 = (~(G1xnv6 & Y1znv6));
assign Exznv6 = (Nyznv6 & Uyznv6);
assign Uyznv6 = (~(I2xnv6 & D1znv6));
assign Nyznv6 = (~(W2xnv6 & Pdc7z6[9]));
assign Jll8v6 = (~(Bzznv6 & Izznv6));
assign Izznv6 = (Pzznv6 & Wzznv6);
assign Wzznv6 = (D00ov6 & Aywnv6);
assign D00ov6 = (~(Hywnv6 & K00ov6));
assign Pzznv6 = (R00ov6 & Y00ov6);
assign Y00ov6 = (~(Czwnv6 & Fhc7z6[8]));
assign R00ov6 = (~(Jzwnv6 & Pic7z6[8]));
assign Bzznv6 = (F10ov6 & M10ov6);
assign M10ov6 = (T10ov6 & A20ov6);
assign A20ov6 = (S0xnv6 | H20ov6);
assign T10ov6 = (~(G1xnv6 & N6znv6));
assign F10ov6 = (O20ov6 & V20ov6);
assign V20ov6 = (~(I2xnv6 & S5znv6));
assign O20ov6 = (~(W2xnv6 & Pdc7z6[8]));
assign Cll8v6 = (~(C30ov6 & J30ov6));
assign J30ov6 = (Q30ov6 & X30ov6);
assign X30ov6 = (E40ov6 & Aywnv6);
assign E40ov6 = (~(Hywnv6 & L40ov6));
assign Q30ov6 = (S40ov6 & Z40ov6);
assign Z40ov6 = (~(Czwnv6 & Fhc7z6[7]));
assign S40ov6 = (~(Jzwnv6 & Pic7z6[7]));
assign C30ov6 = (G50ov6 & N50ov6);
assign N50ov6 = (U50ov6 & B60ov6);
assign B60ov6 = (S0xnv6 | I60ov6);
assign U50ov6 = (~(G1xnv6 & P2xnv6));
assign G50ov6 = (P60ov6 & W60ov6);
assign W60ov6 = (~(I2xnv6 & N1xnv6));
assign P60ov6 = (~(W2xnv6 & Pdc7z6[7]));
assign Vkl8v6 = (~(D70ov6 & K70ov6));
assign K70ov6 = (R70ov6 & Y70ov6);
assign Y70ov6 = (F80ov6 & Aywnv6);
assign F80ov6 = (~(Hywnv6 & M80ov6));
assign R70ov6 = (T80ov6 & A90ov6);
assign A90ov6 = (~(Czwnv6 & Fhc7z6[6]));
assign T80ov6 = (~(Jzwnv6 & Pic7z6[6]));
assign D70ov6 = (H90ov6 & O90ov6);
assign O90ov6 = (V90ov6 & Ca0ov6);
assign Ca0ov6 = (S0xnv6 | Ja0ov6);
assign V90ov6 = (~(G1xnv6 & Zexnv6));
assign H90ov6 = (Qa0ov6 & Xa0ov6);
assign Xa0ov6 = (~(I2xnv6 & Eexnv6));
assign Qa0ov6 = (~(W2xnv6 & Pdc7z6[6]));
assign Okl8v6 = (~(Eb0ov6 & Lb0ov6));
assign Lb0ov6 = (Sb0ov6 & Zb0ov6);
assign Zb0ov6 = (Gc0ov6 & Aywnv6);
assign Gc0ov6 = (~(Hywnv6 & Nc0ov6));
assign Sb0ov6 = (Uc0ov6 & Bd0ov6);
assign Bd0ov6 = (~(Czwnv6 & Fhc7z6[5]));
assign Uc0ov6 = (~(Jzwnv6 & Pic7z6[5]));
assign Eb0ov6 = (Id0ov6 & Pd0ov6);
assign Pd0ov6 = (Wd0ov6 & De0ov6);
assign De0ov6 = (S0xnv6 | Ke0ov6);
assign Wd0ov6 = (~(G1xnv6 & Ojxnv6));
assign Id0ov6 = (Re0ov6 & Ye0ov6);
assign Ye0ov6 = (~(I2xnv6 & Tixnv6));
assign Re0ov6 = (~(W2xnv6 & Pdc7z6[5]));
assign Hkl8v6 = (~(Ff0ov6 & Mf0ov6));
assign Mf0ov6 = (Tf0ov6 & Ag0ov6);
assign Ag0ov6 = (Hg0ov6 & Aywnv6);
assign Hg0ov6 = (~(Hywnv6 & Og0ov6));
assign Tf0ov6 = (Vg0ov6 & Ch0ov6);
assign Ch0ov6 = (~(Czwnv6 & E3c7z6[4]));
assign Vg0ov6 = (~(Jzwnv6 & Pic7z6[4]));
assign Ff0ov6 = (Jh0ov6 & Qh0ov6);
assign Qh0ov6 = (Xh0ov6 & Ei0ov6);
assign Ei0ov6 = (S0xnv6 | Li0ov6);
assign Xh0ov6 = (~(G1xnv6 & Doxnv6));
assign Jh0ov6 = (Si0ov6 & Zi0ov6);
assign Zi0ov6 = (~(I2xnv6 & Inxnv6));
assign Si0ov6 = (~(W2xnv6 & Pdc7z6[4]));
assign Akl8v6 = (~(Gj0ov6 & Nj0ov6));
assign Nj0ov6 = (Uj0ov6 & Bk0ov6);
assign Bk0ov6 = (Ik0ov6 & Aywnv6);
assign Ik0ov6 = (~(Hywnv6 & Pk0ov6));
assign Uj0ov6 = (Wk0ov6 & Dl0ov6);
assign Dl0ov6 = (~(Czwnv6 & E3c7z6[3]));
assign Wk0ov6 = (~(Jzwnv6 & Pic7z6[3]));
assign Gj0ov6 = (Kl0ov6 & Rl0ov6);
assign Rl0ov6 = (Yl0ov6 & Fm0ov6);
assign Fm0ov6 = (S0xnv6 | Mm0ov6);
assign Yl0ov6 = (~(G1xnv6 & Ssxnv6));
assign Kl0ov6 = (Tm0ov6 & An0ov6);
assign An0ov6 = (~(I2xnv6 & Xrxnv6));
assign Tm0ov6 = (~(W2xnv6 & Pdc7z6[3]));
assign Tjl8v6 = (~(Hn0ov6 & On0ov6));
assign On0ov6 = (Vn0ov6 & Co0ov6);
assign Co0ov6 = (Jo0ov6 & Aywnv6);
assign Jo0ov6 = (~(Hywnv6 & Qo0ov6));
assign Hywnv6 = (Xo0ov6 & Ep0ov6);
assign Xo0ov6 = (~(W2xnv6 | Lp0ov6));
assign Vn0ov6 = (Sp0ov6 & Zp0ov6);
assign Zp0ov6 = (~(Czwnv6 & E3c7z6[2]));
assign Czwnv6 = (Gq0ov6 & Nq0ov6);
assign Gq0ov6 = (Lp0ov6 & Qdcdt6);
assign Sp0ov6 = (~(Jzwnv6 & Pic7z6[2]));
assign Jzwnv6 = (Uq0ov6 & Nq0ov6);
assign Nq0ov6 = (Ep0ov6 & Br0ov6);
assign Uq0ov6 = (Lp0ov6 & Ir0ov6);
assign Hn0ov6 = (Pr0ov6 & Wr0ov6);
assign Wr0ov6 = (Ds0ov6 & Ks0ov6);
assign Ks0ov6 = (S0xnv6 | Rs0ov6);
assign S0xnv6 = (~(Ys0ov6 & Br0ov6));
assign Ys0ov6 = (Ft0ov6 | Mt0ov6);
assign Mt0ov6 = (Tt0ov6 & Au0ov6);
assign Tt0ov6 = (Lp0ov6 & Ep0ov6);
assign Ep0ov6 = (~(Hu0ov6 & Ou0ov6));
assign Ou0ov6 = (~(Vu0ov6 & Cv0ov6));
assign Cv0ov6 = (~(Jv0ov6 & Qv0ov6));
assign Ds0ov6 = (~(G1xnv6 & Hxxnv6));
assign Pr0ov6 = (Xv0ov6 & Ew0ov6);
assign Ew0ov6 = (~(I2xnv6 & Mwxnv6));
assign Xv0ov6 = (~(W2xnv6 & Pdc7z6[2]));
assign Mjl8v6 = (~(Lw0ov6 & Sw0ov6));
assign Sw0ov6 = (Zw0ov6 & Aywnv6);
assign Aywnv6 = (~(Gx0ov6 & Br0ov6));
assign Gx0ov6 = (~(Nx0ov6 & Ux0ov6));
assign Ux0ov6 = (~(Sgcdt6 & By0ov6));
assign Zw0ov6 = (~(G1xnv6 & W1ynv6));
assign G1xnv6 = (Iy0ov6 & Evadt6);
assign Iy0ov6 = (Br0ov6 & By0ov6);
assign Lw0ov6 = (Py0ov6 & Wy0ov6);
assign Wy0ov6 = (~(I2xnv6 & B1ynv6));
assign I2xnv6 = (Dz0ov6 & Br0ov6);
assign Dz0ov6 = (By0ov6 & Euonv6);
assign Py0ov6 = (~(W2xnv6 & Pdc7z6[1]));
assign W2xnv6 = (!Br0ov6);
assign Br0ov6 = (~(Kz0ov6 & Rz0ov6));
assign Rz0ov6 = (Yz0ov6 & F01ov6);
assign F01ov6 = (~(M01ov6 & Vu0ov6));
assign M01ov6 = (Q0wnv6 & T01ov6);
assign T01ov6 = (~(Qv0ov6 & A11ov6));
assign Yz0ov6 = (~(H11ov6 & O11ov6));
assign O11ov6 = (~(Nx0ov6 & V11ov6));
assign V11ov6 = (~(Ywcdt6 & By0ov6));
assign By0ov6 = (C21ov6 | J21ov6);
assign Kz0ov6 = (Q21ov6 & X21ov6);
assign X21ov6 = (~(Ft0ov6 & E31ov6));
assign Ft0ov6 = (L31ov6 & S31ov6);
assign S31ov6 = (Z31ov6 & Jv0ov6);
assign Z31ov6 = (Ldo7v6 & Qv0ov6);
assign L31ov6 = (G41ov6 & Vu0ov6);
assign Vu0ov6 = (N41ov6 & U41ov6);
assign U41ov6 = (~(B51ov6 | I51ov6));
assign N41ov6 = (P51ov6 & W51ov6);
assign Q21ov6 = (Hu0ov6 | D61ov6);
assign Fjl8v6 = (~(K61ov6 & R61ov6));
assign R61ov6 = (Y61ov6 & F71ov6);
assign F71ov6 = (M71ov6 & T71ov6);
assign T71ov6 = (~(A81ov6 & Y9o7v6));
assign M71ov6 = (H81ov6 & O81ov6);
assign O81ov6 = (~(Byc7z6[15] & V81ov6));
assign H81ov6 = (~(C91ov6 & R9ynv6));
assign Y61ov6 = (J91ov6 & Q91ov6);
assign Q91ov6 = (~(X91ov6 & Fao7v6));
assign J91ov6 = (~(Ea1ov6 & W8o7v6));
assign K61ov6 = (La1ov6 & Sa1ov6);
assign Sa1ov6 = (Za1ov6 & Gb1ov6);
assign Gb1ov6 = (~(Nb1ov6 & P8o7v6));
assign Za1ov6 = (~(Byc7z6[31] & Ub1ov6));
assign La1ov6 = (Bc1ov6 & Ic1ov6);
assign Ic1ov6 = (~(Pc1ov6 & P2xnv6));
assign Bc1ov6 = (~(Zec7z6[31] & Wc1ov6));
assign Yil8v6 = (~(Dd1ov6 ^ Kd1ov6));
assign Dd1ov6 = (~(Rd1ov6 & Yd1ov6));
assign Yd1ov6 = (~(Wzcdt6 & Fe1ov6));
assign Fe1ov6 = (~(Me1ov6 & Te1ov6));
assign Te1ov6 = (A11ov6 | G41ov6);
assign A11ov6 = (~(A9mnv6 & Af1ov6));
assign Rd1ov6 = (Hf1ov6 & Of1ov6);
assign Of1ov6 = (~(Vf1ov6 & Cg1ov6));
assign Vf1ov6 = (Jv0ov6 & Jg1ov6);
assign Jg1ov6 = (~(Qg1ov6 & Xg1ov6));
assign Qg1ov6 = (Eh1ov6 & Lh1ov6);
assign Hf1ov6 = (~(Me1ov6 & Sh1ov6));
assign Sh1ov6 = (~(Zh1ov6 & Gi1ov6));
assign Gi1ov6 = (~(Ni1ov6 & Ui1ov6));
assign Ui1ov6 = (Af1ov6 ? A9mnv6 : Eh1ov6);
assign Ni1ov6 = (G41ov6 & Kd1ov6);
assign G41ov6 = (N8xnv6 & Lh1ov6);
assign Zh1ov6 = (Bj1ov6 | A9mnv6);
assign Bj1ov6 = (Ij1ov6 | Jv0ov6);
assign Me1ov6 = (Qv0ov6 & Pj1ov6);
assign Ril8v6 = (Aocdt6 | Wj1ov6);
assign Kil8v6 = (~(Dk1ov6 & Kk1ov6));
assign Kk1ov6 = (~(Rk1ov6 & Yk1ov6));
assign Rk1ov6 = (DNOTITRANS & Fl1ov6);
assign Dk1ov6 = (~(U4zet6 & Ml1ov6));
assign Ml1ov6 = (~(DNOTITRANS & Tl1ov6));
assign Tl1ov6 = (~(Am1ov6 & Fl1ov6));
assign Fl1ov6 = (!HREADYI);
assign Dil8v6 = (Om1ov6 ? Hm1ov6 : Ysn7z6[0]);
assign Whl8v6 = (Om1ov6 ? Vm1ov6 : Ysn7z6[1]);
assign Om1ov6 = (!Cn1ov6);
assign Phl8v6 = (Cn1ov6 ? Ysn7z6[2] : Jn1ov6);
assign Cn1ov6 = (~(Ihl8v6 | N7zet6));
assign Ihl8v6 = (HTRANSD[1] & Goonv6);
assign Bhl8v6 = (~(Qn1ov6 & Xn1ov6));
assign Xn1ov6 = (~(Qsinv6 & O5a7z6));
assign Qn1ov6 = (~(Wbxdt6 & Vrinv6));
assign Ugl8v6 = (Eo1ov6 & Lo1ov6);
assign Eo1ov6 = (Ir7et6 | So1ov6);
assign So1ov6 = (Zo1ov6 & Gp1ov6);
assign Ngl8v6 = (Np1ov6 | Up1ov6);
assign Up1ov6 = (Bq1ov6 & Iq1ov6);
assign Iq1ov6 = (Pq1ov6 | Y8uet6);
assign Pq1ov6 = (~(E2wet6 | Wq1ov6));
assign Wq1ov6 = (!Vbo7v6);
assign Np1ov6 = (Kr1ov6 ? Dr1ov6 : Tim7z6[31]);
assign Dr1ov6 = (~(Rr1ov6 & Yr1ov6));
assign Yr1ov6 = (~(Fs1ov6 & Itb7z6[31]));
assign Rr1ov6 = (Ms1ov6 & Ts1ov6);
assign Ts1ov6 = (~(At1ov6 & Vbo7v6));
assign Ms1ov6 = (~(Ht1ov6 & Ot1ov6));
assign Ggl8v6 = (~(Vt1ov6 & Cu1ov6));
assign Cu1ov6 = (~(Ju1ov6 & Qu1ov6));
assign Vt1ov6 = (Xu1ov6 & Uginv6);
assign Uginv6 = (~(Ev1ov6 & Lv1ov6));
assign Lv1ov6 = (Sv1ov6 | Mtkdt6);
assign Sv1ov6 = (Gw1ov6 ? Zv1ov6 : L0g7z6[31]);
assign Zv1ov6 = (~(Nw1ov6 & Uw1ov6));
assign Uw1ov6 = (Bx1ov6 & Ix1ov6);
assign Ix1ov6 = (~(Px1ov6 & Fhc7z6[31]));
assign Bx1ov6 = (~(Wx1ov6 & Dy1ov6));
assign Nw1ov6 = (Ky1ov6 & Ry1ov6);
assign Xu1ov6 = (~(O4gdt6 & Yy1ov6));
assign Zfl8v6 = (~(Fz1ov6 & Mz1ov6));
assign Mz1ov6 = (Tz1ov6 & A02ov6);
assign A02ov6 = (~(H02ov6 & Wt97z6));
assign Tz1ov6 = (O02ov6 & V02ov6);
assign V02ov6 = (C12ov6 | Ckjnv6);
assign Ckjnv6 = (J12ov6 & Q12ov6);
assign Q12ov6 = (X12ov6 & E22ov6);
assign E22ov6 = (L22ov6 & S22ov6);
assign S22ov6 = (Z22ov6 & G32ov6);
assign G32ov6 = (~(vis_psp_o[31] & N32ov6));
assign Z22ov6 = (~(U32ov6 & Pic7z6[31]));
assign L22ov6 = (B42ov6 & I42ov6);
assign I42ov6 = (~(vis_msp_o[31] & P42ov6));
assign B42ov6 = (~(vis_r12_o[31] & W42ov6));
assign X12ov6 = (D52ov6 & K52ov6);
assign K52ov6 = (R52ov6 & Y52ov6);
assign Y52ov6 = (~(vis_r11_o[31] & F62ov6));
assign R52ov6 = (~(vis_r10_o[31] & M62ov6));
assign D52ov6 = (T62ov6 & A72ov6);
assign A72ov6 = (~(vis_r9_o[31] & H72ov6));
assign T62ov6 = (~(vis_r8_o[31] & O72ov6));
assign J12ov6 = (V72ov6 & C82ov6);
assign C82ov6 = (J82ov6 & Q82ov6);
assign Q82ov6 = (X82ov6 & E92ov6);
assign E92ov6 = (~(vis_r7_o[31] & L92ov6));
assign X82ov6 = (~(vis_r6_o[31] & S92ov6));
assign J82ov6 = (Z92ov6 & Ga2ov6);
assign Ga2ov6 = (~(vis_r5_o[31] & Na2ov6));
assign Z92ov6 = (~(vis_r4_o[31] & Ua2ov6));
assign V72ov6 = (Bb2ov6 & Ib2ov6);
assign Ib2ov6 = (Pb2ov6 & Wb2ov6);
assign Wb2ov6 = (~(vis_r3_o[31] & Dc2ov6));
assign Pb2ov6 = (~(vis_r2_o[31] & Kc2ov6));
assign Bb2ov6 = (Rc2ov6 & Yc2ov6);
assign Yc2ov6 = (~(vis_r1_o[31] & Fd2ov6));
assign Rc2ov6 = (~(vis_r0_o[31] & Md2ov6));
assign O02ov6 = (~(Td2ov6 & Ae2ov6));
assign Fz1ov6 = (He2ov6 & Oe2ov6);
assign Oe2ov6 = (~(Ve2ov6 & vis_pc_o[31]));
assign He2ov6 = (~(Fhc7z6[31] & Cf2ov6));
assign Sfl8v6 = (Jf2ov6 & Qf2ov6);
assign Jf2ov6 = (Xf2ov6 & Eg2ov6);
assign Eg2ov6 = (!Lg2ov6);
assign Xf2ov6 = (~(Sg2ov6 & Zg2ov6));
assign Zg2ov6 = (~(Gh2ov6 & Nh2ov6));
assign Sg2ov6 = (~(Uh2ov6 & Bi2ov6));
assign Lfl8v6 = (~(Ii2ov6 & Pi2ov6));
assign Pi2ov6 = (Wi2ov6 | Zfg7z6[32]);
assign Ii2ov6 = (Dj2ov6 & Kj2ov6);
assign Kj2ov6 = (~(Rj2ov6 & Vimdt6));
assign Dj2ov6 = (~(Yj2ov6 & Yxf7z6[2]));
assign Efl8v6 = (~(Fk2ov6 & Mk2ov6));
assign Mk2ov6 = (~(Tk2ov6 & Qu1ov6));
assign Fk2ov6 = (Al2ov6 & Phinv6);
assign Phinv6 = (~(Ev1ov6 & Hl2ov6));
assign Hl2ov6 = (Ol2ov6 | Vl2ov6);
assign Vl2ov6 = (Jm2ov6 ? Iphdt6 : Cm2ov6);
assign Cm2ov6 = (~(Qm2ov6 & Xm2ov6));
assign Xm2ov6 = (En2ov6 & Ln2ov6);
assign Ln2ov6 = (~(Sn2ov6 & Zn2ov6));
assign Zn2ov6 = (Go2ov6 & No2ov6);
assign No2ov6 = (Uo2ov6 & Bp2ov6);
assign Bp2ov6 = (Ip2ov6 & Pp2ov6);
assign Pp2ov6 = (Wp2ov6 & Dq2ov6);
assign Wp2ov6 = (Kq2ov6 & Ky1ov6);
assign Ip2ov6 = (Rq2ov6 & Yq2ov6);
assign Uo2ov6 = (Fr2ov6 & Mr2ov6);
assign Mr2ov6 = (Tr2ov6 & As2ov6);
assign Fr2ov6 = (Hs2ov6 & Os2ov6);
assign Go2ov6 = (Vs2ov6 & Ct2ov6);
assign Ct2ov6 = (Jt2ov6 & Qt2ov6);
assign Qt2ov6 = (Xt2ov6 & Eu2ov6);
assign Jt2ov6 = (Lu2ov6 & Su2ov6);
assign Vs2ov6 = (Zu2ov6 & Gv2ov6);
assign Gv2ov6 = (Nv2ov6 & Uv2ov6);
assign Zu2ov6 = (Bw2ov6 & Iw2ov6);
assign Sn2ov6 = (Pw2ov6 & Ww2ov6);
assign Ww2ov6 = (Dx2ov6 & Kx2ov6);
assign Kx2ov6 = (Rx2ov6 & Yx2ov6);
assign Yx2ov6 = (Fy2ov6 & My2ov6);
assign Rx2ov6 = (Ty2ov6 & Az2ov6);
assign Dx2ov6 = (Hz2ov6 & Oz2ov6);
assign Oz2ov6 = (Vz2ov6 & C03ov6);
assign Hz2ov6 = (J03ov6 & Q03ov6);
assign Pw2ov6 = (X03ov6 & E13ov6);
assign E13ov6 = (L13ov6 & S13ov6);
assign S13ov6 = (Z13ov6 & G23ov6);
assign L13ov6 = (N23ov6 & U23ov6);
assign X03ov6 = (B33ov6 & I33ov6);
assign I33ov6 = (P33ov6 & W33ov6);
assign B33ov6 = (Fennv6 & D43ov6);
assign En2ov6 = (~(K43ov6 & R43ov6));
assign R43ov6 = (Y43ov6 & F53ov6);
assign F53ov6 = (M53ov6 & T53ov6);
assign T53ov6 = (A63ov6 & H63ov6);
assign H63ov6 = (~(O63ov6 & V63ov6));
assign V63ov6 = (C73ov6 | J73ov6);
assign A63ov6 = (~(Q73ov6 & X73ov6));
assign X73ov6 = (~(E83ov6 & L83ov6));
assign L83ov6 = (S83ov6 & Z83ov6);
assign Z83ov6 = (G93ov6 & N93ov6);
assign N93ov6 = (U93ov6 & Ba3ov6);
assign G93ov6 = (~(Ia3ov6 | Pa3ov6));
assign S83ov6 = (~(Wa3ov6 | Db3ov6));
assign Wa3ov6 = (Kb3ov6 | Rb3ov6);
assign E83ov6 = (Yb3ov6 & Fc3ov6);
assign Fc3ov6 = (Mc3ov6 & Tc3ov6);
assign Tc3ov6 = (~(Ad3ov6 | Hd3ov6));
assign Mc3ov6 = (~(Od3ov6 | Vd3ov6));
assign Yb3ov6 = (~(Ce3ov6 | Je3ov6));
assign Ce3ov6 = (Qe3ov6 | Xe3ov6);
assign Q73ov6 = (~(Ef3ov6 & Lf3ov6));
assign Ef3ov6 = (Sf3ov6 & Zf3ov6);
assign M53ov6 = (Gg3ov6 & Ng3ov6);
assign Ng3ov6 = (~(O63ov6 & Ug3ov6));
assign O63ov6 = (~(Bh3ov6 & Ih3ov6));
assign Ih3ov6 = (Ph3ov6 & Wh3ov6);
assign Wh3ov6 = (~(Di3ov6 | Ki3ov6));
assign Ph3ov6 = (~(Ri3ov6 | Yi3ov6));
assign Bh3ov6 = (Fj3ov6 & Mj3ov6);
assign Mj3ov6 = (~(Tj3ov6 | Ak3ov6));
assign Fj3ov6 = (~(Hk3ov6 | Ok3ov6));
assign Y43ov6 = (Vk3ov6 & Cl3ov6);
assign Cl3ov6 = (Jl3ov6 & Ry1ov6);
assign Jl3ov6 = (!Ql3ov6);
assign Vk3ov6 = (~(Xl3ov6 | Em3ov6));
assign K43ov6 = (Lm3ov6 & Sm3ov6);
assign Sm3ov6 = (Zm3ov6 & Gn3ov6);
assign Gn3ov6 = (~(Nn3ov6 | Un3ov6));
assign Zm3ov6 = (~(Bo3ov6 | Io3ov6));
assign Lm3ov6 = (Po3ov6 & Wo3ov6);
assign Po3ov6 = (Dp3ov6 & Kp3ov6);
assign Qm2ov6 = (Rp3ov6 & Yp3ov6);
assign Yp3ov6 = (~(Fq3ov6 & Mq3ov6));
assign Mq3ov6 = (Tq3ov6 & Ar3ov6);
assign Ar3ov6 = (Hr3ov6 & Or3ov6);
assign Or3ov6 = (Vr3ov6 & Cs3ov6);
assign Cs3ov6 = (~(Js3ov6 | Qs3ov6));
assign Js3ov6 = (Xs3ov6 | Et3ov6);
assign Vr3ov6 = (~(Lt3ov6 | St3ov6));
assign Hr3ov6 = (Zt3ov6 & Gu3ov6);
assign Gu3ov6 = (~(Nu3ov6 | Uu3ov6));
assign Zt3ov6 = (~(Bv3ov6 | Iv3ov6));
assign Tq3ov6 = (Pv3ov6 & Wv3ov6);
assign Wv3ov6 = (Dw3ov6 & Kw3ov6);
assign Kw3ov6 = (~(Rw3ov6 | Wx1ov6));
assign Dw3ov6 = (Yw3ov6 & Fx3ov6);
assign Pv3ov6 = (Mx3ov6 & Tx3ov6);
assign Tx3ov6 = (Ay3ov6 & Hy3ov6);
assign Mx3ov6 = (Oy3ov6 & Vy3ov6);
assign Fq3ov6 = (Cz3ov6 & Jz3ov6);
assign Jz3ov6 = (Qz3ov6 & Xz3ov6);
assign Xz3ov6 = (E04ov6 & L04ov6);
assign L04ov6 = (S04ov6 & Z04ov6);
assign E04ov6 = (G14ov6 & N14ov6);
assign Qz3ov6 = (U14ov6 & B24ov6);
assign B24ov6 = (I24ov6 & P24ov6);
assign U14ov6 = (W24ov6 & D34ov6);
assign Cz3ov6 = (K34ov6 & R34ov6);
assign R34ov6 = (Y34ov6 & F44ov6);
assign F44ov6 = (M44ov6 & T44ov6);
assign Y34ov6 = (A54ov6 & H54ov6);
assign K34ov6 = (O54ov6 & V54ov6);
assign V54ov6 = (C64ov6 & J64ov6);
assign O54ov6 = (Q64ov6 & X64ov6);
assign Rp3ov6 = (~(Px1ov6 & Fhc7z6[30]));
assign Ol2ov6 = (E74ov6 & L74ov6);
assign L74ov6 = (S74ov6 & Z74ov6);
assign Z74ov6 = (G84ov6 & N84ov6);
assign N84ov6 = (U84ov6 & B94ov6);
assign B94ov6 = (~(I94ov6 | Sxkdt6));
assign I94ov6 = (Pvkdt6 | Mtkdt6);
assign U84ov6 = (~(Y1ldt6 | Vzkdt6));
assign G84ov6 = (P94ov6 & W94ov6);
assign W94ov6 = (~(E6ldt6 | B4ldt6));
assign P94ov6 = (~(Kaldt6 | H8ldt6));
assign S74ov6 = (Da4ov6 & Ka4ov6);
assign Ka4ov6 = (Ra4ov6 & Ya4ov6);
assign Ya4ov6 = (~(Qeldt6 | Ncldt6));
assign Ra4ov6 = (~(Wildt6 | Tgldt6));
assign Da4ov6 = (Fb4ov6 & Mb4ov6);
assign Mb4ov6 = (~(Cnldt6 | Zkldt6));
assign Fb4ov6 = (~(Irldt6 | Fpldt6));
assign E74ov6 = (Tb4ov6 & Ac4ov6);
assign Ac4ov6 = (Hc4ov6 & Oc4ov6);
assign Oc4ov6 = (Vc4ov6 & Cd4ov6);
assign Cd4ov6 = (~(Ovldt6 | Ltldt6));
assign Vc4ov6 = (~(Uzldt6 | Rxldt6));
assign Hc4ov6 = (Jd4ov6 & Qd4ov6);
assign Qd4ov6 = (~(A4mdt6 | X1mdt6));
assign Jd4ov6 = (~(G8mdt6 | D6mdt6));
assign Tb4ov6 = (Xd4ov6 & Ee4ov6);
assign Ee4ov6 = (Le4ov6 & Se4ov6);
assign Se4ov6 = (~(Mcmdt6 | Jamdt6));
assign Le4ov6 = (~(Sgmdt6 | Pemdt6));
assign Xd4ov6 = (Ze4ov6 & Gf4ov6);
assign Gf4ov6 = (~(Ykmdt6 | Vimdt6));
assign Ze4ov6 = (~(Nf4ov6 | Bnmdt6));
assign Ev1ov6 = (!Ihinv6);
assign Ihinv6 = (~(Uf4ov6 & Bg4ov6));
assign Al2ov6 = (~(D6gdt6 & Yy1ov6));
assign Yy1ov6 = (~(Ig4ov6 & Pg4ov6));
assign Pg4ov6 = (Wg4ov6 | Bg4ov6);
assign Xel8v6 = (~(Dh4ov6 & Kh4ov6));
assign Kh4ov6 = (Rh4ov6 & Yh4ov6);
assign Yh4ov6 = (~(Td2ov6 & Fi4ov6));
assign Rh4ov6 = (Mi4ov6 & Ti4ov6);
assign Ti4ov6 = (C12ov6 | Sljnv6);
assign Sljnv6 = (Aj4ov6 & Hj4ov6);
assign Hj4ov6 = (Oj4ov6 & Vj4ov6);
assign Vj4ov6 = (Ck4ov6 & Jk4ov6);
assign Jk4ov6 = (Qk4ov6 & Xk4ov6);
assign Xk4ov6 = (~(vis_psp_o[30] & N32ov6));
assign Qk4ov6 = (~(U32ov6 & Pic7z6[30]));
assign Ck4ov6 = (El4ov6 & Ll4ov6);
assign Ll4ov6 = (~(vis_msp_o[30] & P42ov6));
assign El4ov6 = (~(vis_r12_o[30] & W42ov6));
assign Oj4ov6 = (Sl4ov6 & Zl4ov6);
assign Zl4ov6 = (Gm4ov6 & Nm4ov6);
assign Nm4ov6 = (~(vis_r11_o[30] & F62ov6));
assign Gm4ov6 = (~(vis_r10_o[30] & M62ov6));
assign Sl4ov6 = (Um4ov6 & Bn4ov6);
assign Bn4ov6 = (~(vis_r9_o[30] & H72ov6));
assign Um4ov6 = (~(vis_r8_o[30] & O72ov6));
assign Aj4ov6 = (In4ov6 & Pn4ov6);
assign Pn4ov6 = (Wn4ov6 & Do4ov6);
assign Do4ov6 = (Ko4ov6 & Ro4ov6);
assign Ro4ov6 = (~(vis_r7_o[30] & L92ov6));
assign Ko4ov6 = (~(vis_r6_o[30] & S92ov6));
assign Wn4ov6 = (Yo4ov6 & Fp4ov6);
assign Fp4ov6 = (~(vis_r5_o[30] & Na2ov6));
assign Yo4ov6 = (~(vis_r4_o[30] & Ua2ov6));
assign In4ov6 = (Mp4ov6 & Tp4ov6);
assign Tp4ov6 = (Aq4ov6 & Hq4ov6);
assign Hq4ov6 = (~(vis_r3_o[30] & Dc2ov6));
assign Aq4ov6 = (~(vis_r2_o[30] & Kc2ov6));
assign Mp4ov6 = (Oq4ov6 & Vq4ov6);
assign Vq4ov6 = (~(vis_r1_o[30] & Fd2ov6));
assign Oq4ov6 = (~(vis_r0_o[30] & Md2ov6));
assign Mi4ov6 = (~(H02ov6 & Eu97z6));
assign Dh4ov6 = (Cr4ov6 & Jr4ov6);
assign Jr4ov6 = (~(Ve2ov6 & vis_pc_o[30]));
assign Cr4ov6 = (~(Fhc7z6[30] & Cf2ov6));
assign Qel8v6 = (~(Qr4ov6 & Xr4ov6));
assign Qr4ov6 = (Es4ov6 & Ls4ov6);
assign Ls4ov6 = (~(Dpo8v6 & Ss4ov6));
assign Es4ov6 = (~(Oyh7z6[31] & Zs4ov6));
assign Jel8v6 = (~(Gt4ov6 & Nt4ov6));
assign Nt4ov6 = (Ut4ov6 | C397z6);
assign Gt4ov6 = (~(Bu4ov6 & Iu4ov6));
assign Cel8v6 = (~(Pu4ov6 & Wu4ov6));
assign Wu4ov6 = (Dv4ov6 & Kv4ov6);
assign Kv4ov6 = (~(Rv4ov6 & Yv4ov6));
assign Dv4ov6 = (Fw4ov6 & Mw4ov6);
assign Mw4ov6 = (~(Tw4ov6 & Ax4ov6));
assign Fw4ov6 = (~(Hx4ov6 & Ox4ov6));
assign Pu4ov6 = (Vx4ov6 & Cy4ov6);
assign Cy4ov6 = (~(Jy4ov6 & Qy4ov6));
assign Vx4ov6 = (~(Wlr7z6[31] & Xy4ov6));
assign Vdl8v6 = (Lz4ov6 ? K0wmz6[7] : Ez4ov6);
assign Odl8v6 = (~(Sz4ov6 & Zz4ov6));
assign Zz4ov6 = (~(Nsvmz6[7] & G05ov6));
assign Sz4ov6 = (N05ov6 & U05ov6);
assign U05ov6 = (~(Gyvmz6[7] & B15ov6));
assign N05ov6 = (~(I15ov6 & K0wmz6[7]));
assign Hdl8v6 = (W15ov6 ? P15ov6 : V7xmz6[7]);
assign W15ov6 = (!D25ov6);
assign Adl8v6 = (~(K25ov6 & R25ov6));
assign R25ov6 = (~(D25ov6 & La6ft6));
assign Tcl8v6 = (!Y25ov6);
assign Y25ov6 = (T35ov6 ? M35ov6 : F35ov6);
assign Mcl8v6 = (A45ov6 | H45ov6);
assign H45ov6 = (O45ov6 & Fbxmz6[1]);
assign O45ov6 = (Fbxmz6[3] & V45ov6);
assign V45ov6 = (~(C55ov6 & J55ov6));
assign J55ov6 = (~(Q55ov6 & I347v6));
assign Q55ov6 = (~(T35ov6 | O9xmz6[1]));
assign A45ov6 = (T35ov6 ? Fbxmz6[2] : X55ov6);
assign X55ov6 = (~(E65ov6 & L65ov6));
assign L65ov6 = (S65ov6 & Z65ov6);
assign E65ov6 = (G75ov6 & N75ov6);
assign G75ov6 = (~(U75ov6 & B85ov6));
assign Fcl8v6 = (~(I85ov6 & P85ov6));
assign P85ov6 = (~(T35ov6 & Fbxmz6[3]));
assign T35ov6 = (!W85ov6);
assign Ybl8v6 = (W85ov6 ? D95ov6 : Fbxmz6[0]);
assign Rbl8v6 = (~(K95ov6 & R95ov6));
assign R95ov6 = (Y95ov6 | Fa5ov6);
assign K95ov6 = (~(O9xmz6[1] & Ma5ov6));
assign Kbl8v6 = (Ab5ov6 ? Ta5ov6 : Pp1nz6[1]);
assign Ta5ov6 = (~(Hb5ov6 & Ob5ov6));
assign Ob5ov6 = (~(Vb5ov6 & Cc5ov6));
assign Dbl8v6 = (~(Jc5ov6 & Qc5ov6));
assign Qc5ov6 = (~(Xc5ov6 & Ed5ov6));
assign Ed5ov6 = (Hb5ov6 ^ Ld5ov6);
assign Jc5ov6 = (~(U81nz6[0] & Sd5ov6));
assign Wal8v6 = (Ge5ov6 ? Zd5ov6 : Oo1nz6[0]);
assign Pal8v6 = (Ge5ov6 ? Vb5ov6 : Oo1nz6[1]);
assign Ial8v6 = (Ne5ov6 ? Zd5ov6 : Nn1nz6[0]);
assign Bal8v6 = (Ne5ov6 ? Vb5ov6 : Nn1nz6[1]);
assign U9l8v6 = (Ue5ov6 ? Zd5ov6 : Mm1nz6[0]);
assign N9l8v6 = (Ue5ov6 ? Vb5ov6 : Mm1nz6[1]);
assign Vb5ov6 = (~(Bf5ov6 & If5ov6));
assign If5ov6 = (~(V7xmz6[1] & Pf5ov6));
assign Bf5ov6 = (I347v6 ? Dg5ov6 : Wf5ov6);
assign Dg5ov6 = (Kg5ov6 & Rg5ov6);
assign Rg5ov6 = (Yg5ov6 & Fh5ov6);
assign Fh5ov6 = (~(Mh5ov6 & Vcxmz6[22]));
assign Yg5ov6 = (~(Vcxmz6[1] & Gjfnv6));
assign Kg5ov6 = (Th5ov6 & Ai5ov6);
assign Ai5ov6 = (~(Hi5ov6 & Vcxmz6[15]));
assign Th5ov6 = (~(Oi5ov6 & Vcxmz6[8]));
assign Wf5ov6 = (Vi5ov6 & Cj5ov6);
assign Cj5ov6 = (~(Oi5ov6 & Vcxmz6[34]));
assign Vi5ov6 = (Jj5ov6 & Qj5ov6);
assign Qj5ov6 = (~(Gjfnv6 & Vcxmz6[27]));
assign Jj5ov6 = (~(Hi5ov6 & Vcxmz6[41]));
assign G9l8v6 = (~(Xj5ov6 & Ek5ov6));
assign Ek5ov6 = (~(Xc5ov6 & Lk5ov6));
assign Lk5ov6 = (~(Hb5ov6 ^ Sk5ov6));
assign Hb5ov6 = (~(Zk5ov6 & Gl5ov6));
assign Zk5ov6 = (Nl5ov6 ^ Ul5ov6);
assign Xj5ov6 = (~(U81nz6[1] & Sd5ov6));
assign Z8l8v6 = (Im5ov6 ? Bm5ov6 : Md1nz6[0]);
assign Bm5ov6 = (~(Pm5ov6 ^ Wm5ov6));
assign S8l8v6 = (Im5ov6 ? Dn5ov6 : Md1nz6[1]);
assign Dn5ov6 = (Kn5ov6 ^ Pm5ov6);
assign Pm5ov6 = (Rn5ov6 ^ Wm5ov6);
assign L8l8v6 = (Im5ov6 ? Kn5ov6 : Md1nz6[2]);
assign Im5ov6 = (Yn5ov6 & Fo5ov6);
assign Yn5ov6 = (~(Mo5ov6 & To5ov6));
assign To5ov6 = (~(Ap5ov6 & Hp5ov6));
assign Ap5ov6 = (~(Op5ov6 | Vp5ov6));
assign Kn5ov6 = (~(Cq5ov6 ^ Md1nz6[2]));
assign Cq5ov6 = (~(Rn5ov6 & Wm5ov6));
assign Wm5ov6 = (Jq5ov6 | Qq5ov6);
assign E8l8v6 = (Xq5ov6 | Er5ov6);
assign Er5ov6 = (Lr5ov6 & W197z6);
assign Xq5ov6 = (At67v6 ? Zr5ov6 : Sr5ov6);
assign Zr5ov6 = (Gs5ov6 & U42nv6);
assign X7l8v6 = (Ns5ov6 & Us5ov6);
assign Us5ov6 = (Bt5ov6 & It5ov6);
assign It5ov6 = (~(Pt5ov6 & Wt5ov6));
assign Wt5ov6 = (Du5ov6 & Ku5ov6);
assign Ku5ov6 = (~(Ru5ov6 & Ea2ft6));
assign Ru5ov6 = (Cq2ft6 & Yu5ov6);
assign Yu5ov6 = (~(Fv5ov6 & Mv5ov6));
assign Mv5ov6 = (~(Bup7z6[0] & Tv5ov6));
assign Fv5ov6 = (~(Wrp7z6[0] & Aw5ov6));
assign Du5ov6 = (~(Y52ft6 & Hw5ov6));
assign Pt5ov6 = (Ow5ov6 & Vw5ov6);
assign Vw5ov6 = (~(Hc2ft6 & Cx5ov6));
assign Ow5ov6 = (~(B82ft6 & Jx5ov6));
assign Bt5ov6 = (~(Qx5ov6 & Xx5ov6));
assign Xx5ov6 = (~(Ey5ov6 & Ly5ov6));
assign Ly5ov6 = (Gwp7z6[0] ? Zy5ov6 : Sy5ov6);
assign Zy5ov6 = (~(Gz5ov6 & Nz5ov6));
assign Nz5ov6 = (~(Uz5ov6 & B06ov6));
assign B06ov6 = (I06ov6 & P06ov6);
assign P06ov6 = (W06ov6 & D16ov6);
assign D16ov6 = (K16ov6 & R16ov6);
assign W06ov6 = (Y16ov6 & F26ov6);
assign I06ov6 = (M26ov6 & T26ov6);
assign T26ov6 = (~(B2q7z6[9] ^ A36ov6));
assign M26ov6 = (H36ov6 & O36ov6);
assign O36ov6 = (~(B2q7z6[13] ^ V36ov6));
assign H36ov6 = (~(B2q7z6[11] ^ C46ov6));
assign Uz5ov6 = (J46ov6 & Q46ov6);
assign Q46ov6 = (X46ov6 & E56ov6);
assign E56ov6 = (L56ov6 & S56ov6);
assign S56ov6 = (Z56ov6 ^ G66ov6);
assign L56ov6 = (N66ov6 ^ U66ov6);
assign X46ov6 = (B76ov6 & I76ov6);
assign I76ov6 = (~(B2q7z6[8] ^ P76ov6));
assign B76ov6 = (~(B2q7z6[14] ^ W76ov6));
assign J46ov6 = (D86ov6 & K86ov6);
assign D86ov6 = (R86ov6 & Y86ov6);
assign Y86ov6 = (~(B2q7z6[12] ^ F96ov6));
assign Gz5ov6 = (~(M96ov6 & T96ov6));
assign T96ov6 = (Aa6ov6 & Ha6ov6);
assign Ha6ov6 = (Oa6ov6 & Va6ov6);
assign Va6ov6 = (~(B2q7z6[9] ^ Cb6ov6));
assign Aa6ov6 = (Jb6ov6 & Qb6ov6);
assign Qb6ov6 = (~(B2q7z6[10] ^ Xb6ov6));
assign Jb6ov6 = (Ec6ov6 & Lc6ov6);
assign Lc6ov6 = (~(B2q7z6[13] ^ Sc6ov6));
assign Ec6ov6 = (~(B2q7z6[11] ^ Zc6ov6));
assign M96ov6 = (Gd6ov6 & Nd6ov6);
assign Nd6ov6 = (Ud6ov6 & Be6ov6);
assign Be6ov6 = (~(B2q7z6[14] ^ Ie6ov6));
assign Ud6ov6 = (Pe6ov6 & We6ov6);
assign We6ov6 = (~(B2q7z6[15] ^ Df6ov6));
assign Pe6ov6 = (~(B2q7z6[12] ^ Kf6ov6));
assign Gd6ov6 = (Rf6ov6 & Yf6ov6);
assign Rf6ov6 = (Fg6ov6 & Mg6ov6);
assign Mg6ov6 = (~(B2q7z6[8] ^ Tg6ov6));
assign Sy5ov6 = (~(Ah6ov6 & Hh6ov6));
assign Hh6ov6 = (~(Oh6ov6 & Vh6ov6));
assign Vh6ov6 = (Ci6ov6 & Ji6ov6);
assign Ji6ov6 = (Qi6ov6 & Xi6ov6);
assign Xi6ov6 = (Ej6ov6 ^ Sc6ov6);
assign Qi6ov6 = (~(B2q7z6[3] ^ Zc6ov6));
assign Ci6ov6 = (Lj6ov6 & Sj6ov6);
assign Sj6ov6 = (Zj6ov6 ^ Df6ov6);
assign Lj6ov6 = (Gk6ov6 ^ Xb6ov6);
assign Oh6ov6 = (Nk6ov6 & Uk6ov6);
assign Uk6ov6 = (Bl6ov6 & Il6ov6);
assign Il6ov6 = (Pl6ov6 ^ Ie6ov6);
assign Bl6ov6 = (~(B2q7z6[4] ^ Kf6ov6));
assign Nk6ov6 = (Wl6ov6 & Dm6ov6);
assign Dm6ov6 = (~(B2q7z6[0] ^ Tg6ov6));
assign Wl6ov6 = (~(B2q7z6[1] ^ Cb6ov6));
assign Ah6ov6 = (~(Km6ov6 & Oa6ov6));
assign Oa6ov6 = (Rm6ov6 & Ym6ov6);
assign Ym6ov6 = (~(G66ov6 ^ B2q7z6[7]));
assign Rm6ov6 = (~(U66ov6 ^ B2q7z6[2]));
assign Km6ov6 = (Yf6ov6 & Fg6ov6);
assign Fg6ov6 = (Fn6ov6 & Mn6ov6);
assign Mn6ov6 = (Tn6ov6 & Ao6ov6);
assign Ao6ov6 = (Ej6ov6 ^ V36ov6);
assign Tn6ov6 = (~(B2q7z6[3] ^ C46ov6));
assign Fn6ov6 = (Ho6ov6 & Oo6ov6);
assign Oo6ov6 = (Pl6ov6 ^ W76ov6);
assign Ho6ov6 = (~(B2q7z6[4] ^ F96ov6));
assign Yf6ov6 = (Vo6ov6 & Cp6ov6);
assign Cp6ov6 = (~(B2q7z6[0] ^ P76ov6));
assign Vo6ov6 = (~(B2q7z6[1] ^ A36ov6));
assign Ey5ov6 = (Jp6ov6 & Bbp7z6[1]);
assign Qx5ov6 = (Qp6ov6 & Xp6ov6);
assign Xp6ov6 = (~(Eq6ov6 & Lq6ov6));
assign Lq6ov6 = (Sq6ov6 & Zq6ov6);
assign Sq6ov6 = (Gr6ov6 & Nr6ov6);
assign Nr6ov6 = (~(Ur6ov6 & Bs6ov6));
assign Bs6ov6 = (~(Is6ov6 & Ps6ov6));
assign Ps6ov6 = (Ws6ov6 & Dt6ov6);
assign Dt6ov6 = (Kt6ov6 & Rt6ov6);
assign Rt6ov6 = (Yt6ov6 & Fu6ov6);
assign Fu6ov6 = (~(B2q7z6[31] ^ Df6ov6));
assign Df6ov6 = (~(Mu6ov6 & Tu6ov6));
assign Tu6ov6 = (Av6ov6 & Hv6ov6);
assign Hv6ov6 = (~(Ov6ov6 & Ox4ov6));
assign Av6ov6 = (~(Vv6ov6 & Yv4ov6));
assign Mu6ov6 = (Cw6ov6 & Jw6ov6);
assign Jw6ov6 = (~(Qw6ov6 & Ax4ov6));
assign Cw6ov6 = (~(Xw6ov6 & Qy4ov6));
assign Yt6ov6 = (~(Ex6ov6 | Lx6ov6));
assign Kt6ov6 = (Sx6ov6 & Zx6ov6);
assign Zx6ov6 = (~(B2q7z6[26] ^ Xb6ov6));
assign Xb6ov6 = (~(Gy6ov6 & Ny6ov6));
assign Ny6ov6 = (Uy6ov6 & Bz6ov6);
assign Bz6ov6 = (~(Ov6ov6 & Iz6ov6));
assign Uy6ov6 = (~(Vv6ov6 & Pz6ov6));
assign Gy6ov6 = (Wz6ov6 & D07ov6);
assign D07ov6 = (~(Qw6ov6 & K07ov6));
assign Wz6ov6 = (~(Xw6ov6 & R07ov6));
assign Sx6ov6 = (~(B2q7z6[24] ^ Tg6ov6));
assign Tg6ov6 = (~(Y07ov6 & F17ov6));
assign F17ov6 = (M17ov6 & T17ov6);
assign T17ov6 = (~(Ov6ov6 & A27ov6));
assign M17ov6 = (~(Vv6ov6 & H27ov6));
assign Y07ov6 = (O27ov6 & V27ov6);
assign V27ov6 = (~(Qw6ov6 & C37ov6));
assign O27ov6 = (~(Xw6ov6 & J37ov6));
assign Ws6ov6 = (Q37ov6 & X37ov6);
assign X37ov6 = (E47ov6 & L47ov6);
assign L47ov6 = (~(B2q7z6[28] ^ Kf6ov6));
assign Kf6ov6 = (~(S47ov6 & Z47ov6));
assign Z47ov6 = (G57ov6 & N57ov6);
assign N57ov6 = (~(Ov6ov6 & U57ov6));
assign G57ov6 = (~(Vv6ov6 & B67ov6));
assign S47ov6 = (I67ov6 & P67ov6);
assign P67ov6 = (~(Qw6ov6 & W67ov6));
assign I67ov6 = (~(Xw6ov6 & D77ov6));
assign E47ov6 = (K77ov6 & R77ov6);
assign R77ov6 = (~(B2q7z6[25] ^ Cb6ov6));
assign Cb6ov6 = (~(Y77ov6 & F87ov6));
assign F87ov6 = (M87ov6 & T87ov6);
assign T87ov6 = (~(Ov6ov6 & A97ov6));
assign M87ov6 = (~(Vv6ov6 & H97ov6));
assign Y77ov6 = (O97ov6 & V97ov6);
assign V97ov6 = (~(Qw6ov6 & Ca7ov6));
assign O97ov6 = (~(Xw6ov6 & Ja7ov6));
assign K77ov6 = (~(B2q7z6[27] ^ Zc6ov6));
assign Zc6ov6 = (~(Qa7ov6 & Xa7ov6));
assign Xa7ov6 = (Eb7ov6 & Lb7ov6);
assign Lb7ov6 = (~(Ov6ov6 & Sb7ov6));
assign Eb7ov6 = (~(Vv6ov6 & Zb7ov6));
assign Qa7ov6 = (Gc7ov6 & Nc7ov6);
assign Nc7ov6 = (~(Qw6ov6 & Uc7ov6));
assign Gc7ov6 = (~(Xw6ov6 & Bd7ov6));
assign Q37ov6 = (Id7ov6 & Pd7ov6);
assign Pd7ov6 = (~(B2q7z6[23] ^ G66ov6));
assign G66ov6 = (~(Wd7ov6 & De7ov6));
assign De7ov6 = (Ke7ov6 & Re7ov6);
assign Re7ov6 = (~(Ov6ov6 & Yv4ov6));
assign Ke7ov6 = (~(Vv6ov6 & Ax4ov6));
assign Wd7ov6 = (Ye7ov6 & Ff7ov6);
assign Ff7ov6 = (~(Qw6ov6 & Qy4ov6));
assign Ye7ov6 = (~(Xw6ov6 & Ox4ov6));
assign Id7ov6 = (~(B2q7z6[29] ^ Sc6ov6));
assign Sc6ov6 = (~(Mf7ov6 & Tf7ov6));
assign Tf7ov6 = (Ag7ov6 & Hg7ov6);
assign Hg7ov6 = (~(Ov6ov6 & Og7ov6));
assign Ag7ov6 = (~(Vv6ov6 & Vg7ov6));
assign Mf7ov6 = (Ch7ov6 & Jh7ov6);
assign Jh7ov6 = (~(Qw6ov6 & Qh7ov6));
assign Ch7ov6 = (~(Xw6ov6 & Xh7ov6));
assign Is6ov6 = (Ei7ov6 & Li7ov6);
assign Li7ov6 = (Si7ov6 & Zi7ov6);
assign Zi7ov6 = (Gj7ov6 & Nj7ov6);
assign Nj7ov6 = (~(B2q7z6[17] ^ A36ov6));
assign A36ov6 = (~(Uj7ov6 & Bk7ov6));
assign Bk7ov6 = (Ik7ov6 & Pk7ov6);
assign Pk7ov6 = (~(Ov6ov6 & H97ov6));
assign Ik7ov6 = (~(Vv6ov6 & Ca7ov6));
assign Uj7ov6 = (Wk7ov6 & Dl7ov6);
assign Dl7ov6 = (~(Qw6ov6 & Ja7ov6));
assign Wk7ov6 = (~(Xw6ov6 & A97ov6));
assign Gj7ov6 = (Kl7ov6 & Rl7ov6);
assign Rl7ov6 = (~(B2q7z6[30] ^ Ie6ov6));
assign Ie6ov6 = (~(Yl7ov6 & Fm7ov6));
assign Fm7ov6 = (Mm7ov6 & Tm7ov6);
assign Tm7ov6 = (~(Ov6ov6 & An7ov6));
assign Mm7ov6 = (~(Vv6ov6 & Hn7ov6));
assign Yl7ov6 = (On7ov6 & Vn7ov6);
assign Vn7ov6 = (~(Qw6ov6 & Co7ov6));
assign On7ov6 = (~(Xw6ov6 & Jo7ov6));
assign Kl7ov6 = (~(B2q7z6[16] ^ P76ov6));
assign P76ov6 = (~(Qo7ov6 & Xo7ov6));
assign Xo7ov6 = (Ep7ov6 & Lp7ov6);
assign Lp7ov6 = (~(Ov6ov6 & H27ov6));
assign Ep7ov6 = (~(Vv6ov6 & C37ov6));
assign Qo7ov6 = (Sp7ov6 & Zp7ov6);
assign Zp7ov6 = (~(Qw6ov6 & J37ov6));
assign Sp7ov6 = (~(Xw6ov6 & A27ov6));
assign Si7ov6 = (Gq7ov6 & Nq7ov6);
assign Nq7ov6 = (~(B2q7z6[20] ^ F96ov6));
assign F96ov6 = (~(Uq7ov6 & Br7ov6));
assign Br7ov6 = (Ir7ov6 & Pr7ov6);
assign Pr7ov6 = (~(Ov6ov6 & B67ov6));
assign Ir7ov6 = (~(Vv6ov6 & W67ov6));
assign Uq7ov6 = (Wr7ov6 & Ds7ov6);
assign Ds7ov6 = (~(Qw6ov6 & D77ov6));
assign Wr7ov6 = (~(Xw6ov6 & U57ov6));
assign Gq7ov6 = (~(B2q7z6[18] ^ U66ov6));
assign U66ov6 = (~(Ks7ov6 & Rs7ov6));
assign Rs7ov6 = (Ys7ov6 & Ft7ov6);
assign Ft7ov6 = (~(Ov6ov6 & Pz6ov6));
assign Ys7ov6 = (~(Vv6ov6 & K07ov6));
assign Ks7ov6 = (Mt7ov6 & Tt7ov6);
assign Tt7ov6 = (~(Qw6ov6 & R07ov6));
assign Mt7ov6 = (~(Xw6ov6 & Iz6ov6));
assign Ei7ov6 = (Au7ov6 & Hu7ov6);
assign Hu7ov6 = (Ou7ov6 & Vu7ov6);
assign Vu7ov6 = (~(B2q7z6[22] ^ W76ov6));
assign W76ov6 = (~(Cv7ov6 & Jv7ov6));
assign Jv7ov6 = (Qv7ov6 & Xv7ov6);
assign Xv7ov6 = (~(Ov6ov6 & Hn7ov6));
assign Qv7ov6 = (~(Vv6ov6 & Co7ov6));
assign Cv7ov6 = (Ew7ov6 & Lw7ov6);
assign Lw7ov6 = (~(Qw6ov6 & Jo7ov6));
assign Ew7ov6 = (~(Xw6ov6 & An7ov6));
assign Ou7ov6 = (Sw7ov6 & Zw7ov6);
assign Zw7ov6 = (~(B2q7z6[19] ^ C46ov6));
assign C46ov6 = (~(Gx7ov6 & Nx7ov6));
assign Nx7ov6 = (Ux7ov6 & By7ov6);
assign By7ov6 = (~(Ov6ov6 & Zb7ov6));
assign Ux7ov6 = (~(Vv6ov6 & Uc7ov6));
assign Gx7ov6 = (Iy7ov6 & Py7ov6);
assign Py7ov6 = (~(Qw6ov6 & Bd7ov6));
assign Iy7ov6 = (~(Xw6ov6 & Sb7ov6));
assign Sw7ov6 = (~(B2q7z6[21] ^ V36ov6));
assign V36ov6 = (~(Wy7ov6 & Dz7ov6));
assign Dz7ov6 = (Kz7ov6 & Rz7ov6);
assign Rz7ov6 = (~(Ov6ov6 & Vg7ov6));
assign Kz7ov6 = (~(Vv6ov6 & Qh7ov6));
assign Wy7ov6 = (Yz7ov6 & F08ov6);
assign F08ov6 = (~(Qw6ov6 & Xh7ov6));
assign Yz7ov6 = (~(Xw6ov6 & Og7ov6));
assign Au7ov6 = (M08ov6 & Gwp7z6[1]);
assign Ur6ov6 = (~(Jp6ov6 & T08ov6));
assign Qp6ov6 = (~(A18ov6 & Jp6ov6));
assign Jp6ov6 = (~(H18ov6 | Ex6ov6));
assign Ex6ov6 = (L42ft6 ? V18ov6 : O18ov6);
assign H18ov6 = (Lx6ov6 | Gwp7z6[1]);
assign A18ov6 = (C28ov6 & J28ov6);
assign J28ov6 = (~(Q28ov6 & X28ov6));
assign X28ov6 = (~(E38ov6 & L38ov6));
assign L38ov6 = (S38ov6 & Z38ov6);
assign Z38ov6 = (R16ov6 & T08ov6);
assign R16ov6 = (~(G48ov6 ^ B2q7z6[5]));
assign S38ov6 = (F26ov6 & K16ov6);
assign K16ov6 = (~(N48ov6 ^ B2q7z6[7]));
assign F26ov6 = (~(U48ov6 ^ B2q7z6[2]));
assign E38ov6 = (B58ov6 & K86ov6);
assign K86ov6 = (I58ov6 & P58ov6);
assign P58ov6 = (~(B2q7z6[3] ^ W58ov6));
assign I58ov6 = (~(B2q7z6[4] ^ D68ov6));
assign B58ov6 = (R86ov6 & Y16ov6);
assign Y16ov6 = (~(K68ov6 ^ B2q7z6[6]));
assign R86ov6 = (R68ov6 & Y68ov6);
assign Y68ov6 = (~(B2q7z6[0] ^ F78ov6));
assign R68ov6 = (~(B2q7z6[1] ^ M78ov6));
assign Q28ov6 = (~(Eq6ov6 & T78ov6));
assign T78ov6 = (A88ov6 & M08ov6);
assign M08ov6 = (H88ov6 & O88ov6);
assign O88ov6 = (V88ov6 & C98ov6);
assign C98ov6 = (J98ov6 & Q98ov6);
assign Q98ov6 = (~(B2q7z6[13] ^ G48ov6));
assign G48ov6 = (~(X98ov6 & Ea8ov6));
assign Ea8ov6 = (La8ov6 & Sa8ov6);
assign Sa8ov6 = (~(Ov6ov6 & Qh7ov6));
assign La8ov6 = (~(Vv6ov6 & Xh7ov6));
assign X98ov6 = (Za8ov6 & Gb8ov6);
assign Gb8ov6 = (~(Qw6ov6 & Og7ov6));
assign Za8ov6 = (~(Xw6ov6 & Vg7ov6));
assign J98ov6 = (~(B2q7z6[11] ^ W58ov6));
assign W58ov6 = (~(Nb8ov6 & Ub8ov6));
assign Ub8ov6 = (Bc8ov6 & Ic8ov6);
assign Ic8ov6 = (~(Ov6ov6 & Uc7ov6));
assign Bc8ov6 = (~(Vv6ov6 & Bd7ov6));
assign Nb8ov6 = (Pc8ov6 & Wc8ov6);
assign Wc8ov6 = (~(Qw6ov6 & Sb7ov6));
assign Pc8ov6 = (~(Xw6ov6 & Zb7ov6));
assign V88ov6 = (Dd8ov6 & Kd8ov6);
assign Kd8ov6 = (Z56ov6 ^ N48ov6);
assign N48ov6 = (~(Rd8ov6 & Yd8ov6));
assign Yd8ov6 = (Fe8ov6 & Me8ov6);
assign Me8ov6 = (~(Ov6ov6 & Ax4ov6));
assign Fe8ov6 = (~(Vv6ov6 & Qy4ov6));
assign Rd8ov6 = (Te8ov6 & Af8ov6);
assign Af8ov6 = (~(Qw6ov6 & Ox4ov6));
assign Te8ov6 = (~(Xw6ov6 & Yv4ov6));
assign Z56ov6 = (!B2q7z6[15]);
assign Dd8ov6 = (N66ov6 ^ U48ov6);
assign U48ov6 = (~(Hf8ov6 & Of8ov6));
assign Of8ov6 = (Vf8ov6 & Cg8ov6);
assign Cg8ov6 = (~(Ov6ov6 & K07ov6));
assign Vf8ov6 = (~(Vv6ov6 & R07ov6));
assign Hf8ov6 = (Jg8ov6 & Qg8ov6);
assign Qg8ov6 = (~(Qw6ov6 & Iz6ov6));
assign Jg8ov6 = (~(Xw6ov6 & Pz6ov6));
assign N66ov6 = (!B2q7z6[10]);
assign H88ov6 = (Xg8ov6 & Eh8ov6);
assign Eh8ov6 = (Lh8ov6 & Sh8ov6);
assign Sh8ov6 = (~(B2q7z6[14] ^ K68ov6));
assign K68ov6 = (~(Zh8ov6 & Gi8ov6));
assign Gi8ov6 = (Ni8ov6 & Ui8ov6);
assign Ui8ov6 = (~(Ov6ov6 & Co7ov6));
assign Ni8ov6 = (~(Vv6ov6 & Jo7ov6));
assign Zh8ov6 = (Bj8ov6 & Ij8ov6);
assign Ij8ov6 = (~(Qw6ov6 & An7ov6));
assign Bj8ov6 = (~(Xw6ov6 & Hn7ov6));
assign Lh8ov6 = (~(B2q7z6[12] ^ D68ov6));
assign D68ov6 = (~(Pj8ov6 & Wj8ov6));
assign Wj8ov6 = (Dk8ov6 & Kk8ov6);
assign Kk8ov6 = (~(Ov6ov6 & W67ov6));
assign Dk8ov6 = (~(Vv6ov6 & D77ov6));
assign Pj8ov6 = (Rk8ov6 & Yk8ov6);
assign Yk8ov6 = (~(Qw6ov6 & U57ov6));
assign Rk8ov6 = (~(Xw6ov6 & B67ov6));
assign Xg8ov6 = (Fl8ov6 & Ml8ov6);
assign Ml8ov6 = (Tl8ov6 ^ F78ov6);
assign F78ov6 = (~(Am8ov6 & Hm8ov6));
assign Hm8ov6 = (Om8ov6 & Vm8ov6);
assign Vm8ov6 = (~(Ov6ov6 & C37ov6));
assign Om8ov6 = (~(Vv6ov6 & J37ov6));
assign Am8ov6 = (Cn8ov6 & Jn8ov6);
assign Jn8ov6 = (~(Qw6ov6 & A27ov6));
assign Cn8ov6 = (~(Xw6ov6 & H27ov6));
assign Tl8ov6 = (!B2q7z6[8]);
assign Fl8ov6 = (~(B2q7z6[9] ^ M78ov6));
assign M78ov6 = (~(Qn8ov6 & Xn8ov6));
assign Xn8ov6 = (Eo8ov6 & Lo8ov6);
assign Lo8ov6 = (~(Ov6ov6 & Ca7ov6));
assign Eo8ov6 = (~(Vv6ov6 & Ja7ov6));
assign Qn8ov6 = (So8ov6 & Zo8ov6);
assign Zo8ov6 = (~(Qw6ov6 & A97ov6));
assign So8ov6 = (~(Xw6ov6 & H97ov6));
assign A88ov6 = (Zq6ov6 & Gr6ov6);
assign Gr6ov6 = (Gp8ov6 ^ Pl6ov6);
assign Pl6ov6 = (!B2q7z6[6]);
assign Gp8ov6 = (~(Np8ov6 & Up8ov6));
assign Up8ov6 = (Bq8ov6 & Iq8ov6);
assign Iq8ov6 = (~(Ov6ov6 & Jo7ov6));
assign Bq8ov6 = (~(Vv6ov6 & An7ov6));
assign Np8ov6 = (Pq8ov6 & Wq8ov6);
assign Wq8ov6 = (~(Qw6ov6 & Hn7ov6));
assign Pq8ov6 = (~(Xw6ov6 & Co7ov6));
assign Zq6ov6 = (Dr8ov6 ^ Ej6ov6);
assign Ej6ov6 = (!B2q7z6[5]);
assign Dr8ov6 = (~(Kr8ov6 & Rr8ov6));
assign Rr8ov6 = (Yr8ov6 & Fs8ov6);
assign Fs8ov6 = (~(Ov6ov6 & Xh7ov6));
assign Yr8ov6 = (~(Vv6ov6 & Og7ov6));
assign Kr8ov6 = (Ms8ov6 & Ts8ov6);
assign Ts8ov6 = (~(Qw6ov6 & Vg7ov6));
assign Ms8ov6 = (~(Xw6ov6 & Qh7ov6));
assign Eq6ov6 = (~(At8ov6 | Ht8ov6));
assign Ht8ov6 = (~(Ot8ov6 & Vt8ov6));
assign Vt8ov6 = (Cu8ov6 & Ju8ov6);
assign Ju8ov6 = (~(Zj6ov6 ^ Qu8ov6));
assign Qu8ov6 = (Xu8ov6 & Ev8ov6);
assign Ev8ov6 = (Lv8ov6 & Sv8ov6);
assign Sv8ov6 = (~(Ov6ov6 & Qy4ov6));
assign Lv8ov6 = (~(Vv6ov6 & Ox4ov6));
assign Xu8ov6 = (Zv8ov6 & Gw8ov6);
assign Gw8ov6 = (~(Qw6ov6 & Yv4ov6));
assign Zv8ov6 = (~(Xw6ov6 & Ax4ov6));
assign Zj6ov6 = (!B2q7z6[7]);
assign Cu8ov6 = (~(Gk6ov6 ^ Nw8ov6));
assign Nw8ov6 = (Uw8ov6 & Bx8ov6);
assign Bx8ov6 = (Ix8ov6 & Px8ov6);
assign Px8ov6 = (~(Ov6ov6 & R07ov6));
assign Ix8ov6 = (~(Vv6ov6 & Iz6ov6));
assign Uw8ov6 = (Wx8ov6 & Dy8ov6);
assign Dy8ov6 = (~(Qw6ov6 & Pz6ov6));
assign Wx8ov6 = (~(Xw6ov6 & K07ov6));
assign Gk6ov6 = (!B2q7z6[2]);
assign Ot8ov6 = (Ky8ov6 & Ry8ov6);
assign Ry8ov6 = (B2q7z6[0] ^ Yy8ov6);
assign Yy8ov6 = (Fz8ov6 & Mz8ov6);
assign Mz8ov6 = (Tz8ov6 & A09ov6);
assign A09ov6 = (~(Ov6ov6 & J37ov6));
assign Tz8ov6 = (~(Vv6ov6 & A27ov6));
assign Fz8ov6 = (H09ov6 & O09ov6);
assign O09ov6 = (~(Qw6ov6 & H27ov6));
assign H09ov6 = (~(Xw6ov6 & C37ov6));
assign Ky8ov6 = (B2q7z6[1] ^ V09ov6);
assign V09ov6 = (C19ov6 & J19ov6);
assign J19ov6 = (Q19ov6 & X19ov6);
assign X19ov6 = (~(Ov6ov6 & Ja7ov6));
assign Q19ov6 = (~(Vv6ov6 & A97ov6));
assign C19ov6 = (E29ov6 & L29ov6);
assign L29ov6 = (~(Qw6ov6 & H97ov6));
assign E29ov6 = (~(Xw6ov6 & Ca7ov6));
assign At8ov6 = (~(S29ov6 & Z29ov6));
assign Z29ov6 = (B2q7z6[3] ^ G39ov6);
assign G39ov6 = (N39ov6 & U39ov6);
assign U39ov6 = (B49ov6 & I49ov6);
assign I49ov6 = (~(Ov6ov6 & Bd7ov6));
assign B49ov6 = (~(Vv6ov6 & Sb7ov6));
assign N39ov6 = (P49ov6 & W49ov6);
assign W49ov6 = (~(Qw6ov6 & Zb7ov6));
assign P49ov6 = (~(Xw6ov6 & Uc7ov6));
assign S29ov6 = (B2q7z6[4] ^ D59ov6);
assign D59ov6 = (K59ov6 & R59ov6);
assign R59ov6 = (Y59ov6 & F69ov6);
assign F69ov6 = (~(Ov6ov6 & D77ov6));
assign Ov6ov6 = (~(M69ov6 | Ncp7z6[0]));
assign Y59ov6 = (~(Vv6ov6 & U57ov6));
assign Vv6ov6 = (~(T69ov6 | Ncp7z6[1]));
assign K59ov6 = (A79ov6 & H79ov6);
assign H79ov6 = (~(Qw6ov6 & B67ov6));
assign Qw6ov6 = (~(Ncp7z6[0] | Ncp7z6[1]));
assign A79ov6 = (~(Xw6ov6 & W67ov6));
assign Xw6ov6 = (~(T69ov6 | M69ov6));
assign C28ov6 = (Bbp7z6[1] | Bbp7z6[0]);
assign Ns5ov6 = (O5a7z6 & O79ov6);
assign O79ov6 = (~(Gwp7z6[1] & V79ov6));
assign V79ov6 = (~(Bbp7z6[1] & C89ov6));
assign C89ov6 = (T08ov6 | Bbp7z6[0]);
assign T08ov6 = (!Gwp7z6[0]);
assign Q7l8v6 = (~(J89ov6 & Q89ov6));
assign Q89ov6 = (X89ov6 & E99ov6);
assign X89ov6 = (~(L99ov6 | Mb88v6));
assign J89ov6 = (S99ov6 & Z99ov6);
assign Z99ov6 = (~(Gg2ft6 & Ga9ov6));
assign Ga9ov6 = (~(Na9ov6 & Ua9ov6));
assign S99ov6 = (~(Kg5ft6 & Bb9ov6));
assign C7l8v6 = (Pb9ov6 ? D6c7z6[0] : Ib9ov6);
assign Ib9ov6 = (~(Wb9ov6 & Dc9ov6));
assign Dc9ov6 = (Kc9ov6 & Rc9ov6);
assign Rc9ov6 = (~(Yc9ov6 & Fd9ov6));
assign Kc9ov6 = (~(Md9ov6 & Td9ov6));
assign Wb9ov6 = (Ae9ov6 & He9ov6);
assign He9ov6 = (~(Oe9ov6 & Ve9ov6));
assign Ae9ov6 = (~(Cf9ov6 & Jf9ov6));
assign O6l8v6 = (~(Qf9ov6 & Xf9ov6));
assign Xf9ov6 = (Eg9ov6 | Mulnv6);
assign Qf9ov6 = (~(Lg9ov6 & Sg9ov6));
assign Sg9ov6 = (Zg9ov6 & Gh9ov6);
assign Gh9ov6 = (~(Nh9ov6 & Uh9ov6));
assign Uh9ov6 = (Bi9ov6 & Ii9ov6);
assign Nh9ov6 = (Gr2et6 & Pi9ov6);
assign Zg9ov6 = (Xmvnv6 & Dxvnv6);
assign Xmvnv6 = (~(Wi9ov6 & Dj9ov6));
assign Wi9ov6 = (Q0wnv6 & Ldo7v6);
assign Lg9ov6 = (S7xdt6 & Kj9ov6);
assign Kj9ov6 = (~(Ecc7z6[14] & Pbadt6));
assign A6l8v6 = (Yj9ov6 ? Rj9ov6 : Kyn7z6[0]);
assign T5l8v6 = (Yj9ov6 ? Fk9ov6 : Kyn7z6[1]);
assign Yj9ov6 = (!Mk9ov6);
assign M5l8v6 = (~(Tk9ov6 & Al9ov6));
assign Al9ov6 = (~(Hl9ov6 & Ol9ov6));
assign Ol9ov6 = (~(Vl9ov6 & Cm9ov6));
assign Cm9ov6 = (Jm9ov6 & Qm9ov6);
assign Jm9ov6 = (Xm9ov6 & En9ov6);
assign Vl9ov6 = (Ln9ov6 & Sn9ov6);
assign Sn9ov6 = (Zn9ov6 | Go9ov6);
assign Ln9ov6 = (No9ov6 & Uo9ov6);
assign Uo9ov6 = (~(Bp9ov6 & Ip9ov6));
assign Ip9ov6 = (~(Pp9ov6 & Wp9ov6));
assign Tk9ov6 = (~(Dq9ov6 & Qln7z6[1]));
assign F5l8v6 = (~(Kq9ov6 & Rq9ov6));
assign Rq9ov6 = (~(Hl9ov6 & Yq9ov6));
assign Kq9ov6 = (~(Dq9ov6 & Xnnet6));
assign Y4l8v6 = (Rconv6 ? Yk1ov6 : Meoet6);
assign R4l8v6 = (Mr9ov6 ? Hrb7z6[0] : Fr9ov6);
assign K4l8v6 = (As9ov6 ? L9d7z6[2] : Tr9ov6);
assign D4l8v6 = (~(Hs9ov6 & Os9ov6));
assign Os9ov6 = (~(W9edt6 & Vs9ov6));
assign W3l8v6 = (~(Ct9ov6 & Jt9ov6));
assign Jt9ov6 = (Qt9ov6 & Xt9ov6);
assign Xt9ov6 = (Eu9ov6 | Lu9ov6);
assign Qt9ov6 = (Su9ov6 & Zu9ov6);
assign Zu9ov6 = (~(Gv9ov6 & Nv9ov6));
assign Su9ov6 = (~(Uv9ov6 & Mu97z6));
assign Ct9ov6 = (Bw9ov6 & Iw9ov6);
assign Iw9ov6 = (~(Pw9ov6 & Kxb7z6[1]));
assign Bw9ov6 = (Ww9ov6 & Dx9ov6);
assign Dx9ov6 = (~(Kx9ov6 & vis_pc_o[1]));
assign Ww9ov6 = (~(Rx9ov6 & Gli7z6[1]));
assign P3l8v6 = (~(Yx9ov6 & Fy9ov6));
assign Fy9ov6 = (~(My9ov6 & Qu1ov6));
assign Yx9ov6 = (Ty9ov6 & Az9ov6);
assign Az9ov6 = (~(Hz9ov6 & H9gdt6));
assign Ty9ov6 = (~(Uf4ov6 & Pfgdt6));
assign Pfgdt6 = (Vz9ov6 ? Oz9ov6 : H9gdt6);
assign Vz9ov6 = (Uf4ov6 & C0aov6);
assign C0aov6 = (~(J0aov6 & Q0aov6));
assign J0aov6 = (~(Dte7z6[19] & Dte7z6[18]));
assign Oz9ov6 = (!X0aov6);
assign X0aov6 = (Jm2ov6 ? L1aov6 : E1aov6);
assign L1aov6 = (~(S1aov6 & Z1aov6));
assign Z1aov6 = (~(X2g7z6[31] & G2aov6));
assign S1aov6 = (J5g7z6[31] ? X2g7z6[31] : G2aov6);
assign J5g7z6[31] = (N2aov6 & Aumnv6);
assign Aumnv6 = (!Sannv6);
assign Sannv6 = (~(U2aov6 | Dte7z6[2]));
assign X2g7z6[31] = (B3aov6 & Gbnnv6);
assign Gbnnv6 = (!Oumnv6);
assign Oumnv6 = (~(U2aov6 | Dte7z6[3]));
assign U2aov6 = (~(I3aov6 & P3aov6));
assign P3aov6 = (~(W3aov6 & D4aov6));
assign W3aov6 = (~(K4aov6 & R4aov6));
assign I3aov6 = (Y4aov6 & F5aov6);
assign F5aov6 = (!M5aov6);
assign G2aov6 = (T5aov6 | L0g7z6[31]);
assign T5aov6 = (!Ky1ov6);
assign E1aov6 = (~(Px1ov6 & Fhc7z6[28]));
assign I3l8v6 = (~(A6aov6 & H6aov6));
assign H6aov6 = (O6aov6 & V6aov6);
assign V6aov6 = (~(Td2ov6 & C7aov6));
assign O6aov6 = (J7aov6 & Q7aov6);
assign Q7aov6 = (C12ov6 | Oqjnv6);
assign Oqjnv6 = (X7aov6 & E8aov6);
assign E8aov6 = (L8aov6 & S8aov6);
assign S8aov6 = (Z8aov6 & G9aov6);
assign G9aov6 = (N9aov6 & U9aov6);
assign U9aov6 = (~(vis_psp_o[28] & N32ov6));
assign N9aov6 = (~(U32ov6 & Pic7z6[28]));
assign Z8aov6 = (Baaov6 & Iaaov6);
assign Iaaov6 = (~(vis_msp_o[28] & P42ov6));
assign Baaov6 = (~(vis_r12_o[28] & W42ov6));
assign L8aov6 = (Paaov6 & Waaov6);
assign Waaov6 = (Dbaov6 & Kbaov6);
assign Kbaov6 = (~(vis_r11_o[28] & F62ov6));
assign Dbaov6 = (~(vis_r10_o[28] & M62ov6));
assign Paaov6 = (Rbaov6 & Ybaov6);
assign Ybaov6 = (~(vis_r9_o[28] & H72ov6));
assign Rbaov6 = (~(vis_r8_o[28] & O72ov6));
assign X7aov6 = (Fcaov6 & Mcaov6);
assign Mcaov6 = (Tcaov6 & Adaov6);
assign Adaov6 = (Hdaov6 & Odaov6);
assign Odaov6 = (~(vis_r7_o[28] & L92ov6));
assign Hdaov6 = (~(vis_r6_o[28] & S92ov6));
assign Tcaov6 = (Vdaov6 & Ceaov6);
assign Ceaov6 = (~(vis_r5_o[28] & Na2ov6));
assign Vdaov6 = (~(vis_r4_o[28] & Ua2ov6));
assign Fcaov6 = (Jeaov6 & Qeaov6);
assign Qeaov6 = (Xeaov6 & Efaov6);
assign Efaov6 = (~(vis_r3_o[28] & Dc2ov6));
assign Xeaov6 = (~(vis_r2_o[28] & Kc2ov6));
assign Jeaov6 = (Lfaov6 & Sfaov6);
assign Sfaov6 = (~(vis_r1_o[28] & Fd2ov6));
assign Lfaov6 = (~(vis_r0_o[28] & Md2ov6));
assign J7aov6 = (~(H02ov6 & Uu97z6));
assign A6aov6 = (Zfaov6 & Ggaov6);
assign Ggaov6 = (~(Ve2ov6 & vis_pc_o[28]));
assign Zfaov6 = (~(Fhc7z6[28] & Cf2ov6));
assign B3l8v6 = (Ngaov6 & Ugaov6);
assign Ugaov6 = (~(Bhaov6 | Pacdt6));
assign Ngaov6 = (Snvnv6 & Ihaov6);
assign U2l8v6 = (~(Phaov6 & Whaov6));
assign Whaov6 = (Diaov6 | G597z6);
assign N2l8v6 = (~(Ij1ov6 & Kiaov6));
assign Kiaov6 = (~(Riaov6 & Lpc7z6[1]));
assign G2l8v6 = (Diaov6 ? Yiaov6 : Pmc7z6[0]);
assign Z1l8v6 = (Diaov6 ? Fjaov6 : Pmc7z6[1]);
assign S1l8v6 = (~(Mjaov6 & Tjaov6));
assign Tjaov6 = (Akaov6 & Hkaov6);
assign Hkaov6 = (~(Ohe7z6[7] & Okaov6));
assign Akaov6 = (Vkaov6 & Claov6);
assign Claov6 = (~(Jlaov6 & Zec7z6[7]));
assign Vkaov6 = (~(Qlaov6 & Xlaov6));
assign Mjaov6 = (Emaov6 & Lmaov6);
assign Lmaov6 = (Smaov6 | Zmaov6);
assign Emaov6 = (~(Gnaov6 & Zec7z6[23]));
assign L1l8v6 = (~(Unaov6 & Boaov6));
assign Boaov6 = (Ioaov6 & Poaov6);
assign Poaov6 = (~(Ohe7z6[6] & Okaov6));
assign Ioaov6 = (Woaov6 & Dpaov6);
assign Dpaov6 = (~(Jlaov6 & Zec7z6[6]));
assign Woaov6 = (~(Qlaov6 & Kpaov6));
assign Unaov6 = (Rpaov6 & Ypaov6);
assign Ypaov6 = (Smaov6 | Fqaov6);
assign Rpaov6 = (~(Gnaov6 & Zec7z6[22]));
assign E1l8v6 = (!Mqaov6);
assign Mqaov6 = (Nnaov6 ? Qtvnv6 : Tqaov6);
assign Tqaov6 = (Araov6 & Hraov6);
assign Hraov6 = (Oraov6 & Vraov6);
assign Vraov6 = (Csaov6 & Jsaov6);
assign Csaov6 = (Qsaov6 & Srknv6);
assign Oraov6 = (Xsaov6 & Etaov6);
assign Xsaov6 = (~(Ltaov6 & Staov6));
assign Ltaov6 = (Ztaov6 & Guaov6);
assign Guaov6 = (~(Nuaov6 & Uuaov6));
assign Uuaov6 = (Fqaov6 & Zmaov6);
assign Nuaov6 = (Bvaov6 & Ivaov6);
assign Araov6 = (Pvaov6 & Wvaov6);
assign Wvaov6 = (Dwaov6 & Kwaov6);
assign Kwaov6 = (~(Rwaov6 & Yl2et6));
assign Rwaov6 = (Ywaov6 & Fxaov6);
assign Dwaov6 = (~(Xtvnv6 & Mxaov6));
assign Mxaov6 = (~(Txaov6 & Ayaov6));
assign Pvaov6 = (Hyaov6 & Oyaov6);
assign Oyaov6 = (Vyaov6 | Txinv6);
assign Vyaov6 = (Czaov6 & Jzaov6);
assign Czaov6 = (Qzaov6 & Xzaov6);
assign Qzaov6 = (~(E0bov6 & Lxydt6));
assign E0bov6 = (~(Euvnv6 & L0bov6));
assign Hyaov6 = (~(S0bov6 & Qg2nv6));
assign X0l8v6 = (~(Z0bov6 & G1bov6));
assign G1bov6 = (~(Pw9ov6 & Kxb7z6[0]));
assign Z0bov6 = (N1bov6 & U1bov6);
assign U1bov6 = (~(Gv9ov6 & B2bov6));
assign N1bov6 = (Eu9ov6 | I2bov6);
assign Q0l8v6 = (~(P2bov6 & W2bov6));
assign W2bov6 = (~(D3bov6 & S7f7z6[5]));
assign J0l8v6 = (~(K3bov6 & R3bov6));
assign R3bov6 = (~(Y3bov6 & Yxf7z6[27]));
assign K3bov6 = (F4bov6 & M4bov6);
assign M4bov6 = (~(Rj2ov6 & Mtkdt6));
assign F4bov6 = (~(Yj2ov6 & Yxf7z6[31]));
assign C0l8v6 = (~(T4bov6 & A5bov6));
assign A5bov6 = (H5bov6 & O5bov6);
assign O5bov6 = (~(V5bov6 & C6bov6));
assign H5bov6 = (~(J6bov6 & Alf7z6[31]));
assign T4bov6 = (Q6bov6 & X6bov6);
assign X6bov6 = (~(Cqf7z6[15] & E7bov6));
assign Q6bov6 = (~(L0g7z6[31] & L7bov6));
assign Vzk8v6 = (~(S7bov6 & Z7bov6));
assign Z7bov6 = (G8bov6 & N8bov6);
assign N8bov6 = (~(Ubpdt6 & U8bov6));
assign G8bov6 = (B9bov6 & I9bov6);
assign I9bov6 = (~(Epmdt6 & P9bov6));
assign B9bov6 = (~(W9bov6 & Onf7z6[31]));
assign S7bov6 = (Dabov6 & Kabov6);
assign Kabov6 = (~(Rabov6 & L0g7z6[31]));
assign Dabov6 = (Yabov6 & Fbbov6);
assign Fbbov6 = (~(Mtkdt6 & Mbbov6));
assign Yabov6 = (~(L0g7z6[15] & Gcmnv6));
assign Ozk8v6 = (Tbbov6 ? vis_r0_o[31] : Ae2ov6);
assign Hzk8v6 = (~(Acbov6 & Hcbov6));
assign Hcbov6 = (Ocbov6 & Vcbov6);
assign Vcbov6 = (~(H02ov6 & Cv97z6));
assign Ocbov6 = (Cdbov6 & Jdbov6);
assign Jdbov6 = (C12ov6 | Yojnv6);
assign Yojnv6 = (Qdbov6 & Xdbov6);
assign Xdbov6 = (Eebov6 & Lebov6);
assign Lebov6 = (Sebov6 & Zebov6);
assign Zebov6 = (Gfbov6 & Nfbov6);
assign Nfbov6 = (~(vis_psp_o[29] & N32ov6));
assign Gfbov6 = (~(U32ov6 & Pic7z6[29]));
assign Sebov6 = (Ufbov6 & Bgbov6);
assign Bgbov6 = (~(vis_msp_o[29] & P42ov6));
assign Ufbov6 = (~(vis_r12_o[29] & W42ov6));
assign Eebov6 = (Igbov6 & Pgbov6);
assign Pgbov6 = (Wgbov6 & Dhbov6);
assign Dhbov6 = (~(vis_r11_o[29] & F62ov6));
assign Wgbov6 = (~(vis_r10_o[29] & M62ov6));
assign Igbov6 = (Khbov6 & Rhbov6);
assign Rhbov6 = (~(vis_r9_o[29] & H72ov6));
assign Khbov6 = (~(vis_r8_o[29] & O72ov6));
assign Qdbov6 = (Yhbov6 & Fibov6);
assign Fibov6 = (Mibov6 & Tibov6);
assign Tibov6 = (Ajbov6 & Hjbov6);
assign Hjbov6 = (~(vis_r7_o[29] & L92ov6));
assign Ajbov6 = (~(vis_r6_o[29] & S92ov6));
assign Mibov6 = (Ojbov6 & Vjbov6);
assign Vjbov6 = (~(vis_r5_o[29] & Na2ov6));
assign Ojbov6 = (~(vis_r4_o[29] & Ua2ov6));
assign Yhbov6 = (Ckbov6 & Jkbov6);
assign Jkbov6 = (Qkbov6 & Xkbov6);
assign Xkbov6 = (~(vis_r3_o[29] & Dc2ov6));
assign Qkbov6 = (~(vis_r2_o[29] & Kc2ov6));
assign Ckbov6 = (Elbov6 & Llbov6);
assign Llbov6 = (~(vis_r1_o[29] & Fd2ov6));
assign Elbov6 = (~(vis_r0_o[29] & Md2ov6));
assign Cdbov6 = (~(Td2ov6 & Slbov6));
assign Acbov6 = (Zlbov6 & Gmbov6);
assign Gmbov6 = (~(Ve2ov6 & vis_pc_o[29]));
assign Zlbov6 = (~(Fhc7z6[29] & Cf2ov6));
assign Azk8v6 = (~(Nmbov6 & Umbov6));
assign Umbov6 = (~(Bnbov6 & Qu1ov6));
assign Nmbov6 = (Inbov6 & Pnbov6);
assign Pnbov6 = (~(Hz9ov6 & S7gdt6));
assign Inbov6 = (~(Uf4ov6 & Aegdt6));
assign Aegdt6 = (~(Wnbov6 & Dobov6));
assign Dobov6 = (Rdnnv6 | Kobov6);
assign Rdnnv6 = (!S7gdt6);
assign Wnbov6 = (Gw1ov6 ? Yobov6 : Robov6);
assign Yobov6 = (~(Fpbov6 & Mpbov6));
assign Fpbov6 = (Uf4ov6 & Tpbov6);
assign Tpbov6 = (~(Aqbov6 & Hqbov6));
assign Hqbov6 = (~(Dte7z6[5] & V1c7z6[31]));
assign Aqbov6 = (Oqbov6 & Vqbov6);
assign Vqbov6 = (~(Crbov6 & Jrbov6));
assign Jrbov6 = (Dy1ov6 | Dte7z6[4]);
assign Crbov6 = (Esbov6 ? Xrbov6 : Qrbov6);
assign Esbov6 = (Lsbov6 & Ssbov6);
assign Ssbov6 = (~(Zsbov6 & Gtbov6));
assign Gtbov6 = (~(Ntbov6 & Utbov6));
assign Qrbov6 = (Iubov6 ? S7gdt6 : Bubov6);
assign Iubov6 = (Pubov6 & Wubov6);
assign Pubov6 = (~(Ntbov6 | Dvbov6));
assign Dvbov6 = (Utbov6 & Kvbov6);
assign Bubov6 = (Fwbov6 ? Yvbov6 : Rvbov6);
assign Oqbov6 = (~(Px1ov6 & Fhc7z6[29]));
assign Robov6 = (~(Mwbov6 & Twbov6));
assign Twbov6 = (~(Dte7z6[4] | Dte7z6[5]));
assign Mwbov6 = (L0g7z6[32] & Kobov6);
assign Kobov6 = (Mpbov6 & Uf4ov6);
assign Tyk8v6 = (~(Axbov6 & Hxbov6));
assign Hxbov6 = (Oxbov6 & Vxbov6);
assign Vxbov6 = (Eu9ov6 | Cybov6);
assign Oxbov6 = (Jybov6 & Qybov6);
assign Qybov6 = (~(Gv9ov6 & Slbov6));
assign Jybov6 = (~(Uv9ov6 & Cv97z6));
assign Axbov6 = (Xybov6 & Ezbov6);
assign Ezbov6 = (~(Pw9ov6 & Kxb7z6[29]));
assign Xybov6 = (Lzbov6 & Szbov6);
assign Szbov6 = (~(Kx9ov6 & vis_pc_o[29]));
assign Lzbov6 = (~(Gli7z6[29] & Rx9ov6));
assign Myk8v6 = (~(Zzbov6 & G0cov6));
assign G0cov6 = (N0cov6 & U0cov6);
assign U0cov6 = (Eu9ov6 | B1cov6);
assign N0cov6 = (I1cov6 & P1cov6);
assign P1cov6 = (~(Gv9ov6 & Ae2ov6));
assign I1cov6 = (~(Uv9ov6 & Wt97z6));
assign Zzbov6 = (W1cov6 & D2cov6);
assign D2cov6 = (~(Pw9ov6 & Kxb7z6[31]));
assign W1cov6 = (K2cov6 & R2cov6);
assign R2cov6 = (~(Kx9ov6 & vis_pc_o[31]));
assign K2cov6 = (~(Rx9ov6 & Gli7z6[31]));
assign Fyk8v6 = (~(Y2cov6 & F3cov6));
assign F3cov6 = (M3cov6 & T3cov6);
assign T3cov6 = (~(H02ov6 & Kv97z6));
assign M3cov6 = (A4cov6 & H4cov6);
assign H4cov6 = (C12ov6 | Sdknv6);
assign Sdknv6 = (O4cov6 & V4cov6);
assign V4cov6 = (C5cov6 & J5cov6);
assign J5cov6 = (Q5cov6 & X5cov6);
assign X5cov6 = (E6cov6 & L6cov6);
assign L6cov6 = (~(vis_psp_o[15] & N32ov6));
assign E6cov6 = (~(U32ov6 & Pic7z6[15]));
assign Q5cov6 = (S6cov6 & Z6cov6);
assign Z6cov6 = (~(vis_msp_o[15] & P42ov6));
assign S6cov6 = (~(vis_r12_o[15] & W42ov6));
assign C5cov6 = (G7cov6 & N7cov6);
assign N7cov6 = (U7cov6 & B8cov6);
assign B8cov6 = (~(vis_r11_o[15] & F62ov6));
assign U7cov6 = (~(vis_r10_o[15] & M62ov6));
assign G7cov6 = (I8cov6 & P8cov6);
assign P8cov6 = (~(vis_r9_o[15] & H72ov6));
assign I8cov6 = (~(vis_r8_o[15] & O72ov6));
assign O4cov6 = (W8cov6 & D9cov6);
assign D9cov6 = (K9cov6 & R9cov6);
assign R9cov6 = (Y9cov6 & Facov6);
assign Facov6 = (~(vis_r7_o[15] & L92ov6));
assign Y9cov6 = (~(vis_r6_o[15] & S92ov6));
assign K9cov6 = (Macov6 & Tacov6);
assign Tacov6 = (~(vis_r5_o[15] & Na2ov6));
assign Macov6 = (~(vis_r4_o[15] & Ua2ov6));
assign W8cov6 = (Abcov6 & Hbcov6);
assign Hbcov6 = (Obcov6 & Vbcov6);
assign Vbcov6 = (~(vis_r3_o[15] & Dc2ov6));
assign Obcov6 = (~(vis_r2_o[15] & Kc2ov6));
assign Abcov6 = (Cccov6 & Jccov6);
assign Jccov6 = (~(vis_r1_o[15] & Fd2ov6));
assign Cccov6 = (~(vis_r0_o[15] & Md2ov6));
assign A4cov6 = (~(Td2ov6 & Qccov6));
assign Y2cov6 = (Xccov6 & Edcov6);
assign Edcov6 = (~(Ve2ov6 & vis_pc_o[15]));
assign Xccov6 = (~(Fhc7z6[15] & Cf2ov6));
assign Yxk8v6 = (~(Ldcov6 & Sdcov6));
assign Sdcov6 = (~(B987v6 & I0snv6));
assign Ldcov6 = (~(Zdcov6 & Gecov6));
assign Zdcov6 = (~(Necov6 & Uecov6));
assign Uecov6 = (Bfcov6 & Ifcov6);
assign Ifcov6 = (~(Pfcov6 | Wfcov6));
assign Pfcov6 = (TSVALUEB[10] ^ Gnzmz6[11]);
assign Bfcov6 = (Dgcov6 & Kgcov6);
assign Kgcov6 = (~(TSVALUEB[11] ^ Gnzmz6[12]));
assign Dgcov6 = (~(TSVALUEB[12] ^ Gnzmz6[13]));
assign Necov6 = (Rgcov6 & Ygcov6);
assign Ygcov6 = (Fhcov6 & Mhcov6);
assign Mhcov6 = (~(TSVALUEB[13] ^ Gnzmz6[14]));
assign Fhcov6 = (~(TSVALUEB[7] ^ Gnzmz6[8]));
assign Rgcov6 = (Thcov6 & Aicov6);
assign Aicov6 = (~(TSVALUEB[8] ^ Gnzmz6[9]));
assign Thcov6 = (~(TSVALUEB[9] ^ Gnzmz6[10]));
assign Rxk8v6 = (~(Hicov6 & Oicov6));
assign Oicov6 = (~(Vicov6 & Fed7v6));
assign Hicov6 = (~(Cjcov6 & Jjcov6));
assign Jjcov6 = (Qjcov6 & Xjcov6);
assign Xjcov6 = (~(Ekcov6 & Lkcov6));
assign Ekcov6 = (Xfd7v6 ^ Ocd7v6);
assign Cjcov6 = (Skcov6 & Zkcov6);
assign Zkcov6 = (~(Glcov6 & Nlcov6));
assign Glcov6 = (~(Ulcov6 & Bmcov6));
assign Bmcov6 = (Imcov6 & Pmcov6);
assign Pmcov6 = (Wmcov6 & Fftnv6);
assign Imcov6 = (Dncov6 & Kncov6);
assign Kncov6 = (E11nz6[0] ^ E5d7v6);
assign Dncov6 = (~(Rncov6 ^ E11nz6[4]));
assign Ulcov6 = (Yncov6 & Focov6);
assign Focov6 = (Mocov6 ^ Tocov6);
assign Yncov6 = (Apcov6 & Hpcov6);
assign Hpcov6 = (~(Opcov6 ^ E11nz6[3]));
assign Apcov6 = (~(Y3d7v6 ^ E11nz6[1]));
assign Kxk8v6 = (~(Lyrnv6 ^ Wmcov6));
assign Dxk8v6 = (Wmcov6 ? Rncov6 : Rr0nz6[1]);
assign Rncov6 = (Vpcov6 & Lkcov6);
assign Vpcov6 = (~(Owrnv6 ^ Cqcov6));
assign Cqcov6 = (Jqcov6 & Rr0nz6[0]);
assign Wwk8v6 = (Wmcov6 ? Y3d7v6 : Hw0nz6[1]);
assign Y3d7v6 = (Lyrnv6 ^ Qqcov6);
assign Pwk8v6 = (Wmcov6 ? Tocov6 : Hw0nz6[2]);
assign Tocov6 = (~(Xqcov6 & Eyrnv6));
assign Xqcov6 = (Lyrnv6 ? Ercov6 : Xxrnv6);
assign Iwk8v6 = (Wmcov6 ? Opcov6 : Rr0nz6[0]);
assign Opcov6 = (Lrcov6 & Lkcov6);
assign Lrcov6 = (~(Cxrnv6 ^ Jqcov6));
assign Jqcov6 = (~(Srcov6 | Lyrnv6));
assign Bwk8v6 = (~(Zrcov6 & Gscov6));
assign Gscov6 = (~(Ft0nz6[4] & Nscov6));
assign Nscov6 = (~(Uscov6 & Btcov6));
assign Btcov6 = (~(Ft0nz6[3] & Itcov6));
assign Zrcov6 = (~(Spc7v6 & Ptcov6));
assign Ptcov6 = (~(Wtcov6 ^ Tvrnv6));
assign Wtcov6 = (Ducov6 & Fvrnv6);
assign Uvk8v6 = (~(Kucov6 & Rucov6));
assign Rucov6 = (~(Spc7v6 & Yucov6));
assign Yucov6 = (Fvcov6 ^ Durnv6);
assign Kucov6 = (Ft0nz6[1] ? Tvcov6 : Mvcov6);
assign Mvcov6 = (Awcov6 | Ft0nz6[0]);
assign Nvk8v6 = (~(Hwcov6 & Owcov6));
assign Hwcov6 = (Vwcov6 & Cxcov6);
assign Cxcov6 = (~(Ft0nz6[2] & Jxcov6));
assign Jxcov6 = (~(Tvcov6 & Qxcov6));
assign Qxcov6 = (~(Ft0nz6[1] & Itcov6));
assign Tvcov6 = (Xxcov6 & Eycov6);
assign Eycov6 = (~(Itcov6 & Ft0nz6[0]));
assign Vwcov6 = (~(Spc7v6 & Lycov6));
assign Lycov6 = (Sycov6 ^ Qqrnv6);
assign Gvk8v6 = (~(Zycov6 & Gzcov6));
assign Gzcov6 = (~(Spc7v6 & Nzcov6));
assign Nzcov6 = (~(Ducov6 ^ Imrnv6));
assign Ducov6 = (~(Sycov6 | Qqrnv6));
assign Sycov6 = (Fvcov6 | Durnv6);
assign Fvcov6 = (Gsrnv6 | Uzcov6);
assign Zycov6 = (Ft0nz6[3] ? Uscov6 : Owcov6);
assign Uscov6 = (Xxcov6 & B0dov6);
assign B0dov6 = (Awcov6 | I0dov6);
assign Owcov6 = (~(Itcov6 & I0dov6));
assign Itcov6 = (!Awcov6);
assign Zuk8v6 = (~(P0dov6 & W0dov6));
assign W0dov6 = (~(D1dov6 & Spc7v6));
assign D1dov6 = (~(Errnv6 ^ Uzcov6));
assign P0dov6 = (K1dov6 ? Awcov6 : Xxcov6);
assign Awcov6 = (~(R1dov6 & Qjrnv6));
assign Qjrnv6 = (~(Y1dov6 & I0dov6));
assign I0dov6 = (F2dov6 & K1dov6);
assign F2dov6 = (~(Ft0nz6[1] | Ft0nz6[2]));
assign Y1dov6 = (~(Ft0nz6[3] | Ft0nz6[4]));
assign R1dov6 = (~(M2dov6 | Spc7v6));
assign Xxcov6 = (!M2dov6);
assign M2dov6 = (~(T2dov6 | Spc7v6));
assign T2dov6 = (~(A3dov6 | H3dov6));
assign Suk8v6 = (V3dov6 ? H71nz6[1] : O3dov6);
assign O3dov6 = (Tvd7v6 | C4dov6);
assign Luk8v6 = (V3dov6 ? H71nz6[8] : J4dov6);
assign J4dov6 = (Bmd7v6 | C4dov6);
assign Euk8v6 = (V3dov6 ? H71nz6[7] : Q4dov6);
assign Q4dov6 = (Lnd7v6 | C4dov6);
assign Xtk8v6 = (V3dov6 ? H71nz6[6] : X4dov6);
assign X4dov6 = (Vod7v6 | C4dov6);
assign Qtk8v6 = (V3dov6 ? H71nz6[5] : E5dov6);
assign E5dov6 = (Fqd7v6 | C4dov6);
assign Jtk8v6 = (V3dov6 ? H71nz6[4] : L5dov6);
assign L5dov6 = (Prd7v6 | C4dov6);
assign Ctk8v6 = (V3dov6 ? H71nz6[3] : S5dov6);
assign S5dov6 = (Zsd7v6 | C4dov6);
assign Vsk8v6 = (V3dov6 ? H71nz6[2] : Z5dov6);
assign Z5dov6 = (Jud7v6 | C4dov6);
assign Osk8v6 = (V3dov6 ? H71nz6[0] : G6dov6);
assign V3dov6 = (~(N6dov6 | U6dov6));
assign U6dov6 = (Sr5ov6 & Jrqnv6);
assign G6dov6 = (Dxd7v6 | C4dov6);
assign Hsk8v6 = (I7dov6 ? B7dov6 : Uh77v6);
assign B7dov6 = (P7dov6 & W7dov6);
assign W7dov6 = (D8dov6 & K8dov6);
assign K8dov6 = (R8dov6 & Y8dov6);
assign Y8dov6 = (~(F9dov6 | Ruymz6[7]));
assign F9dov6 = (Ruymz6[8] | Ruymz6[9]);
assign R8dov6 = (~(Ruymz6[5] | Ruymz6[6]));
assign D8dov6 = (M9dov6 & T9dov6);
assign T9dov6 = (~(Ruymz6[3] | Ruymz6[4]));
assign M9dov6 = (~(Ruymz6[1] | Ruymz6[2]));
assign P7dov6 = (Aadov6 & Hadov6);
assign Hadov6 = (Oadov6 & Vadov6);
assign Vadov6 = (~(Ruymz6[14] | Ruymz6[15]));
assign Oadov6 = (~(Ruymz6[12] | Ruymz6[13]));
assign Aadov6 = (Cbdov6 & Jbdov6);
assign Jbdov6 = (~(Ruymz6[10] | Ruymz6[11]));
assign Cbdov6 = (Ruymz6[0] & Y9rnv6);
assign Ask8v6 = (~(Qbdov6 & Xbdov6));
assign Xbdov6 = (Ecdov6 & Lcdov6);
assign Lcdov6 = (Scdov6 & Zcdov6);
assign Zcdov6 = (Gddov6 & Nddov6);
assign Nddov6 = (Uddov6 & Bedov6);
assign Bedov6 = (Iedov6 & Pedov6);
assign Pedov6 = (~(Hvw7v6 & Wedov6));
assign Iedov6 = (Dfdov6 & Kfdov6);
assign Kfdov6 = (~(Rtw7v6 & Rfdov6));
assign Dfdov6 = (~(Avw7v6 & Yfdov6));
assign Uddov6 = (Fgdov6 & Mgdov6);
assign Mgdov6 = (~(Vvw7v6 & Tgdov6));
assign Fgdov6 = (~(Jww7v6 & Ahdov6));
assign Gddov6 = (Hhdov6 & Ohdov6);
assign Ohdov6 = (Vhdov6 & Cidov6);
assign Cidov6 = (~(Zxw7v6 & Jidov6));
assign Vhdov6 = (Qidov6 & Xidov6);
assign Xidov6 = (~(Xww7v6 & Ejdov6));
assign Qidov6 = (~(Lxw7v6 & Ljdov6));
assign Hhdov6 = (Sjdov6 & Zjdov6);
assign Zjdov6 = (~(Nyw7v6 & Gkdov6));
assign Sjdov6 = (~(Bzw7v6 & Nkdov6));
assign Scdov6 = (Ukdov6 & Bldov6);
assign Bldov6 = (Ildov6 & Pldov6);
assign Pldov6 = (Wldov6 & Dmdov6);
assign Dmdov6 = (~(R0x7v6 & Kmdov6));
assign Wldov6 = (Rmdov6 & Ymdov6);
assign Ymdov6 = (~(Pzw7v6 & Fndov6));
assign Rmdov6 = (~(D0x7v6 & Mndov6));
assign Ildov6 = (Tndov6 & Aodov6);
assign Aodov6 = (~(F1x7v6 & Hodov6));
assign Tndov6 = (~(T1x7v6 & Oodov6));
assign Ukdov6 = (Vodov6 & Cpdov6);
assign Cpdov6 = (Jpdov6 & Qpdov6);
assign Qpdov6 = (~(H2x7v6 & Xpdov6));
assign Jpdov6 = (~(V2x7v6 & Eqdov6));
assign Vodov6 = (Lqdov6 & Sqdov6);
assign Sqdov6 = (~(J3x7v6 & Zqdov6));
assign Lqdov6 = (~(X3x7v6 & Grdov6));
assign Ecdov6 = (Nrdov6 & Urdov6);
assign Urdov6 = (Bsdov6 & Isdov6);
assign Isdov6 = (Psdov6 & Wsdov6);
assign Wsdov6 = (Dtdov6 & Ktdov6);
assign Ktdov6 = (~(N5x7v6 & Rtdov6));
assign Dtdov6 = (Ytdov6 & Fudov6);
assign Fudov6 = (~(L4x7v6 & Mudov6));
assign Ytdov6 = (~(Z4x7v6 & Tudov6));
assign Psdov6 = (Avdov6 & Hvdov6);
assign Hvdov6 = (~(B6x7v6 & Ovdov6));
assign Avdov6 = (~(P6x7v6 & Vvdov6));
assign Bsdov6 = (Cwdov6 & Jwdov6);
assign Jwdov6 = (Qwdov6 & Xwdov6);
assign Xwdov6 = (~(D7x7v6 & Exdov6));
assign Qwdov6 = (~(R7x7v6 & Lxdov6));
assign Cwdov6 = (Sxdov6 & Zxdov6);
assign Zxdov6 = (~(F8x7v6 & Gydov6));
assign Sxdov6 = (~(T8x7v6 & Nydov6));
assign Nrdov6 = (Uydov6 & Bzdov6);
assign Bzdov6 = (Izdov6 & Pzdov6);
assign Pzdov6 = (Wzdov6 & D0eov6);
assign D0eov6 = (~(Jax7v6 & K0eov6));
assign Wzdov6 = (R0eov6 & Y0eov6);
assign Y0eov6 = (~(H9x7v6 & F1eov6));
assign R0eov6 = (~(V9x7v6 & M1eov6));
assign Izdov6 = (T1eov6 & A2eov6);
assign A2eov6 = (~(Xax7v6 & H2eov6));
assign T1eov6 = (~(Lbx7v6 & O2eov6));
assign Uydov6 = (V2eov6 & C3eov6);
assign C3eov6 = (J3eov6 & Q3eov6);
assign Q3eov6 = (~(Zbx7v6 & X3eov6));
assign J3eov6 = (~(Ncx7v6 & E4eov6));
assign V2eov6 = (L4eov6 & S4eov6);
assign S4eov6 = (Z4eov6 | Zfcet6);
assign L4eov6 = (~(Pdx7v6 & G5eov6));
assign Qbdov6 = (N5eov6 & U5eov6);
assign U5eov6 = (B6eov6 & I6eov6);
assign I6eov6 = (P6eov6 & W6eov6);
assign W6eov6 = (D7eov6 & K7eov6);
assign K7eov6 = (R7eov6 & Y7eov6);
assign Y7eov6 = (~(Nr38v6 & F8eov6));
assign R7eov6 = (M8eov6 & T8eov6);
assign T8eov6 = (~(Lq38v6 & A9eov6));
assign M8eov6 = (~(Zq38v6 & H9eov6));
assign D7eov6 = (O9eov6 & V9eov6);
assign V9eov6 = (~(Bs38v6 & Caeov6));
assign O9eov6 = (~(Ps38v6 & Jaeov6));
assign P6eov6 = (Qaeov6 & Xaeov6);
assign Xaeov6 = (Ebeov6 & Lbeov6);
assign Lbeov6 = (~(Dt38v6 & Sbeov6));
assign Ebeov6 = (~(Rt38v6 & Zbeov6));
assign Qaeov6 = (Gceov6 & Nceov6);
assign Nceov6 = (~(Fu38v6 & Uceov6));
assign Gceov6 = (~(Tu38v6 & Bdeov6));
assign B6eov6 = (Ideov6 & Pdeov6);
assign Pdeov6 = (Wdeov6 & Deeov6);
assign Deeov6 = (Keeov6 & Reeov6);
assign Reeov6 = (~(Jw38v6 & Yeeov6));
assign Keeov6 = (Ffeov6 & Mfeov6);
assign Mfeov6 = (~(Hv38v6 & Tfeov6));
assign Ffeov6 = (~(Vv38v6 & Ageov6));
assign Wdeov6 = (Hgeov6 & Ogeov6);
assign Ogeov6 = (~(Xw38v6 & Vgeov6));
assign Hgeov6 = (~(Lx38v6 & Cheov6));
assign Ideov6 = (Jheov6 & Qheov6);
assign Qheov6 = (Xheov6 & Eieov6);
assign Eieov6 = (~(Zx38v6 & Lieov6));
assign Xheov6 = (~(Ny38v6 & Sieov6));
assign Jheov6 = (Zieov6 & Gjeov6);
assign Gjeov6 = (~(Bz38v6 & Njeov6));
assign Zieov6 = (~(Pz38v6 & Ujeov6));
assign N5eov6 = (Bkeov6 & Ikeov6);
assign Ikeov6 = (Pkeov6 & Wkeov6);
assign Wkeov6 = (Dleov6 & Kleov6);
assign Kleov6 = (Rleov6 & Yleov6);
assign Yleov6 = (~(F148v6 & Fmeov6));
assign Rleov6 = (Mmeov6 & Tmeov6);
assign Tmeov6 = (~(D048v6 & Aneov6));
assign Mmeov6 = (~(R048v6 & Hneov6));
assign Dleov6 = (Oneov6 & Vneov6);
assign Vneov6 = (~(T148v6 & Coeov6));
assign Oneov6 = (~(H248v6 & Joeov6));
assign Pkeov6 = (Qoeov6 & Xoeov6);
assign Xoeov6 = (Epeov6 & Lpeov6);
assign Lpeov6 = (~(V248v6 & Speov6));
assign Epeov6 = (~(J348v6 & Zpeov6));
assign Qoeov6 = (Gqeov6 & Nqeov6);
assign Nqeov6 = (~(X348v6 & Uqeov6));
assign Gqeov6 = (~(L448v6 & Breov6));
assign Bkeov6 = (Ireov6 & Preov6);
assign Preov6 = (Wreov6 & Dseov6);
assign Dseov6 = (Kseov6 & Rseov6);
assign Rseov6 = (~(Qfk8v6 & Yseov6));
assign Kseov6 = (Fteov6 & Mteov6);
assign Mteov6 = (~(Z448v6 & Tteov6));
assign Fteov6 = (~(Vek8v6 & Aueov6));
assign Wreov6 = (Hueov6 & Oueov6);
assign Oueov6 = (~(Xfk8v6 & Vueov6));
assign Hueov6 = (~(Sgk8v6 & Cveov6));
assign Ireov6 = (Jveov6 & Qveov6);
assign Qveov6 = (Xveov6 & Eweov6);
assign Eweov6 = (~(Nhk8v6 & Lweov6));
assign Xveov6 = (~(Djk8v6 & Sweov6));
assign Jveov6 = (Zweov6 & Gxeov6);
assign Gxeov6 = (~(Yjk8v6 & Nxeov6));
assign Zweov6 = (~(Yqk8v6 & Uxeov6));
assign Trk8v6 = (~(Byeov6 & Iyeov6));
assign Iyeov6 = (Pyeov6 | Wyeov6);
assign Mrk8v6 = (Dzeov6 & Kzeov6);
assign Kzeov6 = (Wyeov6 ? Yzeov6 : Rzeov6);
assign Yzeov6 = (D2fet6 & F0fov6);
assign F0fov6 = (Tnzdt6 | SLEEPHOLDREQn);
assign Rzeov6 = (M0fov6 & T0fov6);
assign Frk8v6 = (~(A1fov6 & H1fov6));
assign H1fov6 = (~(INTISR[63] & O1fov6));
assign A1fov6 = (~(U697z6 & V1fov6));
assign Yqk8v6 = (~(C2fov6 & J2fov6));
assign J2fov6 = (~(Q2fov6 & X2fov6));
assign X2fov6 = (~(Jqj7z6[1] & X3get6));
assign Q2fov6 = (Qmj7z6[1] & Uxeov6);
assign C2fov6 = (~(V5get6 & E3fov6));
assign E3fov6 = (~(L3fov6 & Cn2nv6));
assign Rqk8v6 = (Cn2nv6 ? L3fov6 : S3fov6);
assign S3fov6 = (~(Z3fov6 & G4fov6));
assign G4fov6 = (~(N4fov6 & U4fov6));
assign Kqk8v6 = (Zs4ov6 ? Xz7et6 : B5fov6);
assign B5fov6 = (~(Dtadt6 & I5fov6));
assign Dqk8v6 = (W5fov6 ? Pjb7z6[19] : P5fov6);
assign Ppk8v6 = (~(Wfo7v6 & D6fov6));
assign D6fov6 = (~(K6fov6 & Ke2ft6));
assign Ipk8v6 = (~(R6fov6 & Y6fov6));
assign Y6fov6 = (~(F7fov6 & Em5ft6));
assign F7fov6 = (M7fov6 & Wdtnv6);
assign M7fov6 = (Hk5ft6 | V1gnv6);
assign R6fov6 = (~(K6fov6 & Hk5ft6));
assign Bpk8v6 = (~(T7fov6 & A8fov6));
assign A8fov6 = (~(Bxi7z6[2] & H8fov6));
assign H8fov6 = (~(O8fov6 & I52nv6));
assign T7fov6 = (~(V8fov6 & C9fov6));
assign V8fov6 = (~(J9fov6 & Q9fov6));
assign Q9fov6 = (~(X9fov6 | Eafov6));
assign J9fov6 = (~(L99ov6 | Lafov6));
assign Uok8v6 = (Pb9ov6 ? D6c7z6[2] : Safov6);
assign Safov6 = (~(Zafov6 & Gbfov6));
assign Gbfov6 = (Nbfov6 & Ubfov6);
assign Ubfov6 = (~(Yc9ov6 & Bcfov6));
assign Nbfov6 = (~(Md9ov6 & Icfov6));
assign Zafov6 = (Pcfov6 & Wcfov6);
assign Wcfov6 = (~(Oe9ov6 & Ddfov6));
assign Pcfov6 = (~(Cf9ov6 & Kdfov6));
assign Nok8v6 = (~(Rdfov6 & Ydfov6));
assign Ydfov6 = (~(E3c7z6[0] & Cf2ov6));
assign Rdfov6 = (Fefov6 & Mefov6);
assign Mefov6 = (C12ov6 | Tefov6);
assign Fefov6 = (~(Td2ov6 & B2bov6));
assign Gok8v6 = (Hffov6 ? Inadt6 : Affov6);
assign Hffov6 = (Offov6 & Vffov6);
assign Vffov6 = (~(Cgfov6 & Jgfov6));
assign Jgfov6 = (~(Qgfov6 & Xgfov6));
assign Qgfov6 = (Ehfov6 & Lhfov6);
assign Ehfov6 = (~(Shfov6 & Zhfov6));
assign Zhfov6 = (~(Gifov6 & Nifov6));
assign Nifov6 = (~(I9e7z6[1] & Uifov6));
assign Uifov6 = (~(I9e7z6[0] & Xsinv6));
assign Gifov6 = (~(Ibe7z6[3] & Bjfov6));
assign Bjfov6 = (~(E3c7z6[0] & Xsinv6));
assign Affov6 = (Ijfov6 & Offov6);
assign Ijfov6 = (~(Pjfov6 & Wjfov6));
assign Wjfov6 = (Dkfov6 & Kkfov6);
assign Dkfov6 = (~(Rkfov6 & Ykfov6));
assign Pjfov6 = (Flfov6 & Xgfov6);
assign Xgfov6 = (~(Ieadt6 & Mlfov6));
assign Znk8v6 = (~(Tlfov6 & Amfov6));
assign Amfov6 = (~(Hmfov6 & Omfov6));
assign Omfov6 = (Vmfov6 & Cnfov6);
assign Cnfov6 = (Jnfov6 | Qnfov6);
assign Vmfov6 = (Xnfov6 & SLEEPHOLDACKn);
assign Hmfov6 = (Eofov6 & Lofov6);
assign Lofov6 = (F02nv6 | Cwadt6);
assign Tlfov6 = (~(Sofov6 & Zofov6));
assign Sofov6 = (Nneet6 & Ldo7v6);
assign Snk8v6 = (~(Gpfov6 & Npfov6));
assign Npfov6 = (~(Upfov6 & Ohe7z6[2]));
assign Lnk8v6 = (~(Bqfov6 & Iqfov6));
assign Iqfov6 = (~(Gnaov6 & Tcinv6));
assign Tcinv6 = (~(Pqfov6 & Qg2nv6));
assign Pqfov6 = (Hdinv6 | Wqfov6);
assign Hdinv6 = (~(Drfov6 & Krfov6));
assign Krfov6 = (Rrfov6 | Yrfov6);
assign Rrfov6 = (Fsfov6 & Msfov6);
assign Msfov6 = (!Cmbdt6);
assign Bqfov6 = (~(Iufdt6 & Vs9ov6));
assign Enk8v6 = (~(Tsfov6 & Atfov6));
assign Atfov6 = (~(Htfov6 & Qu1ov6));
assign Tsfov6 = (Otfov6 & Vtfov6);
assign Vtfov6 = (~(Cufov6 & Jufov6));
assign Cufov6 = (Uf4ov6 & Qufov6);
assign Qufov6 = (~(Px1ov6 & Xufov6));
assign Xufov6 = (!Fhc7z6[27]);
assign Uf4ov6 = (!Wg4ov6);
assign Otfov6 = (~(Lsfdt6 & Evfov6));
assign Evfov6 = (~(Ig4ov6 & Lvfov6));
assign Lvfov6 = (Wg4ov6 | Jufov6);
assign Ig4ov6 = (!Hz9ov6);
assign Hz9ov6 = (Svfov6 & Wg4ov6);
assign Wg4ov6 = (~(Zvfov6 & Gwfov6));
assign Gwfov6 = (~(Nwfov6 & Uwfov6));
assign Uwfov6 = (~(Iufdt6 & Knbdt6));
assign Nwfov6 = (~(Yrfov6 | Lwfdt6));
assign Zvfov6 = (Bg4ov6 | Jufov6);
assign Jufov6 = (Bxfov6 & Ixfov6);
assign Bxfov6 = (Pxfov6 & Wxfov6);
assign Wxfov6 = (~(Dyfov6 & Q0aov6));
assign Q0aov6 = (~(Px1ov6 & I0c7z6[1]));
assign Dyfov6 = (Kyfov6 & Ryfov6);
assign Kyfov6 = (~(Yyfov6 & Fzfov6));
assign Yyfov6 = (Mzfov6 & V5bov6);
assign Bg4ov6 = (Mpbov6 | Tzfov6);
assign Tzfov6 = (A0gov6 & Dte7z6[18]);
assign A0gov6 = (Ixfov6 & Pxfov6);
assign Mpbov6 = (H0gov6 & Ixfov6);
assign H0gov6 = (Pxfov6 & O0gov6);
assign O0gov6 = (V0gov6 | Dte7z6[19]);
assign V0gov6 = (Px1ov6 & I0c7z6[1]);
assign Px1ov6 = (C1gov6 & J1gov6);
assign Xmk8v6 = (~(Q1gov6 & X1gov6));
assign X1gov6 = (E2gov6 & L2gov6);
assign L2gov6 = (~(Td2ov6 & S2gov6));
assign E2gov6 = (Z2gov6 & G3gov6);
assign G3gov6 = (C12ov6 | Esjnv6);
assign Esjnv6 = (N3gov6 & U3gov6);
assign U3gov6 = (B4gov6 & I4gov6);
assign I4gov6 = (P4gov6 & W4gov6);
assign W4gov6 = (D5gov6 & K5gov6);
assign K5gov6 = (~(vis_psp_o[27] & N32ov6));
assign D5gov6 = (~(U32ov6 & Pic7z6[27]));
assign P4gov6 = (R5gov6 & Y5gov6);
assign Y5gov6 = (~(vis_msp_o[27] & P42ov6));
assign R5gov6 = (~(vis_r12_o[27] & W42ov6));
assign B4gov6 = (F6gov6 & M6gov6);
assign M6gov6 = (T6gov6 & A7gov6);
assign A7gov6 = (~(vis_r11_o[27] & F62ov6));
assign T6gov6 = (~(vis_r10_o[27] & M62ov6));
assign F6gov6 = (H7gov6 & O7gov6);
assign O7gov6 = (~(vis_r9_o[27] & H72ov6));
assign H7gov6 = (~(vis_r8_o[27] & O72ov6));
assign N3gov6 = (V7gov6 & C8gov6);
assign C8gov6 = (J8gov6 & Q8gov6);
assign Q8gov6 = (X8gov6 & E9gov6);
assign E9gov6 = (~(vis_r7_o[27] & L92ov6));
assign X8gov6 = (~(vis_r6_o[27] & S92ov6));
assign J8gov6 = (L9gov6 & S9gov6);
assign S9gov6 = (~(vis_r5_o[27] & Na2ov6));
assign L9gov6 = (~(vis_r4_o[27] & Ua2ov6));
assign V7gov6 = (Z9gov6 & Gagov6);
assign Gagov6 = (Nagov6 & Uagov6);
assign Uagov6 = (~(vis_r3_o[27] & Dc2ov6));
assign Nagov6 = (~(vis_r2_o[27] & Kc2ov6));
assign Z9gov6 = (Bbgov6 & Ibgov6);
assign Ibgov6 = (~(vis_r1_o[27] & Fd2ov6));
assign Bbgov6 = (~(vis_r0_o[27] & Md2ov6));
assign Z2gov6 = (~(H02ov6 & Sv97z6));
assign Q1gov6 = (Pbgov6 & Wbgov6);
assign Wbgov6 = (~(Ve2ov6 & vis_pc_o[27]));
assign Pbgov6 = (~(Fhc7z6[27] & Cf2ov6));
assign Qmk8v6 = (~(Dcgov6 & Kcgov6));
assign Kcgov6 = (Rcgov6 & Ycgov6);
assign Ycgov6 = (~(H02ov6 & Mu97z6));
assign Rcgov6 = (Fdgov6 & Mdgov6);
assign Mdgov6 = (C12ov6 | H4knv6);
assign H4knv6 = (Tdgov6 & Aegov6);
assign Aegov6 = (Hegov6 & Oegov6);
assign Oegov6 = (Vegov6 & Cfgov6);
assign Cfgov6 = (Jfgov6 & Qfgov6);
assign Qfgov6 = (~(Pic7z6[1] & U32ov6));
assign Jfgov6 = (~(vis_r12_o[1] & W42ov6));
assign Vegov6 = (Xfgov6 & Eggov6);
assign Eggov6 = (~(vis_r11_o[1] & F62ov6));
assign Xfgov6 = (~(vis_r10_o[1] & M62ov6));
assign Hegov6 = (Lggov6 & Sggov6);
assign Sggov6 = (~(vis_r7_o[1] & L92ov6));
assign Lggov6 = (Zggov6 & Ghgov6);
assign Ghgov6 = (~(vis_r9_o[1] & H72ov6));
assign Zggov6 = (~(vis_r8_o[1] & O72ov6));
assign Tdgov6 = (Nhgov6 & Uhgov6);
assign Uhgov6 = (Bigov6 & Iigov6);
assign Iigov6 = (Pigov6 & Wigov6);
assign Wigov6 = (~(vis_r6_o[1] & S92ov6));
assign Pigov6 = (~(vis_r5_o[1] & Na2ov6));
assign Bigov6 = (Djgov6 & Kjgov6);
assign Kjgov6 = (~(vis_r4_o[1] & Ua2ov6));
assign Djgov6 = (~(vis_r3_o[1] & Dc2ov6));
assign Nhgov6 = (Rjgov6 & Yjgov6);
assign Yjgov6 = (~(vis_r0_o[1] & Md2ov6));
assign Rjgov6 = (Fkgov6 & Mkgov6);
assign Mkgov6 = (~(vis_r2_o[1] & Kc2ov6));
assign Fkgov6 = (~(vis_r1_o[1] & Fd2ov6));
assign Fdgov6 = (~(Td2ov6 & Nv9ov6));
assign Dcgov6 = (Tkgov6 & Algov6);
assign Algov6 = (~(Ve2ov6 & vis_pc_o[1]));
assign Tkgov6 = (~(E3c7z6[1] & Cf2ov6));
assign Jmk8v6 = (~(Hlgov6 & Olgov6));
assign Olgov6 = (~(Vlgov6 & Ppb7z6[7]));
assign Hlgov6 = (Cmgov6 & Jmgov6);
assign Jmgov6 = (Qmgov6 | Zmaov6);
assign Cmgov6 = (~(Xmgov6 & Fhc7z6[7]));
assign Cmk8v6 = (~(Engov6 & Lngov6));
assign Lngov6 = (~(Vlgov6 & Ppb7z6[5]));
assign Engov6 = (Sngov6 & Zngov6);
assign Zngov6 = (Qmgov6 | Ivaov6);
assign Sngov6 = (~(Xmgov6 & Fhc7z6[5]));
assign Vlk8v6 = (~(Gogov6 & Nogov6));
assign Nogov6 = (~(Vlgov6 & Ppb7z6[6]));
assign Gogov6 = (Uogov6 & Bpgov6);
assign Bpgov6 = (Qmgov6 | Fqaov6);
assign Qmgov6 = (Ipgov6 | Vlgov6);
assign Uogov6 = (~(Xmgov6 & Fhc7z6[6]));
assign Xmgov6 = (Ipgov6 & Ppgov6);
assign Ppgov6 = (!Vlgov6);
assign Vlgov6 = (Wpgov6 & Dqgov6);
assign Wpgov6 = (~(Kqgov6 & Rqgov6));
assign Rqgov6 = (Yqgov6 | Ibe7z6[1]);
assign Yqgov6 = (Ibe7z6[2] & Frgov6);
assign Olk8v6 = (Trgov6 ? Mrgov6 : Moj7z6[2]);
assign Hlk8v6 = (Trgov6 ? Asgov6 : Moj7z6[1]);
assign Alk8v6 = (S93nv6 ? P2j7z6[6] : Hsgov6);
assign Tkk8v6 = (S93nv6 ? P2j7z6[5] : Osgov6);
assign Mkk8v6 = (Vsgov6 & Ctgov6);
assign Ctgov6 = (~(Jtgov6 & Qtgov6));
assign Qtgov6 = (~(Xtgov6 & X7get6));
assign Xtgov6 = (Eugov6 & Lugov6);
assign Jtgov6 = (~(Ib3nv6 & Sugov6));
assign Fkk8v6 = (Fjadt6 ? Gvgov6 : Zugov6);
assign Gvgov6 = (~(Z3fov6 & Nvgov6));
assign Nvgov6 = (~(Uvgov6 & U4fov6));
assign Zugov6 = (~(Bwgov6 & Iwgov6));
assign Iwgov6 = (~(Pwgov6 & X7get6));
assign Pwgov6 = (~(Wwgov6 | Dxgov6));
assign Bwgov6 = (Kxgov6 | Rxgov6);
assign Yjk8v6 = (~(Yxgov6 & Fygov6));
assign Fygov6 = (~(Mygov6 & Fjadt6));
assign Mygov6 = (S3a7z6 & Tygov6);
assign Tygov6 = (!Jqj7z6[0]);
assign Yxgov6 = (Hdcet6 ? Hzgov6 : Azgov6);
assign Hzgov6 = (Ozgov6 & Vzgov6);
assign Ozgov6 = (~(Rxgov6 | Fjadt6));
assign Azgov6 = (C0hov6 & J0hov6);
assign J0hov6 = (~(Q0hov6 & X0hov6));
assign C0hov6 = (~(S3a7z6 & Ev2nv6));
assign Rjk8v6 = (S93nv6 ? P2j7z6[0] : E1hov6);
assign Kjk8v6 = (~(L1hov6 & S1hov6));
assign S1hov6 = (~(G5j7z6[63] & Z1hov6));
assign Z1hov6 = (~(G2hov6 & N2hov6));
assign Djk8v6 = (!U2hov6);
assign U2hov6 = (M6j7z6[63] ? I3hov6 : B3hov6);
assign I3hov6 = (~(L1hov6 & P3hov6));
assign P3hov6 = (~(W3hov6 & X0hov6));
assign L1hov6 = (~(D4hov6 & K4hov6));
assign D4hov6 = (R4hov6 & Y4hov6);
assign B3hov6 = (F5hov6 & M5hov6);
assign M5hov6 = (~(T5hov6 & X0hov6));
assign F5hov6 = (~(Qkj7z6[63] | A6hov6));
assign A6hov6 = (H6hov6 & Tib7z6[63]);
assign H6hov6 = (~(Jqj7z6[72] & G5j7z6[63]));
assign Wik8v6 = (Trgov6 ? O6hov6 : Moj7z6[0]);
assign Trgov6 = (~(S93nv6 & V6hov6));
assign O6hov6 = (!C7hov6);
assign Pik8v6 = (J7hov6 & Q7hov6);
assign J7hov6 = (X7hov6 & E8hov6);
assign E8hov6 = (~(Tnzdt6 & L8hov6));
assign X7hov6 = (~(Vzvnv6 & S8hov6));
assign S8hov6 = (~(Vzbet6 & Z8hov6));
assign Z8hov6 = (~(L8hov6 & G9hov6));
assign G9hov6 = (~(N3onv6 & Ga3nv6));
assign L8hov6 = (~(N9hov6 & U9hov6));
assign U9hov6 = (Bahov6 & Iahov6);
assign Bahov6 = (~(Pahov6 & Wahov6));
assign Wahov6 = (Dbhov6 | Kbhov6);
assign N9hov6 = (Tnzdt6 & Rbhov6);
assign Rbhov6 = (~(Kbhov6 & Dbhov6));
assign Dbhov6 = (!Ybhov6);
assign Kbhov6 = (Fchov6 & Mchov6);
assign Mchov6 = (~(Tchov6 & Adhov6));
assign Fchov6 = (~(Hdhov6 & Odhov6));
assign Odhov6 = (Vdhov6 & Cehov6);
assign Vdhov6 = (~(Jehov6 & Qehov6));
assign Hdhov6 = (Moj7z6[0] & Rwl8v6);
assign Iik8v6 = (Efhov6 ? Xehov6 : Oac7z6[1]);
assign Bik8v6 = (Lfhov6 | Sfhov6);
assign Sfhov6 = (Zfhov6 & Qu1ov6);
assign Lfhov6 = (Ughov6 ? Nghov6 : Gghov6);
assign Ughov6 = (Bhhov6 & Ihhov6);
assign Ihhov6 = (~(Phhov6 & Whhov6));
assign Bhhov6 = (Dihov6 & Kihov6);
assign Dihov6 = (Rihov6 | Sb77z6);
assign Nghov6 = (Svfov6 & Lybdt6);
assign Uhk8v6 = (~(Yihov6 | Fjhov6));
assign Yihov6 = (~(Mjhov6 & Tjhov6));
assign Nhk8v6 = (~(Akhov6 & Hkhov6));
assign Hkhov6 = (~(Okhov6 & Qmj7z6[4]));
assign Okhov6 = (Vkhov6 & Lweov6);
assign Vkhov6 = (~(Jqj7z6[4] & Z3j7z6[3]));
assign Akhov6 = (Qlhov6 ? Jlhov6 : Clhov6);
assign Jlhov6 = (~(Xlhov6 & Emhov6));
assign Xlhov6 = (Lmhov6 | Lweov6);
assign Lweov6 = (!Z3j7z6[12]);
assign Clhov6 = (~(Z3j7z6[12] & Lmhov6));
assign Ghk8v6 = (~(Smhov6 & Lmhov6));
assign Lmhov6 = (~(Zmhov6 & Gnhov6));
assign Zmhov6 = (~(Kxgov6 | Z3j7z6[3]));
assign Smhov6 = (Z3j7z6[3] ? Unhov6 : Nnhov6);
assign Unhov6 = (~(Bohov6 & Iohov6));
assign Iohov6 = (~(Pohov6 & Wohov6));
assign Bohov6 = (Dphov6 & U4fov6);
assign Dphov6 = (~(Kphov6 & Rphov6));
assign Nnhov6 = (~(Wohov6 & P52nv6));
assign Zgk8v6 = (~(Yphov6 & Fqhov6));
assign Yphov6 = (Z3j7z6[0] ? Tqhov6 : Mqhov6);
assign Tqhov6 = (~(Arhov6 & Hrhov6));
assign Hrhov6 = (~(Orhov6 & Wohov6));
assign Arhov6 = (Vrhov6 & U4fov6);
assign Vrhov6 = (~(Kphov6 & Cshov6));
assign Mqhov6 = (~(Wohov6 & U42nv6));
assign Sgk8v6 = (~(Jshov6 & Qshov6));
assign Qshov6 = (~(Xshov6 & Pnfet6));
assign Xshov6 = (Ethov6 & Cveov6);
assign Ethov6 = (~(Jqj7z6[2] & Z3j7z6[0]));
assign Jshov6 = (Qlhov6 ? Sthov6 : Lthov6);
assign Sthov6 = (~(Zthov6 & Guhov6));
assign Zthov6 = (Fqhov6 | Cveov6);
assign Cveov6 = (!Z3j7z6[13]);
assign Lthov6 = (~(Z3j7z6[13] & Fqhov6));
assign Fqhov6 = (~(Nuhov6 & Uuhov6));
assign Nuhov6 = (Vzgov6 & Bvhov6);
assign Lgk8v6 = (S93nv6 ? P2j7z6[1] : Ivhov6);
assign Egk8v6 = (~(Pvhov6 & Wvhov6));
assign Wvhov6 = (~(G5j7z6[62] & Dwhov6));
assign Dwhov6 = (Kwhov6 | Rwhov6);
assign Xfk8v6 = (!Ywhov6);
assign Ywhov6 = (Oecet6 ? Mxhov6 : Fxhov6);
assign Mxhov6 = (~(Txhov6 & Ayhov6));
assign Txhov6 = (~(Hyhov6 & Oyhov6));
assign Fxhov6 = (~(Vyhov6 & Zrbet6));
assign Vyhov6 = (~(Jqj7z6[6] & Z3j7z6[8]));
assign Qfk8v6 = (~(Czhov6 & Jzhov6));
assign Jzhov6 = (~(Qzhov6 & Qmj7z6[5]));
assign Qzhov6 = (Xzhov6 & Yseov6);
assign Xzhov6 = (~(Jqj7z6[5] & Z3j7z6[7]));
assign Czhov6 = (Qlhov6 ? L0iov6 : E0iov6);
assign L0iov6 = (~(S0iov6 & Z0iov6));
assign S0iov6 = (G1iov6 | Yseov6);
assign E0iov6 = (~(Z3j7z6[15] & G1iov6));
assign Jfk8v6 = (!N1iov6);
assign N1iov6 = (Na3nv6 ? B2iov6 : U1iov6);
assign Cfk8v6 = (~(I2iov6 & P2iov6));
assign P2iov6 = (~(G5j7z6[47] & W2iov6));
assign W2iov6 = (~(D3iov6 & N2hov6));
assign Vek8v6 = (!K3iov6);
assign K3iov6 = (M6j7z6[47] ? Y3iov6 : R3iov6);
assign Y3iov6 = (~(I2iov6 & F4iov6));
assign F4iov6 = (~(M4iov6 & Z0iov6));
assign I2iov6 = (~(T4iov6 & K4hov6));
assign T4iov6 = (A5iov6 & H5iov6);
assign R3iov6 = (O5iov6 & V5iov6);
assign V5iov6 = (~(C6iov6 & Z0iov6));
assign O5iov6 = (~(Qkj7z6[47] | J6iov6));
assign J6iov6 = (Q6iov6 & Tib7z6[47]);
assign Q6iov6 = (~(Jqj7z6[56] & G5j7z6[47]));
assign Oek8v6 = (!X6iov6);
assign X6iov6 = (Na3nv6 ? L7iov6 : E7iov6);
assign Hek8v6 = (!S7iov6);
assign S7iov6 = (Na3nv6 ? G8iov6 : Z7iov6);
assign Na3nv6 = (!S93nv6);
assign S93nv6 = (~(N8iov6 & U8iov6));
assign U8iov6 = (~(B9iov6 & I9iov6));
assign I9iov6 = (P9iov6 & Nxeov6);
assign P9iov6 = (~(V5get6 & W9iov6));
assign B9iov6 = (Tnzdt6 & Daiov6);
assign Daiov6 = (~(Kaiov6 & Raiov6));
assign Raiov6 = (Yaiov6 | Ybhov6);
assign Kaiov6 = (Fbiov6 & V82nv6);
assign Fbiov6 = (~(Mbiov6 & Tbiov6));
assign Tbiov6 = (~(Ybhov6 & Yaiov6));
assign Yaiov6 = (~(Aciov6 & Hciov6));
assign Hciov6 = (~(Tchov6 & Ociov6));
assign Aciov6 = (~(Vciov6 & Moj7z6[0]));
assign Vciov6 = (Cdiov6 & Jdiov6);
assign Jdiov6 = (~(Qdiov6 & Qehov6));
assign Qehov6 = (!Tchov6);
assign Tchov6 = (Moj7z6[1] & Zyl8v6);
assign Ybhov6 = (Moj7z6[2] & H1m8v6);
assign N8iov6 = (Eugov6 & V6hov6);
assign V6hov6 = (~(Xdiov6 & Eeiov6));
assign Eeiov6 = (Leiov6 & Seiov6);
assign Seiov6 = (Zeiov6 & Gfiov6);
assign Gfiov6 = (~(E7iov6 ^ L7iov6));
assign Zeiov6 = (~(U1iov6 ^ B2iov6));
assign Leiov6 = (Nfiov6 & Ufiov6);
assign Ufiov6 = (~(Z7iov6 ^ G8iov6));
assign Nfiov6 = (Bgiov6 ^ E1hov6);
assign E1hov6 = (~(Igiov6 & Pgiov6));
assign Pgiov6 = (Wgiov6 & Dhiov6);
assign Dhiov6 = (Khiov6 & Rhiov6);
assign Rhiov6 = (~(Yhiov6 & Fiiov6));
assign Yhiov6 = (Miiov6 & Osgov6);
assign Miiov6 = (Hjiov6 ? Ajiov6 : Tiiov6);
assign Khiov6 = (~(Ojiov6 & Vjiov6));
assign Ojiov6 = (Qkiov6 ? Jkiov6 : Ckiov6);
assign Wgiov6 = (Xkiov6 & Eliov6);
assign Eliov6 = (~(Lliov6 & Sliov6));
assign Lliov6 = (Nmiov6 ? Gmiov6 : Zliov6);
assign Xkiov6 = (~(Umiov6 & Bniov6));
assign Umiov6 = (Wniov6 ? Pniov6 : Iniov6);
assign Igiov6 = (Doiov6 & Koiov6);
assign Koiov6 = (Roiov6 & Yoiov6);
assign Yoiov6 = (~(Fpiov6 & Mpiov6));
assign Fpiov6 = (Hqiov6 ? Aqiov6 : Tpiov6);
assign Aqiov6 = (Criov6 ? Vqiov6 : Oqiov6);
assign Tpiov6 = (Xriov6 ? Qriov6 : Jriov6);
assign Roiov6 = (~(Esiov6 & Lsiov6));
assign Esiov6 = (Gtiov6 ? Zsiov6 : Ssiov6);
assign Zsiov6 = (Buiov6 ? Utiov6 : Ntiov6);
assign Ssiov6 = (Wuiov6 ? Puiov6 : Iuiov6);
assign Doiov6 = (Dviov6 & Kviov6);
assign Kviov6 = (~(Rviov6 & Yviov6));
assign Yviov6 = (~(Fwiov6 & Mwiov6));
assign Mwiov6 = (Twiov6 & Axiov6);
assign Axiov6 = (Hxiov6 & Oxiov6);
assign Oxiov6 = (~(Vxiov6 & Cyiov6));
assign Vxiov6 = (Jyiov6 & Qyiov6);
assign Hxiov6 = (~(Xyiov6 & Eziov6));
assign Xyiov6 = (Zziov6 ? Sziov6 : Lziov6);
assign Twiov6 = (G0jov6 & N0jov6);
assign N0jov6 = (~(U0jov6 & B1jov6));
assign U0jov6 = (W1jov6 ? P1jov6 : I1jov6);
assign G0jov6 = (~(D2jov6 & K2jov6));
assign D2jov6 = (F3jov6 ? Y2jov6 : R2jov6);
assign Fwiov6 = (M3jov6 & T3jov6);
assign T3jov6 = (~(A4jov6 & Nxeov6));
assign M3jov6 = (H4jov6 & O4jov6);
assign O4jov6 = (~(V4jov6 & C5jov6));
assign V4jov6 = (X5jov6 ? Q5jov6 : J5jov6);
assign H4jov6 = (~(E6jov6 & L6jov6));
assign L6jov6 = (~(S6jov6 & Z6jov6));
assign Z6jov6 = (~(G7jov6 & N7jov6));
assign Dviov6 = (~(Hsgov6 & U7jov6));
assign U7jov6 = (B8jov6 | I8jov6);
assign I8jov6 = (D9jov6 ? W8jov6 : P8jov6);
assign W8jov6 = (K9jov6 & R9jov6);
assign K9jov6 = (Y9jov6 & Fajov6);
assign P8jov6 = (Abjov6 ? Tajov6 : Majov6);
assign Tajov6 = (Vbjov6 ? Objov6 : Hbjov6);
assign Majov6 = (Qcjov6 ? Jcjov6 : Ccjov6);
assign B8jov6 = (~(Xcjov6 & Edjov6));
assign Edjov6 = (~(Ldjov6 & Sdjov6));
assign Ldjov6 = (Nejov6 ? Gejov6 : Zdjov6);
assign Xcjov6 = (Uejov6 | Bfjov6);
assign Xdiov6 = (Ifjov6 & Pfjov6);
assign Pfjov6 = (Hsgov6 ^ Wfjov6);
assign Ifjov6 = (Dgjov6 & Kgjov6);
assign Kgjov6 = (Rgjov6 ^ Ivhov6);
assign Ivhov6 = (~(Ygjov6 & Fhjov6));
assign Fhjov6 = (Mhjov6 & Thjov6);
assign Thjov6 = (Aijov6 & Hijov6);
assign Hijov6 = (~(Oijov6 & Fiiov6));
assign Fiiov6 = (Vijov6 & Cjjov6);
assign Vijov6 = (Jjjov6 & Qjjov6);
assign Oijov6 = (Osgov6 & Hjiov6);
assign Aijov6 = (~(Xjjov6 & Mpiov6));
assign Xjjov6 = (Ekjov6 ? Xriov6 : Criov6);
assign Mhjov6 = (Lkjov6 & Skjov6);
assign Skjov6 = (~(Zkjov6 & Lsiov6));
assign Zkjov6 = (Gtiov6 ? Buiov6 : Wuiov6);
assign Lkjov6 = (~(Hsgov6 & Gljov6));
assign Gljov6 = (~(Nljov6 & Uljov6));
assign Uljov6 = (~(Sdjov6 & Nejov6));
assign Nljov6 = (Bmjov6 & Uejov6);
assign Uejov6 = (~(Imjov6 & D9jov6));
assign Imjov6 = (Pmjov6 & Y9jov6);
assign Bmjov6 = (~(Wmjov6 & Dnjov6));
assign Wmjov6 = (Abjov6 ? Vbjov6 : Qcjov6);
assign Ygjov6 = (Knjov6 & Rnjov6);
assign Rnjov6 = (Ynjov6 & Fojov6);
assign Fojov6 = (~(Vjiov6 & Qkiov6));
assign Vjiov6 = (Mojov6 & Tojov6);
assign Mojov6 = (~(Apjov6 | Hpjov6));
assign Ynjov6 = (~(Rviov6 & Opjov6));
assign Opjov6 = (~(Vpjov6 & Cqjov6));
assign Cqjov6 = (Jqjov6 & Qqjov6);
assign Qqjov6 = (Xqjov6 & Erjov6);
assign Erjov6 = (~(E6jov6 & Lrjov6));
assign Lrjov6 = (~(S6jov6 & Srjov6));
assign Xqjov6 = (Zrjov6 | Gsjov6);
assign Jqjov6 = (Nsjov6 & Usjov6);
assign Usjov6 = (~(Eziov6 & Zziov6));
assign Eziov6 = (Btjov6 & Itjov6);
assign Btjov6 = (Ptjov6 & Wtjov6);
assign Nsjov6 = (~(B1jov6 & W1jov6));
assign B1jov6 = (Dujov6 & Itjov6);
assign Dujov6 = (Kujov6 & Rujov6);
assign Vpjov6 = (Yujov6 & Fvjov6);
assign Yujov6 = (Mvjov6 & Tvjov6);
assign Tvjov6 = (~(K2jov6 & F3jov6));
assign Mvjov6 = (~(C5jov6 & X5jov6));
assign Knjov6 = (Awjov6 & Hwjov6);
assign Hwjov6 = (~(Sliov6 & Nmiov6));
assign Awjov6 = (~(Bniov6 & Wniov6));
assign Dgjov6 = (Osgov6 ^ Owjov6);
assign Eugov6 = (~(Kkadt6 & Sugov6));
assign Aek8v6 = (~(Vwjov6 & Cxjov6));
assign Cxjov6 = (~(Qmb7z6[8] & Jxjov6));
assign Vwjov6 = (Qxjov6 | Xxjov6);
assign Tdk8v6 = (~(Eyjov6 & Lyjov6));
assign Lyjov6 = (Syjov6 & Zyjov6);
assign Zyjov6 = (~(H02ov6 & Aw97z6));
assign Syjov6 = (Gzjov6 & Nzjov6);
assign Nzjov6 = (C12ov6 | Kajnv6);
assign Kajnv6 = (Uzjov6 & B0kov6);
assign B0kov6 = (I0kov6 & P0kov6);
assign P0kov6 = (W0kov6 & D1kov6);
assign D1kov6 = (K1kov6 & R1kov6);
assign R1kov6 = (~(vis_psp_o[8] & N32ov6));
assign K1kov6 = (~(U32ov6 & Pic7z6[8]));
assign W0kov6 = (Y1kov6 & F2kov6);
assign F2kov6 = (~(vis_msp_o[8] & P42ov6));
assign Y1kov6 = (~(vis_r12_o[8] & W42ov6));
assign I0kov6 = (M2kov6 & T2kov6);
assign T2kov6 = (A3kov6 & H3kov6);
assign H3kov6 = (~(vis_r11_o[8] & F62ov6));
assign A3kov6 = (~(vis_r10_o[8] & M62ov6));
assign M2kov6 = (O3kov6 & V3kov6);
assign V3kov6 = (~(vis_r9_o[8] & H72ov6));
assign O3kov6 = (~(vis_r8_o[8] & O72ov6));
assign Uzjov6 = (C4kov6 & J4kov6);
assign J4kov6 = (Q4kov6 & X4kov6);
assign X4kov6 = (E5kov6 & L5kov6);
assign L5kov6 = (~(vis_r7_o[8] & L92ov6));
assign E5kov6 = (~(vis_r6_o[8] & S92ov6));
assign Q4kov6 = (S5kov6 & Z5kov6);
assign Z5kov6 = (~(vis_r5_o[8] & Na2ov6));
assign S5kov6 = (~(vis_r4_o[8] & Ua2ov6));
assign C4kov6 = (G6kov6 & N6kov6);
assign N6kov6 = (U6kov6 & B7kov6);
assign B7kov6 = (~(vis_r3_o[8] & Dc2ov6));
assign U6kov6 = (~(vis_r2_o[8] & Kc2ov6));
assign G6kov6 = (I7kov6 & P7kov6);
assign P7kov6 = (~(vis_r1_o[8] & Fd2ov6));
assign I7kov6 = (~(vis_r0_o[8] & Md2ov6));
assign Gzjov6 = (~(Td2ov6 & W7kov6));
assign Eyjov6 = (D8kov6 & K8kov6);
assign K8kov6 = (~(Ve2ov6 & vis_pc_o[8]));
assign D8kov6 = (~(Fhc7z6[8] & Cf2ov6));
assign Mdk8v6 = (~(R8kov6 & Y8kov6));
assign Y8kov6 = (F9kov6 & M9kov6);
assign M9kov6 = (~(T9kov6 & C6bov6));
assign F9kov6 = (~(J6bov6 & Alf7z6[24]));
assign R8kov6 = (Aakov6 & Hakov6);
assign Hakov6 = (~(Cqf7z6[8] & E7bov6));
assign Aakov6 = (~(L0g7z6[24] & L7bov6));
assign Fdk8v6 = (~(Oakov6 & Vakov6));
assign Vakov6 = (Cbkov6 & Jbkov6);
assign Jbkov6 = (~(Sepdt6 & U8bov6));
assign Cbkov6 = (Qbkov6 & Xbkov6);
assign Xbkov6 = (~(Dsmdt6 & P9bov6));
assign Qbkov6 = (~(W9bov6 & Onf7z6[30]));
assign Oakov6 = (Eckov6 & Lckov6);
assign Lckov6 = (~(L0g7z6[30] & Rabov6));
assign Eckov6 = (Sckov6 & Zckov6);
assign Zckov6 = (~(Pvkdt6 & Mbbov6));
assign Sckov6 = (~(L0g7z6[14] & Gcmnv6));
assign Yck8v6 = (~(Gdkov6 & Ndkov6));
assign Ndkov6 = (~(Udkov6 & Bekov6));
assign Bekov6 = (~(Iekov6 & Pekov6));
assign Pekov6 = (Wekov6 | Mpe7z6[4]);
assign Iekov6 = (~(Dfkov6 & Kfkov6));
assign Gdkov6 = (Rfkov6 | Udkov6);
assign Rck8v6 = (~(Yfkov6 & Fgkov6));
assign Fgkov6 = (Mgkov6 & Tgkov6);
assign Tgkov6 = (~(Kurdt6 & U8bov6));
assign Mgkov6 = (Ahkov6 & Hhkov6);
assign Hhkov6 = (~(W8pdt6 & P9bov6));
assign Ahkov6 = (~(Onf7z6[0] & Ohkov6));
assign Yfkov6 = (Vhkov6 & Cikov6);
assign Cikov6 = (~(Bnmdt6 & Mbbov6));
assign Vhkov6 = (~(L0g7z6[0] & Rabov6));
assign Kck8v6 = (~(Jikov6 & Qikov6));
assign Qikov6 = (Xikov6 & Ejkov6);
assign Ejkov6 = (~(H02ov6 & As97z6));
assign Xikov6 = (Ljkov6 & Sjkov6);
assign Sjkov6 = (C12ov6 | Injnv6);
assign Injnv6 = (Zjkov6 & Gkkov6);
assign Gkkov6 = (Nkkov6 & Ukkov6);
assign Ukkov6 = (Blkov6 & Ilkov6);
assign Ilkov6 = (Plkov6 & Wlkov6);
assign Wlkov6 = (~(vis_psp_o[2] & N32ov6));
assign Plkov6 = (~(U32ov6 & Pic7z6[2]));
assign Blkov6 = (Dmkov6 & Kmkov6);
assign Kmkov6 = (~(vis_msp_o[2] & P42ov6));
assign Dmkov6 = (~(vis_r12_o[2] & W42ov6));
assign Nkkov6 = (Rmkov6 & Ymkov6);
assign Ymkov6 = (Fnkov6 & Mnkov6);
assign Mnkov6 = (~(vis_r11_o[2] & F62ov6));
assign Fnkov6 = (~(vis_r10_o[2] & M62ov6));
assign Rmkov6 = (Tnkov6 & Aokov6);
assign Aokov6 = (~(vis_r9_o[2] & H72ov6));
assign Tnkov6 = (~(vis_r8_o[2] & O72ov6));
assign Zjkov6 = (Hokov6 & Ookov6);
assign Ookov6 = (Vokov6 & Cpkov6);
assign Cpkov6 = (Jpkov6 & Qpkov6);
assign Qpkov6 = (~(vis_r7_o[2] & L92ov6));
assign Jpkov6 = (~(vis_r6_o[2] & S92ov6));
assign Vokov6 = (Xpkov6 & Eqkov6);
assign Eqkov6 = (~(vis_r5_o[2] & Na2ov6));
assign Xpkov6 = (~(vis_r4_o[2] & Ua2ov6));
assign Hokov6 = (Lqkov6 & Sqkov6);
assign Sqkov6 = (Zqkov6 & Grkov6);
assign Grkov6 = (~(vis_r3_o[2] & Dc2ov6));
assign Zqkov6 = (~(vis_r2_o[2] & Kc2ov6));
assign Lqkov6 = (Nrkov6 & Urkov6);
assign Urkov6 = (~(vis_r1_o[2] & Fd2ov6));
assign Nrkov6 = (~(vis_r0_o[2] & Md2ov6));
assign Ljkov6 = (~(Td2ov6 & Bskov6));
assign Jikov6 = (Iskov6 & Pskov6);
assign Pskov6 = (~(Ve2ov6 & vis_pc_o[2]));
assign Iskov6 = (~(E3c7z6[2] & Cf2ov6));
assign Dck8v6 = (~(Wskov6 & Dtkov6));
assign Dtkov6 = (Ktkov6 & Rtkov6);
assign Rtkov6 = (~(Iv3ov6 & C6bov6));
assign Ktkov6 = (~(J6bov6 & Alf7z6[30]));
assign Wskov6 = (Ytkov6 & Fukov6);
assign Fukov6 = (~(Cqf7z6[14] & E7bov6));
assign Ytkov6 = (~(L0g7z6[30] & L7bov6));
assign Wbk8v6 = (~(Mukov6 & Tukov6));
assign Tukov6 = (Avkov6 & Hvkov6);
assign Hvkov6 = (~(Qhpdt6 & U8bov6));
assign Avkov6 = (Ovkov6 & Vvkov6);
assign Vvkov6 = (~(Cvmdt6 & P9bov6));
assign Ovkov6 = (~(W9bov6 & Onf7z6[29]));
assign Mukov6 = (Cwkov6 & Jwkov6);
assign Jwkov6 = (~(L0g7z6[29] & Rabov6));
assign Cwkov6 = (Qwkov6 & Xwkov6);
assign Xwkov6 = (~(Sxkdt6 & Mbbov6));
assign Qwkov6 = (~(L0g7z6[13] & Gcmnv6));
assign Pbk8v6 = (~(Exkov6 & Lxkov6));
assign Lxkov6 = (Sxkov6 & Zxkov6);
assign Zxkov6 = (~(H02ov6 & Iw97z6));
assign Sxkov6 = (Gykov6 & Nykov6);
assign Nykov6 = (C12ov6 | Wgjnv6);
assign Wgjnv6 = (Uykov6 & Bzkov6);
assign Bzkov6 = (Izkov6 & Pzkov6);
assign Pzkov6 = (Wzkov6 & D0lov6);
assign D0lov6 = (K0lov6 & R0lov6);
assign R0lov6 = (~(vis_psp_o[4] & N32ov6));
assign K0lov6 = (~(U32ov6 & Pic7z6[4]));
assign Wzkov6 = (Y0lov6 & F1lov6);
assign F1lov6 = (~(vis_msp_o[4] & P42ov6));
assign Y0lov6 = (~(vis_r12_o[4] & W42ov6));
assign Izkov6 = (M1lov6 & T1lov6);
assign T1lov6 = (A2lov6 & H2lov6);
assign H2lov6 = (~(vis_r11_o[4] & F62ov6));
assign A2lov6 = (~(vis_r10_o[4] & M62ov6));
assign M1lov6 = (O2lov6 & V2lov6);
assign V2lov6 = (~(vis_r9_o[4] & H72ov6));
assign O2lov6 = (~(vis_r8_o[4] & O72ov6));
assign Uykov6 = (C3lov6 & J3lov6);
assign J3lov6 = (Q3lov6 & X3lov6);
assign X3lov6 = (E4lov6 & L4lov6);
assign L4lov6 = (~(vis_r7_o[4] & L92ov6));
assign E4lov6 = (~(vis_r6_o[4] & S92ov6));
assign Q3lov6 = (S4lov6 & Z4lov6);
assign Z4lov6 = (~(vis_r5_o[4] & Na2ov6));
assign S4lov6 = (~(vis_r4_o[4] & Ua2ov6));
assign C3lov6 = (G5lov6 & N5lov6);
assign N5lov6 = (U5lov6 & B6lov6);
assign B6lov6 = (~(vis_r3_o[4] & Dc2ov6));
assign U5lov6 = (~(vis_r2_o[4] & Kc2ov6));
assign G5lov6 = (I6lov6 & P6lov6);
assign P6lov6 = (~(vis_r1_o[4] & Fd2ov6));
assign I6lov6 = (~(vis_r0_o[4] & Md2ov6));
assign Gykov6 = (~(Td2ov6 & W6lov6));
assign Exkov6 = (D7lov6 & K7lov6);
assign K7lov6 = (~(Ve2ov6 & vis_pc_o[4]));
assign D7lov6 = (~(E3c7z6[4] & Cf2ov6));
assign Ibk8v6 = (~(Wpvnv6 & R7lov6));
assign R7lov6 = (~(Y7lov6 & F02nv6));
assign Y7lov6 = (~(F8lov6 & M8lov6));
assign F8lov6 = (S2onv6 & C0wnv6);
assign Bbk8v6 = (~(T8lov6 & A9lov6));
assign A9lov6 = (~(H9lov6 & X6eet6));
assign H9lov6 = (~(Ldo7v6 | Kdadt6));
assign Uak8v6 = (Kdadt6 ? Bpvnv6 : O9lov6);
assign Bpvnv6 = (V9lov6 | Ldo7v6);
assign O9lov6 = (Calov6 & O5a7z6);
assign Calov6 = (Ztaov6 & Gvvnv6);
assign Nak8v6 = (Jalov6 & Qalov6);
assign Qalov6 = (~(Xalov6 & Eblov6));
assign Eblov6 = (~(Hryet6 & Lblov6));
assign Xalov6 = (~(Sblov6 & Zblov6));
assign Gak8v6 = (~(Gclov6 & Nclov6));
assign Nclov6 = (~(Hl9ov6 & Uclov6));
assign Gclov6 = (~(Dq9ov6 & Ewyet6));
assign Z9k8v6 = (Bdlov6 | A497z6);
assign S9k8v6 = (~(Bdlov6 & Idlov6));
assign Idlov6 = (~(Pdlov6 & Ja1ft6));
assign Bdlov6 = (~(Wdlov6 & Delov6));
assign Delov6 = (~(Kelov6 & Relov6));
assign Kelov6 = (~(Yelov6 | Fflov6));
assign L9k8v6 = (Mflov6 & Kb77z6);
assign Mflov6 = (Aglov6 ? Frzet6 : Tflov6);
assign Tflov6 = (I6oet6 & Hglov6);
assign Hglov6 = (~(Oglov6 & Vglov6));
assign Vglov6 = (Chlov6 & Jhlov6);
assign Jhlov6 = (~(Dtm7z6[3] & Qhlov6));
assign Chlov6 = (~(Dtm7z6[2] & Xhlov6));
assign Oglov6 = (Eilov6 & Lilov6);
assign Lilov6 = (~(Dtm7z6[0] & HRESPD[0]));
assign Eilov6 = (~(Dtm7z6[1] & HRESPS[0]));
assign E9k8v6 = (Silov6 ? Zdh7v6 : Blzet6);
assign X8k8v6 = (~(Zilov6 & Gjlov6));
assign Gjlov6 = (~(Njlov6 & Ujlov6));
assign Zilov6 = (~(Bklov6 & Pvj7z6[0]));
assign Q8k8v6 = (Pklov6 ? Iklov6 : Hfm7z6[25]);
assign J8k8v6 = (Pb9ov6 ? D6c7z6[3] : Wklov6);
assign Wklov6 = (~(Dllov6 & Kllov6));
assign Kllov6 = (Rllov6 & Yllov6);
assign Yllov6 = (~(Yc9ov6 & Fmlov6));
assign Rllov6 = (~(Md9ov6 & Mmlov6));
assign Dllov6 = (Tmlov6 & Anlov6);
assign Anlov6 = (~(Oe9ov6 & Hnlov6));
assign Tmlov6 = (~(Cf9ov6 & Onlov6));
assign C8k8v6 = (~(Vnlov6 & Colov6));
assign Colov6 = (Jolov6 | Qolov6);
assign Vnlov6 = (Xolov6 & Eplov6);
assign Eplov6 = (~(Lplov6 & Splov6));
assign Splov6 = (Zplov6 & Gqlov6);
assign Gqlov6 = (~(Nqlov6 | Qmb7z6[6]));
assign Nqlov6 = (Qmb7z6[7] | Qmb7z6[8]);
assign Zplov6 = (~(Qmb7z6[4] | Qmb7z6[5]));
assign Lplov6 = (Uqlov6 & Brlov6);
assign Brlov6 = (~(Irlov6 | Qmb7z6[1]));
assign Irlov6 = (Qmb7z6[2] | Qmb7z6[3]);
assign Uqlov6 = (~(Prlov6 | Qmb7z6[0]));
assign Prlov6 = (~(Wrlov6 | Lcadt6));
assign Xolov6 = (~(Dslov6 & Kslov6));
assign Dslov6 = (~(Rslov6 | Lcadt6));
assign V7k8v6 = (!Yslov6);
assign Yslov6 = (O5a7z6 ? Mtlov6 : Ftlov6);
assign Mtlov6 = (~(Ttlov6 & Aulov6));
assign Ttlov6 = (Hulov6 & Oulov6);
assign Oulov6 = (~(Rslov6 ^ Vulov6));
assign Vulov6 = (Cvlov6 & Jvlov6);
assign Jvlov6 = (Qvlov6 & Xvlov6);
assign Xvlov6 = (Ewlov6 & Lwlov6);
assign Ewlov6 = (~(Swlov6 | Zwlov6));
assign Qvlov6 = (Gxlov6 & Nxlov6);
assign Cvlov6 = (Uxlov6 & Bylov6);
assign Bylov6 = (Iylov6 & Pylov6);
assign Uxlov6 = (Wylov6 & Dzlov6);
assign O7k8v6 = (~(Kzlov6 & Rzlov6));
assign Rzlov6 = (~(Yzlov6 & F0mov6));
assign F0mov6 = (Svfov6 & Vs9ov6);
assign Yzlov6 = (L2gdt6 & M0mov6);
assign Kzlov6 = (~(T0mov6 & A1mov6));
assign A1mov6 = (~(H1mov6 & O1mov6));
assign O1mov6 = (V1mov6 & Gpfov6);
assign Gpfov6 = (C2mov6 & J2mov6);
assign J2mov6 = (~(Q2mov6 & X2mov6));
assign C2mov6 = (E3mov6 & L3mov6);
assign L3mov6 = (~(S3mov6 & Z3mov6));
assign S3mov6 = (G4mov6 ? Zec7z6[1] : Zec7z6[17]);
assign E3mov6 = (~(N4mov6 & Ohe7z6[1]));
assign H1mov6 = (U4mov6 & B5mov6);
assign T0mov6 = (~(I5mov6 & M0mov6));
assign I5mov6 = (Svfov6 & P5mov6);
assign Svfov6 = (!Qu1ov6);
assign H7k8v6 = (C1onv6 & W5mov6);
assign C1onv6 = (~(Fjhov6 | D6mov6));
assign A7k8v6 = (Tznnv6 & W5mov6);
assign W5mov6 = (~(K6mov6 & R6mov6));
assign R6mov6 = (~(S2onv6 & Geh7v6));
assign Tznnv6 = (~(Fjhov6 | Y6mov6));
assign Fjhov6 = (~(F7mov6 & G3onv6));
assign F7mov6 = (~(M7mov6 | T7mov6));
assign T6k8v6 = (A8mov6 & H8mov6);
assign H8mov6 = (~(O8mov6 & V8mov6));
assign V8mov6 = (~(Loddt6 & C9mov6));
assign O8mov6 = (~(J9mov6 | Pqddt6));
assign M6k8v6 = (Pqddt6 | Q9mov6);
assign Q9mov6 = (X9mov6 & Eamov6);
assign Eamov6 = (~(J9mov6 | C9mov6));
assign J9mov6 = (A8mov6 & Lamov6);
assign X9mov6 = (Loddt6 & Samov6);
assign F6k8v6 = (~(Zamov6 & Gbmov6));
assign Gbmov6 = (~(Dheet6 & Nbmov6));
assign Y5k8v6 = (Ubmov6 ? D62nv6 : Qteet6);
assign Ubmov6 = (~(Bcmov6 | Dheet6));
assign R5k8v6 = (~(Mdonv6 & Icmov6));
assign Icmov6 = (~(Pcmov6 & Wcmov6));
assign Pcmov6 = (Aeonv6 & B2jnv6);
assign K5k8v6 = (!Ddmov6);
assign Ddmov6 = (Kdmov6 ? Y497z6 : Jfonv6);
assign D5k8v6 = (Mdonv6 ? Rj9ov6 : Qboet6);
assign W4k8v6 = (~(Sh2nv6 | Rdmov6));
assign P4k8v6 = (~(Ydmov6 & Femov6));
assign Femov6 = (~(Memov6 & Temov6));
assign Temov6 = (Afmov6 & Hfmov6);
assign Hfmov6 = (Ofmov6 & Cmm7z6[9]);
assign Ofmov6 = (Cmm7z6[6] & Cmm7z6[8]);
assign Afmov6 = (Vfmov6 & Cmm7z6[7]);
assign Memov6 = (Cgmov6 & Jgmov6);
assign Jgmov6 = (Cmm7z6[4] & Cmm7z6[5]);
assign Cgmov6 = (Yefnv6 & Cmm7z6[3]);
assign Ydmov6 = (~(Ex7et6 & Vrinv6));
assign I4k8v6 = (!Qgmov6);
assign Qgmov6 = (Vfmov6 ? Ehmov6 : Xgmov6);
assign Ehmov6 = (~(Evadt6 & Lgonv6));
assign B4k8v6 = (W13et6 | Vfmov6);
assign U3k8v6 = (Shmov6 ? Ow2et6 : Lhmov6);
assign N3k8v6 = (Shmov6 ? Kih7z6[1] : Cmm7z6[1]);
assign G3k8v6 = (Shmov6 ? Kih7z6[0] : Cmm7z6[0]);
assign Z2k8v6 = (!Zhmov6);
assign Zhmov6 = (Vfmov6 ? Nimov6 : Gimov6);
assign Nimov6 = (~(M43et6 & K73et6));
assign S2k8v6 = (Uimov6 ? Xmtet6 : Cmm7z6[1]);
assign L2k8v6 = (Uimov6 ? Yotet6 : Cmm7z6[0]);
assign E2k8v6 = (Bjmov6 & Ypinv6);
assign Bjmov6 = (~(Ijmov6 & Pjmov6));
assign Pjmov6 = (~(W13et6 & Wjmov6));
assign Wjmov6 = (~(Dkmov6 & Kkmov6));
assign Kkmov6 = (~(Rkmov6 & Ykmov6));
assign Ykmov6 = (Flmov6 & Mlmov6);
assign Rkmov6 = (A0onv6 & Tlmov6);
assign Dkmov6 = (~(Ammov6 & Gimov6));
assign Ammov6 = (~(Hmmov6 & Ommov6));
assign Ommov6 = (~(A0onv6 & Whhov6));
assign X1k8v6 = (~(Vmmov6 & Cnmov6));
assign Cnmov6 = (~(Jnmov6 & Kgbdt6));
assign Jnmov6 = (Qnmov6 & Xnmov6);
assign Qnmov6 = (~(O5a7z6 & Eomov6));
assign Eomov6 = (~(Lomov6 & Somov6));
assign Lomov6 = (Zomov6 & Gpmov6);
assign Zomov6 = (~(Npmov6 & Ijmov6));
assign Npmov6 = (~(Upmov6 & Bqmov6));
assign Upmov6 = (Flmov6 & Iqmov6);
assign Vmmov6 = (~(Pqmov6 & Wqmov6));
assign Wqmov6 = (~(Drmov6 & Krmov6));
assign Krmov6 = (~(Rrmov6 & Yrmov6));
assign Yrmov6 = (U1jnv6 & Fsmov6);
assign Rrmov6 = (Msmov6 & N1jnv6);
assign Drmov6 = (~(Tsmov6 & Atmov6));
assign Tsmov6 = (Ypinv6 & Ijmov6);
assign Pqmov6 = (~(Htmov6 | Nhonv6));
assign Q1k8v6 = (~(Otmov6 & Vtmov6));
assign Vtmov6 = (Cumov6 & Jumov6);
assign Jumov6 = (~(Qumov6 & Xumov6));
assign Cumov6 = (Evmov6 & Lvmov6);
assign Lvmov6 = (Svmov6 | Bvaov6);
assign Evmov6 = (~(Zvmov6 & Gwmov6));
assign Otmov6 = (Nwmov6 & Uwmov6);
assign Uwmov6 = (~(Bxmov6 & Ixmov6));
assign Nwmov6 = (~(Nnaov6 & Pxmov6));
assign J1k8v6 = (~(Wxmov6 & Dymov6));
assign Dymov6 = (Kymov6 & 1'b1);
assign Kymov6 = (Rymov6 & Yymov6);
assign Yymov6 = (Svmov6 | Zmaov6);
assign Zmaov6 = (!Fzmov6);
assign Rymov6 = (~(Zvmov6 & Mzmov6));
assign Wxmov6 = (Tzmov6 & A0nov6);
assign A0nov6 = (~(Bxmov6 & H0nov6));
assign Tzmov6 = (~(Nnaov6 & Xlaov6));
assign C1k8v6 = (~(O0nov6 & V0nov6));
assign V0nov6 = (C1nov6 & J1nov6);
assign J1nov6 = (~(Qumov6 & Xlaov6));
assign C1nov6 = (Q1nov6 & X1nov6);
assign X1nov6 = (Svmov6 | Fqaov6);
assign Fqaov6 = (!E2nov6);
assign Q1nov6 = (~(Zvmov6 & L2nov6));
assign O0nov6 = (S2nov6 & Z2nov6);
assign Z2nov6 = (~(Bxmov6 & G3nov6));
assign S2nov6 = (~(Nnaov6 & Kpaov6));
assign V0k8v6 = (~(N3nov6 & U3nov6));
assign U3nov6 = (B4nov6 & I4nov6);
assign I4nov6 = (~(Qumov6 & Kpaov6));
assign Qumov6 = (P4nov6 & Ywaov6);
assign P4nov6 = (Fxaov6 & W4nov6);
assign B4nov6 = (D5nov6 & K5nov6);
assign K5nov6 = (Svmov6 | Ivaov6);
assign Svmov6 = (~(R5nov6 & Staov6));
assign R5nov6 = (Ztaov6 & W4nov6);
assign D5nov6 = (~(Zvmov6 & Y5nov6));
assign Zvmov6 = (W4nov6 & F6nov6);
assign F6nov6 = (~(M6nov6 & Txaov6));
assign M6nov6 = (Etaov6 & Ayaov6);
assign Etaov6 = (~(Xtvnv6 & Lyknv6));
assign N3nov6 = (T6nov6 & A7nov6);
assign A7nov6 = (~(Bxmov6 & H7nov6));
assign Bxmov6 = (O7nov6 & W4nov6);
assign O7nov6 = (~(V7nov6 & C8nov6));
assign V7nov6 = (J8nov6 & Xzaov6);
assign Xzaov6 = (~(Q8nov6 & X8nov6));
assign X8nov6 = (~(Tnzdt6 & E9nov6));
assign Q8nov6 = (L9nov6 & Bfo7v6);
assign T6nov6 = (~(Nnaov6 & Xumov6));
assign O0k8v6 = (~(Vs9ov6 & S9nov6));
assign S9nov6 = (~(Zhbdt6 & Rihov6));
assign H0k8v6 = (~(V1mov6 & Z9nov6));
assign Z9nov6 = (~(Upfov6 & Ohe7z6[3]));
assign V1mov6 = (Ganov6 & Nanov6);
assign Nanov6 = (~(Uanov6 & X2mov6));
assign Ganov6 = (Bbnov6 & Ibnov6);
assign Ibnov6 = (~(Pbnov6 & Z3mov6));
assign Pbnov6 = (G4mov6 ? Zec7z6[2] : Zec7z6[18]);
assign Bbnov6 = (~(N4mov6 & Ohe7z6[2]));
assign A0k8v6 = (~(G4mov6 & Wbnov6));
assign Wbnov6 = (~(Knbdt6 & Dcnov6));
assign Tzj8v6 = (~(Kcnov6 & Rcnov6));
assign Rcnov6 = (Ycnov6 | Hs9ov6);
assign Kcnov6 = (~(I9e7z6[2] & Dcnov6));
assign Mzj8v6 = (Mdnov6 ? Nmadt6 : Fdnov6);
assign Mdnov6 = (Tdnov6 & Dqgov6);
assign Dqgov6 = (~(Rkfov6 & Cgfov6));
assign Tdnov6 = (~(Kqgov6 & Aenov6));
assign Aenov6 = (I9e7z6[2] | Ibe7z6[0]);
assign Kqgov6 = (Shfov6 & Cgfov6);
assign Cgfov6 = (Ib3nv6 | Henov6);
assign Ib3nv6 = (Oenov6 & Lugov6);
assign Lugov6 = (!X83nv6);
assign X83nv6 = (Oxfet6 & SLEEPHOLDACKn);
assign Oxfet6 = (!Jg2nv6);
assign Oenov6 = (~(Venov6 & Cfnov6));
assign Cfnov6 = (~(Sh2nv6 & Qg2nv6));
assign Fdnov6 = (~(Jfnov6 & Qfnov6));
assign Qfnov6 = (~(Rkfov6 & Swlov6));
assign Fzj8v6 = (~(Xfnov6 | Tnzdt6));
assign Yyj8v6 = (Lgnov6 ? Tkbdt6 : Egnov6);
assign Lgnov6 = (Sgnov6 & Lhfov6);
assign Sgnov6 = (!Zgnov6);
assign Egnov6 = (Ibe7z6[4] ? E3c7z6[0] : Zfhov6);
assign Ryj8v6 = (Wj1ov6 ? Ghnov6 : Fsc7z6[1]);
assign Kyj8v6 = (~(Nhnov6 & Uhnov6));
assign Nhnov6 = (~(Ztcdt6 & M4xnv6));
assign Dyj8v6 = (Binov6 & F4xnv6);
assign Binov6 = (Crcdt6 | Wj1ov6);
assign Wxj8v6 = (~(T8ddt6 ^ Iinov6));
assign Iinov6 = (T8ddt6 ? Uhnov6 : Ldo7v6);
assign Uhnov6 = (~(N8xnv6 & Am1ov6));
assign Pxj8v6 = (Qp38v6 | Pinov6);
assign Pinov6 = (Winov6 & Djnov6);
assign Djnov6 = (Kjnov6 & Pj1ov6);
assign Kjnov6 = (~(Iladt6 & J21ov6));
assign Winov6 = (Rjnov6 & Sgcdt6);
assign Ixj8v6 = (Fknov6 ? Yjnov6 : Cgc7z6[1]);
assign Yjnov6 = (~(Mknov6 & Tknov6));
assign Tknov6 = (Alnov6 & Hlnov6);
assign Hlnov6 = (Olnov6 & Nx0ov6);
assign Alnov6 = (Vlnov6 & Cmnov6);
assign Cmnov6 = (~(Jmnov6 & Qg2nv6));
assign Jmnov6 = (Qmnov6 | Xmnov6);
assign Vlnov6 = (~(Ennov6 & J21ov6));
assign Mknov6 = (Lnnov6 & Snnov6);
assign Snnov6 = (~(Znnov6 & Gonov6));
assign Lnnov6 = (Nonov6 & Uonov6);
assign Uonov6 = (~(Bpnov6 & Rgo7v6));
assign Nonov6 = (~(Ipnov6 & Pj1ov6));
assign Bxj8v6 = (~(Ldbdt6 ^ Ppnov6));
assign Ppnov6 = (Ldbdt6 ? Wpnov6 : Dxvnv6);
assign Wpnov6 = (~(Wrlov6 | Dqnov6));
assign Uwj8v6 = (~(Kqnov6 & Rqnov6));
assign Rqnov6 = (~(Yqnov6 & Frnov6));
assign Yqnov6 = (M0edt6 & Mrnov6);
assign Kqnov6 = (~(Trnov6 & Asnov6));
assign Asnov6 = (~(Hsnov6 & Osnov6));
assign Osnov6 = (~(Vsnov6 & Ctnov6));
assign Hsnov6 = (~(Jtnov6 & Qtnov6));
assign Nwj8v6 = (~(Xnfov6 & T0fov6));
assign T0fov6 = (SLEEPHOLDACKn | SLEEPHOLDREQn);
assign Xnfov6 = (~(Xtnov6 & SLEEPING));
assign Xtnov6 = (~(M0fov6 | SLEEPHOLDREQn));
assign M0fov6 = (Eunov6 & Lunov6);
assign Eunov6 = (Pyeov6 & Sunov6);
assign Zvj8v6 = (Fknov6 ? Zunov6 : Cgc7z6[0]);
assign Zunov6 = (~(Gvnov6 & Nvnov6));
assign Nvnov6 = (Uvnov6 & Bwnov6);
assign Uvnov6 = (P51ov6 & Iwnov6);
assign Gvnov6 = (Pwnov6 & Wwnov6);
assign Wwnov6 = (Dxnov6 & Kxnov6);
assign Kxnov6 = (~(Xmnov6 & Qg2nv6));
assign Dxnov6 = (~(Rxnov6 & IFLUSH));
assign Pwnov6 = (Yxnov6 & Fynov6);
assign Fynov6 = (~(Bpnov6 & Gonov6));
assign Svj8v6 = (Fknov6 ? Mynov6 : Cgc7z6[2]);
assign Mynov6 = (~(Tynov6 & Aznov6));
assign Aznov6 = (Hznov6 & Olnov6);
assign Olnov6 = (~(Ennov6 & Oznov6));
assign Hznov6 = (~(Gonov6 & Vznov6));
assign Vznov6 = (~(Hu0ov6 & C0oov6));
assign C0oov6 = (~(Bpnov6 & Aiadt6));
assign Tynov6 = (Yxnov6 & J0oov6);
assign J0oov6 = (~(Q0oov6 & Pj1ov6));
assign Q0oov6 = (~(X0oov6 & P51ov6));
assign Yxnov6 = (E1oov6 & L1oov6);
assign L1oov6 = (S1oov6 | Tnzdt6);
assign E1oov6 = (~(Z1oov6 & G2oov6));
assign Lvj8v6 = (Fknov6 ? N2oov6 : Cgc7z6[3]);
assign Fknov6 = (~(U2oov6 & B3oov6));
assign B3oov6 = (I3oov6 & P3oov6);
assign P3oov6 = (W3oov6 & D4oov6);
assign D4oov6 = (K4oov6 & Iwnov6);
assign K4oov6 = (~(R4oov6 & Bpnov6));
assign R4oov6 = (Ldo7v6 & Y4oov6);
assign Y4oov6 = (~(Dxvnv6 & F5oov6));
assign F5oov6 = (~(O5a7z6 & Tnzdt6));
assign W3oov6 = (M5oov6 & T5oov6);
assign T5oov6 = (~(A6oov6 & H6oov6));
assign H6oov6 = (~(Iladt6 & X0wnv6));
assign M5oov6 = (~(Xmnov6 & O6oov6));
assign O6oov6 = (~(Qg2nv6 & V6oov6));
assign V6oov6 = (~(K3jnv6 & Sh2nv6));
assign Xmnov6 = (!C7oov6);
assign I3oov6 = (J7oov6 & Q7oov6);
assign Q7oov6 = (~(N8xnv6 & X7oov6));
assign X7oov6 = (~(E8oov6 & L8oov6));
assign E8oov6 = (S8oov6 & Z8oov6);
assign S8oov6 = (~(G9oov6 & Pj1ov6));
assign G9oov6 = (Qmnov6 | N9oov6);
assign J7oov6 = (U9oov6 & Baoov6);
assign Baoov6 = (~(J21ov6 & Iaoov6));
assign Iaoov6 = (~(Ennov6 & Paoov6));
assign Paoov6 = (~(Waoov6 & H11ov6));
assign Waoov6 = (~(Dboov6 | Sgcdt6));
assign U9oov6 = (~(Kboov6 & Rboov6));
assign Rboov6 = (~(Gonov6 & Qv0ov6));
assign U2oov6 = (Yboov6 & Fcoov6);
assign Fcoov6 = (Mcoov6 & Tcoov6);
assign Tcoov6 = (Pj1ov6 | L8oov6);
assign Mcoov6 = (Adoov6 & Hdoov6);
assign Hdoov6 = (~(Odoov6 & Wrlov6));
assign Wrlov6 = (!Vsgov6);
assign Adoov6 = (Venov6 | Vdoov6);
assign Yboov6 = (Ceoov6 & Jeoov6);
assign Ceoov6 = (Rjnov6 & Qeoov6);
assign Qeoov6 = (~(Sa2nv6 & Z1oov6));
assign Rjnov6 = (Xeoov6 & P51ov6);
assign Xeoov6 = (~(Efoov6 & Lfoov6));
assign Lfoov6 = (~(Dboov6 | Sfoov6));
assign Dboov6 = (Zfoov6 & Somov6);
assign Somov6 = (~(Ggoov6 & Dwb7z6[1]));
assign Zfoov6 = (Ngoov6 & Ugoov6);
assign Ugoov6 = (~(Bhoov6 & Ihoov6));
assign Ihoov6 = (~(Phoov6 & Whoov6));
assign Whoov6 = (~(Dioov6 & Kioov6));
assign Phoov6 = (~(Fxaov6 & Uvvnv6));
assign Ngoov6 = (~(Rioov6 & Yioov6));
assign Efoov6 = (J21ov6 & H11ov6);
assign N2oov6 = (~(Fjoov6 & Mjoov6));
assign Mjoov6 = (Tjoov6 & C7oov6);
assign C7oov6 = (~(Akoov6 & Cgc7z6[3]));
assign Akoov6 = (Cgc7z6[0] & Cgc7z6[2]);
assign Tjoov6 = (Hu0ov6 & Hkoov6);
assign Fjoov6 = (Vdoov6 & Jeoov6);
assign Jeoov6 = (Okoov6 & Vkoov6);
assign Vkoov6 = (~(Iladt6 & Z1oov6));
assign Okoov6 = (Cloov6 & Jloov6);
assign Jloov6 = (Qg2nv6 | S1oov6);
assign S1oov6 = (~(Qmnov6 | Odoov6));
assign Odoov6 = (Qloov6 & Cgc7z6[0]);
assign Cloov6 = (Z8oov6 | Ennov6);
assign Ennov6 = (G2oov6 & Pj1ov6);
assign Vdoov6 = (X6xnv6 & Xloov6);
assign Evj8v6 = (Wj1ov6 ? Emoov6 : Fsc7z6[0]);
assign Xuj8v6 = (~(Lmoov6 & Smoov6));
assign Smoov6 = (~(N8xnv6 & Emoov6));
assign Lmoov6 = (~(Ywcdt6 & M4xnv6));
assign Quj8v6 = (Zmoov6 & Gnoov6);
assign Gnoov6 = (Nnoov6 & Unoov6);
assign Unoov6 = (Booov6 & Nx0ov6);
assign Booov6 = (Iooov6 & G2oov6);
assign Nnoov6 = (~(Sugov6 | S1wnv6));
assign Zmoov6 = (Pooov6 & Wooov6);
assign Wooov6 = (Dpoov6 & Gpmov6);
assign Dpoov6 = (V5ddt6 | IFLUSH);
assign Juj8v6 = (Rpoov6 ? P6d7z6[1] : Kpoov6);
assign Kpoov6 = (Ypoov6 & P6d7z6[0]);
assign Cuj8v6 = (As9ov6 ? L9d7z6[3] : Ujnet6);
assign Vtj8v6 = (Rpoov6 ? P6d7z6[0] : Fqoov6);
assign Fqoov6 = (Mqoov6 | P6d7z6[2]);
assign Otj8v6 = (Tqoov6 ? L9d7z6[0] : Tr9ov6);
assign Htj8v6 = (Tqoov6 ? L9d7z6[1] : Ujnet6);
assign Atj8v6 = (Rpoov6 ? P6d7z6[2] : Aroov6);
assign Rpoov6 = (Hroov6 & Ij1ov6);
assign Hroov6 = (~(Mqoov6 & Oroov6));
assign Oroov6 = (~(Vroov6 & P6d7z6[0]));
assign Mqoov6 = (!Ypoov6);
assign Aroov6 = (Ypoov6 & P6d7z6[1]);
assign Ypoov6 = (Vroov6 & Csoov6);
assign Csoov6 = (Jsoov6 & Qsoov6);
assign Vroov6 = (D61ov6 & Iwnov6);
assign Tsj8v6 = (~(Xsoov6 & Etoov6));
assign Etoov6 = (~(Tr9ov6 & H5xnv6));
assign Xsoov6 = (~(O5xnv6 & L9d7z6[4]));
assign Msj8v6 = (~(Ltoov6 & Stoov6));
assign Stoov6 = (Ztoov6 & Guoov6);
assign Guoov6 = (Nuoov6 & Uuoov6);
assign Uuoov6 = (~(Bvoov6 & D9o7v6));
assign Nuoov6 = (Ivoov6 & Pvoov6);
assign Pvoov6 = (~(Byc7z6[16] & Wvoov6));
assign Ivoov6 = (~(Dwoov6 & N6znv6));
assign Ztoov6 = (Kwoov6 & Rwoov6);
assign Rwoov6 = (~(X91ov6 & Ke48v6));
assign Kwoov6 = (~(Ea1ov6 & Nvs7v6));
assign Ltoov6 = (Ywoov6 & Fxoov6);
assign Fxoov6 = (Mxoov6 & Txoov6);
assign Txoov6 = (~(Nb1ov6 & De48v6));
assign Mxoov6 = (~(Byc7z6[0] & Ub1ov6));
assign Ywoov6 = (Ayoov6 & Hyoov6);
assign Hyoov6 = (~(Pc1ov6 & Kaxnv6));
assign Ayoov6 = (~(Zec7z6[0] & Wc1ov6));
assign Fsj8v6 = (~(Oyoov6 & Vyoov6));
assign Vyoov6 = (Czoov6 & Jzoov6);
assign Jzoov6 = (Qzoov6 & Xzoov6);
assign Xzoov6 = (~(A81ov6 & Rl48v6));
assign Qzoov6 = (E0pov6 & L0pov6);
assign L0pov6 = (~(Byc7z6[14] & V81ov6));
assign E0pov6 = (~(C91ov6 & Geynv6));
assign Czoov6 = (S0pov6 & Z0pov6);
assign Z0pov6 = (~(X91ov6 & Gos7v6));
assign S0pov6 = (~(Ea1ov6 & R9o7v6));
assign Oyoov6 = (G1pov6 & N1pov6);
assign N1pov6 = (U1pov6 & B2pov6);
assign B2pov6 = (~(Nb1ov6 & K9o7v6));
assign U1pov6 = (~(Byc7z6[30] & Ub1ov6));
assign G1pov6 = (I2pov6 & P2pov6);
assign P2pov6 = (~(Pc1ov6 & Zexnv6));
assign I2pov6 = (~(Zec7z6[30] & Wc1ov6));
assign Yrj8v6 = (~(W2pov6 & D3pov6));
assign D3pov6 = (K3pov6 & R3pov6);
assign R3pov6 = (Y3pov6 & F4pov6);
assign F4pov6 = (~(A81ov6 & Kl48v6));
assign Y3pov6 = (M4pov6 & T4pov6);
assign T4pov6 = (~(Byc7z6[13] & V81ov6));
assign M4pov6 = (~(C91ov6 & Viynv6));
assign K3pov6 = (A5pov6 & H5pov6);
assign H5pov6 = (~(X91ov6 & Uos7v6));
assign A5pov6 = (~(Ea1ov6 & Dl48v6));
assign W2pov6 = (O5pov6 & V5pov6);
assign V5pov6 = (C6pov6 & J6pov6);
assign J6pov6 = (~(Nb1ov6 & Nos7v6));
assign C6pov6 = (~(Byc7z6[29] & Ub1ov6));
assign O5pov6 = (Q6pov6 & X6pov6);
assign X6pov6 = (~(Pc1ov6 & Ojxnv6));
assign Q6pov6 = (~(Zec7z6[29] & Wc1ov6));
assign Rrj8v6 = (~(E7pov6 & L7pov6));
assign L7pov6 = (S7pov6 & Z7pov6);
assign Z7pov6 = (G8pov6 & N8pov6);
assign N8pov6 = (~(A81ov6 & Wk48v6));
assign G8pov6 = (U8pov6 & B9pov6);
assign B9pov6 = (~(Byc7z6[12] & V81ov6));
assign U8pov6 = (~(C91ov6 & Knynv6));
assign S7pov6 = (I9pov6 & P9pov6);
assign P9pov6 = (~(X91ov6 & Ips7v6));
assign I9pov6 = (~(Ea1ov6 & Pk48v6));
assign E7pov6 = (W9pov6 & Dapov6);
assign Dapov6 = (Kapov6 & Rapov6);
assign Rapov6 = (~(Nb1ov6 & Bps7v6));
assign Kapov6 = (~(Byc7z6[28] & Ub1ov6));
assign W9pov6 = (Yapov6 & Fbpov6);
assign Fbpov6 = (~(Pc1ov6 & Doxnv6));
assign Yapov6 = (~(Zec7z6[28] & Wc1ov6));
assign Krj8v6 = (~(Mbpov6 & Tbpov6));
assign Tbpov6 = (Acpov6 & Hcpov6);
assign Hcpov6 = (Ocpov6 & Vcpov6);
assign Vcpov6 = (~(A81ov6 & Ik48v6));
assign Ocpov6 = (Cdpov6 & Jdpov6);
assign Jdpov6 = (~(Byc7z6[11] & V81ov6));
assign Cdpov6 = (~(C91ov6 & Zrynv6));
assign Acpov6 = (Qdpov6 & Xdpov6);
assign Xdpov6 = (~(X91ov6 & Wps7v6));
assign Qdpov6 = (~(Ea1ov6 & Bk48v6));
assign Mbpov6 = (Eepov6 & Lepov6);
assign Lepov6 = (Sepov6 & Zepov6);
assign Zepov6 = (~(Nb1ov6 & Pps7v6));
assign Sepov6 = (~(Byc7z6[27] & Ub1ov6));
assign Eepov6 = (Gfpov6 & Nfpov6);
assign Nfpov6 = (~(Pc1ov6 & Ssxnv6));
assign Gfpov6 = (~(Zec7z6[27] & Wc1ov6));
assign Drj8v6 = (~(Ufpov6 & Bgpov6));
assign Bgpov6 = (Igpov6 & Pgpov6);
assign Pgpov6 = (Wgpov6 & Dhpov6);
assign Dhpov6 = (~(A81ov6 & Uj48v6));
assign Wgpov6 = (Khpov6 & Rhpov6);
assign Rhpov6 = (~(Byc7z6[10] & V81ov6));
assign Khpov6 = (~(C91ov6 & Owynv6));
assign Igpov6 = (Yhpov6 & Fipov6);
assign Fipov6 = (~(X91ov6 & Kqs7v6));
assign Yhpov6 = (~(Ea1ov6 & Nj48v6));
assign Ufpov6 = (Mipov6 & Tipov6);
assign Tipov6 = (Ajpov6 & Hjpov6);
assign Hjpov6 = (~(Nb1ov6 & Dqs7v6));
assign Ajpov6 = (~(Byc7z6[26] & Ub1ov6));
assign Mipov6 = (Ojpov6 & Vjpov6);
assign Vjpov6 = (~(Pc1ov6 & Hxxnv6));
assign Ojpov6 = (~(Zec7z6[26] & Wc1ov6));
assign Wqj8v6 = (~(Ckpov6 & Jkpov6));
assign Jkpov6 = (Qkpov6 & Xkpov6);
assign Xkpov6 = (Elpov6 & Llpov6);
assign Llpov6 = (~(A81ov6 & Gj48v6));
assign Elpov6 = (Slpov6 & Zlpov6);
assign Zlpov6 = (~(Byc7z6[9] & V81ov6));
assign Slpov6 = (~(C91ov6 & D1znv6));
assign Qkpov6 = (Gmpov6 & Nmpov6);
assign Nmpov6 = (~(X91ov6 & Yqs7v6));
assign Gmpov6 = (~(Ea1ov6 & Zi48v6));
assign Ckpov6 = (Umpov6 & Bnpov6);
assign Bnpov6 = (Inpov6 & Pnpov6);
assign Pnpov6 = (~(Nb1ov6 & Rqs7v6));
assign Inpov6 = (~(Byc7z6[25] & Ub1ov6));
assign Umpov6 = (Wnpov6 & Dopov6);
assign Dopov6 = (~(Pc1ov6 & W1ynv6));
assign Wnpov6 = (~(Zec7z6[25] & Wc1ov6));
assign Pqj8v6 = (~(Kopov6 & Ropov6));
assign Ropov6 = (Yopov6 & Fppov6);
assign Fppov6 = (Mppov6 & Tppov6);
assign Tppov6 = (~(A81ov6 & Si48v6));
assign Mppov6 = (Aqpov6 & Hqpov6);
assign Hqpov6 = (~(Byc7z6[8] & V81ov6));
assign Aqpov6 = (~(C91ov6 & S5znv6));
assign Yopov6 = (Oqpov6 & Vqpov6);
assign Vqpov6 = (~(X91ov6 & Mrs7v6));
assign Oqpov6 = (~(Ea1ov6 & Li48v6));
assign Kopov6 = (Crpov6 & Jrpov6);
assign Jrpov6 = (Qrpov6 & Xrpov6);
assign Xrpov6 = (~(Nb1ov6 & Frs7v6));
assign Qrpov6 = (~(Byc7z6[24] & Ub1ov6));
assign Crpov6 = (Espov6 & Lspov6);
assign Lspov6 = (~(Pc1ov6 & P9xnv6));
assign Espov6 = (~(Zec7z6[24] & Wc1ov6));
assign Iqj8v6 = (~(Sspov6 & Zspov6));
assign Zspov6 = (Gtpov6 & Ntpov6);
assign Ntpov6 = (Utpov6 & Bupov6);
assign Bupov6 = (~(A81ov6 & Ei48v6));
assign Utpov6 = (Iupov6 & Pupov6);
assign Pupov6 = (~(Byc7z6[7] & V81ov6));
assign Iupov6 = (~(C91ov6 & N1xnv6));
assign Gtpov6 = (Wupov6 & Dvpov6);
assign Dvpov6 = (~(X91ov6 & Ass7v6));
assign Wupov6 = (~(Ea1ov6 & Xh48v6));
assign Sspov6 = (Kvpov6 & Rvpov6);
assign Rvpov6 = (Yvpov6 & Fwpov6);
assign Fwpov6 = (~(Nb1ov6 & Trs7v6));
assign Yvpov6 = (~(Byc7z6[23] & Ub1ov6));
assign Kvpov6 = (Mwpov6 & Twpov6);
assign Twpov6 = (~(Pc1ov6 & Maynv6));
assign Mwpov6 = (~(Zec7z6[23] & Wc1ov6));
assign Bqj8v6 = (~(Axpov6 & Hxpov6));
assign Hxpov6 = (Oxpov6 & Vxpov6);
assign Vxpov6 = (Cypov6 & Jypov6);
assign Jypov6 = (~(A81ov6 & Qh48v6));
assign Cypov6 = (Qypov6 & Xypov6);
assign Xypov6 = (~(Byc7z6[6] & V81ov6));
assign Qypov6 = (~(C91ov6 & Eexnv6));
assign Oxpov6 = (Ezpov6 & Lzpov6);
assign Lzpov6 = (~(X91ov6 & Oss7v6));
assign Ezpov6 = (~(Ea1ov6 & Jh48v6));
assign Axpov6 = (Szpov6 & Zzpov6);
assign Zzpov6 = (G0qov6 & N0qov6);
assign N0qov6 = (~(Nb1ov6 & Hss7v6));
assign G0qov6 = (~(Byc7z6[22] & Ub1ov6));
assign Szpov6 = (U0qov6 & B1qov6);
assign B1qov6 = (~(Pc1ov6 & Bfynv6));
assign U0qov6 = (~(Zec7z6[22] & Wc1ov6));
assign Upj8v6 = (~(I1qov6 & P1qov6));
assign P1qov6 = (W1qov6 & D2qov6);
assign D2qov6 = (K2qov6 & R2qov6);
assign R2qov6 = (~(A81ov6 & Ch48v6));
assign K2qov6 = (Y2qov6 & F3qov6);
assign F3qov6 = (~(Byc7z6[5] & V81ov6));
assign Y2qov6 = (~(C91ov6 & Tixnv6));
assign W1qov6 = (M3qov6 & T3qov6);
assign T3qov6 = (~(X91ov6 & Cts7v6));
assign M3qov6 = (~(Ea1ov6 & Vg48v6));
assign I1qov6 = (A4qov6 & H4qov6);
assign H4qov6 = (O4qov6 & V4qov6);
assign V4qov6 = (~(Nb1ov6 & Vss7v6));
assign O4qov6 = (~(Byc7z6[21] & Ub1ov6));
assign A4qov6 = (C5qov6 & J5qov6);
assign J5qov6 = (~(Pc1ov6 & Qjynv6));
assign C5qov6 = (~(Zec7z6[21] & Wc1ov6));
assign Npj8v6 = (~(Q5qov6 & X5qov6));
assign X5qov6 = (E6qov6 & L6qov6);
assign L6qov6 = (S6qov6 & Z6qov6);
assign Z6qov6 = (~(A81ov6 & Og48v6));
assign S6qov6 = (G7qov6 & N7qov6);
assign N7qov6 = (~(Byc7z6[4] & V81ov6));
assign G7qov6 = (~(C91ov6 & Inxnv6));
assign E6qov6 = (U7qov6 & B8qov6);
assign B8qov6 = (~(X91ov6 & Qts7v6));
assign U7qov6 = (~(Ea1ov6 & Hg48v6));
assign Q5qov6 = (I8qov6 & P8qov6);
assign P8qov6 = (W8qov6 & D9qov6);
assign D9qov6 = (~(Nb1ov6 & Jts7v6));
assign W8qov6 = (~(Byc7z6[20] & Ub1ov6));
assign I8qov6 = (K9qov6 & R9qov6);
assign R9qov6 = (~(Pc1ov6 & Foynv6));
assign K9qov6 = (~(Zec7z6[20] & Wc1ov6));
assign Gpj8v6 = (~(Y9qov6 & Faqov6));
assign Faqov6 = (Maqov6 & Taqov6);
assign Taqov6 = (Abqov6 & Hbqov6);
assign Hbqov6 = (~(A81ov6 & Ag48v6));
assign Abqov6 = (Obqov6 & Vbqov6);
assign Vbqov6 = (~(Byc7z6[3] & V81ov6));
assign Obqov6 = (~(C91ov6 & Xrxnv6));
assign Maqov6 = (Ccqov6 & Jcqov6);
assign Jcqov6 = (~(X91ov6 & Eus7v6));
assign Ccqov6 = (~(Ea1ov6 & Tf48v6));
assign Y9qov6 = (Qcqov6 & Xcqov6);
assign Xcqov6 = (Edqov6 & Ldqov6);
assign Ldqov6 = (~(Nb1ov6 & Xts7v6));
assign Edqov6 = (~(Byc7z6[19] & Ub1ov6));
assign Qcqov6 = (Sdqov6 & Zdqov6);
assign Zdqov6 = (~(Pc1ov6 & Usynv6));
assign Sdqov6 = (~(Zec7z6[19] & Wc1ov6));
assign Zoj8v6 = (~(Geqov6 & Neqov6));
assign Neqov6 = (Ueqov6 & Bfqov6);
assign Bfqov6 = (Ifqov6 & Pfqov6);
assign Pfqov6 = (~(A81ov6 & Mf48v6));
assign Ifqov6 = (Wfqov6 & Dgqov6);
assign Dgqov6 = (~(Byc7z6[2] & V81ov6));
assign Wfqov6 = (~(C91ov6 & Mwxnv6));
assign Ueqov6 = (Kgqov6 & Rgqov6);
assign Rgqov6 = (~(X91ov6 & Sus7v6));
assign Kgqov6 = (~(Ea1ov6 & Ff48v6));
assign Geqov6 = (Ygqov6 & Fhqov6);
assign Fhqov6 = (Mhqov6 & Thqov6);
assign Thqov6 = (~(Nb1ov6 & Lus7v6));
assign Mhqov6 = (~(Byc7z6[18] & Ub1ov6));
assign Ygqov6 = (Aiqov6 & Hiqov6);
assign Hiqov6 = (~(Pc1ov6 & Jxynv6));
assign Aiqov6 = (~(Zec7z6[18] & Wc1ov6));
assign Soj8v6 = (~(Oiqov6 & Viqov6));
assign Viqov6 = (Cjqov6 & Jjqov6);
assign Jjqov6 = (Qjqov6 & Xjqov6);
assign Xjqov6 = (~(A81ov6 & Ye48v6));
assign Qjqov6 = (Ekqov6 & Lkqov6);
assign Lkqov6 = (~(Byc7z6[1] & V81ov6));
assign Ekqov6 = (~(C91ov6 & B1ynv6));
assign Cjqov6 = (Skqov6 & Zkqov6);
assign Zkqov6 = (~(X91ov6 & Gvs7v6));
assign Skqov6 = (~(Ea1ov6 & Re48v6));
assign Oiqov6 = (Glqov6 & Nlqov6);
assign Nlqov6 = (Ulqov6 & Bmqov6);
assign Bmqov6 = (~(Nb1ov6 & Zus7v6));
assign Ulqov6 = (~(Byc7z6[17] & Ub1ov6));
assign Glqov6 = (Imqov6 & Pmqov6);
assign Pmqov6 = (~(Pc1ov6 & Y1znv6));
assign Imqov6 = (~(Zec7z6[17] & Wc1ov6));
assign Loj8v6 = (~(Wmqov6 & Dnqov6));
assign Dnqov6 = (Knqov6 & Rnqov6);
assign Rnqov6 = (Ynqov6 & Foqov6);
assign Foqov6 = (~(A81ov6 & Ke48v6));
assign Ynqov6 = (Moqov6 & Toqov6);
assign Toqov6 = (~(Byc7z6[0] & V81ov6));
assign V81ov6 = (~(Apqov6 | Hpqov6));
assign Moqov6 = (~(C91ov6 & Kaxnv6));
assign C91ov6 = (~(Opqov6 | Apqov6));
assign Apqov6 = (!Bvoov6);
assign Knqov6 = (Vpqov6 & Cqqov6);
assign Cqqov6 = (~(X91ov6 & Nvs7v6));
assign Vpqov6 = (~(Ea1ov6 & De48v6));
assign Wmqov6 = (Jqqov6 & Qqqov6);
assign Qqqov6 = (Xqqov6 & Erqov6);
assign Erqov6 = (~(Nb1ov6 & D9o7v6));
assign Xqqov6 = (~(Byc7z6[16] & Ub1ov6));
assign Jqqov6 = (Lrqov6 & Srqov6);
assign Srqov6 = (~(Pc1ov6 & N6znv6));
assign Lrqov6 = (~(Zec7z6[16] & Wc1ov6));
assign Eoj8v6 = (~(Zrqov6 & Gsqov6));
assign Gsqov6 = (Nsqov6 & Usqov6);
assign Usqov6 = (Btqov6 & Itqov6);
assign Itqov6 = (~(Bvoov6 & P8o7v6));
assign Btqov6 = (Ptqov6 & Wtqov6);
assign Wtqov6 = (~(Wvoov6 & Byc7z6[31]));
assign Ptqov6 = (~(Dwoov6 & P2xnv6));
assign Nsqov6 = (Duqov6 & Kuqov6);
assign Kuqov6 = (~(X91ov6 & Y9o7v6));
assign Duqov6 = (~(Ea1ov6 & Fao7v6));
assign Zrqov6 = (Ruqov6 & Yuqov6);
assign Yuqov6 = (Fvqov6 & Mvqov6);
assign Mvqov6 = (~(Nb1ov6 & W8o7v6));
assign Fvqov6 = (~(Ub1ov6 & Byc7z6[15]));
assign Ruqov6 = (Tvqov6 & Awqov6);
assign Awqov6 = (~(Pc1ov6 & R9ynv6));
assign Tvqov6 = (~(Zec7z6[15] & Wc1ov6));
assign Xnj8v6 = (~(Hwqov6 & Owqov6));
assign Owqov6 = (Vwqov6 & Cxqov6);
assign Cxqov6 = (Jxqov6 & Qxqov6);
assign Qxqov6 = (~(Bvoov6 & K9o7v6));
assign Jxqov6 = (Xxqov6 & Eyqov6);
assign Eyqov6 = (~(Byc7z6[30] & Wvoov6));
assign Xxqov6 = (~(Dwoov6 & Zexnv6));
assign Vwqov6 = (Lyqov6 & Syqov6);
assign Syqov6 = (~(X91ov6 & Rl48v6));
assign Lyqov6 = (~(Ea1ov6 & Gos7v6));
assign Hwqov6 = (Zyqov6 & Gzqov6);
assign Gzqov6 = (Nzqov6 & Uzqov6);
assign Uzqov6 = (~(Nb1ov6 & R9o7v6));
assign Nzqov6 = (~(Byc7z6[14] & Ub1ov6));
assign Zyqov6 = (B0rov6 & I0rov6);
assign I0rov6 = (~(Pc1ov6 & Geynv6));
assign B0rov6 = (~(Zec7z6[14] & Wc1ov6));
assign Qnj8v6 = (~(P0rov6 & W0rov6));
assign W0rov6 = (D1rov6 & K1rov6);
assign K1rov6 = (R1rov6 & Y1rov6);
assign Y1rov6 = (~(Bvoov6 & Nos7v6));
assign R1rov6 = (F2rov6 & M2rov6);
assign M2rov6 = (~(Byc7z6[29] & Wvoov6));
assign F2rov6 = (~(Dwoov6 & Ojxnv6));
assign D1rov6 = (T2rov6 & A3rov6);
assign A3rov6 = (~(X91ov6 & Kl48v6));
assign T2rov6 = (~(Ea1ov6 & Uos7v6));
assign P0rov6 = (H3rov6 & O3rov6);
assign O3rov6 = (V3rov6 & C4rov6);
assign C4rov6 = (~(Nb1ov6 & Dl48v6));
assign V3rov6 = (~(Byc7z6[13] & Ub1ov6));
assign H3rov6 = (J4rov6 & Q4rov6);
assign Q4rov6 = (~(Pc1ov6 & Viynv6));
assign J4rov6 = (~(Zec7z6[13] & Wc1ov6));
assign Jnj8v6 = (~(X4rov6 & E5rov6));
assign E5rov6 = (L5rov6 & S5rov6);
assign S5rov6 = (Z5rov6 & G6rov6);
assign G6rov6 = (~(Bvoov6 & Bps7v6));
assign Z5rov6 = (N6rov6 & U6rov6);
assign U6rov6 = (~(Byc7z6[28] & Wvoov6));
assign N6rov6 = (~(Dwoov6 & Doxnv6));
assign L5rov6 = (B7rov6 & I7rov6);
assign I7rov6 = (~(X91ov6 & Wk48v6));
assign B7rov6 = (~(Ea1ov6 & Ips7v6));
assign X4rov6 = (P7rov6 & W7rov6);
assign W7rov6 = (D8rov6 & K8rov6);
assign K8rov6 = (~(Nb1ov6 & Pk48v6));
assign D8rov6 = (~(Byc7z6[12] & Ub1ov6));
assign P7rov6 = (R8rov6 & Y8rov6);
assign Y8rov6 = (~(Pc1ov6 & Knynv6));
assign R8rov6 = (~(Zec7z6[12] & Wc1ov6));
assign Cnj8v6 = (~(F9rov6 & M9rov6));
assign M9rov6 = (T9rov6 & Aarov6);
assign Aarov6 = (Harov6 & Oarov6);
assign Oarov6 = (~(Bvoov6 & Pps7v6));
assign Harov6 = (Varov6 & Cbrov6);
assign Cbrov6 = (~(Byc7z6[27] & Wvoov6));
assign Varov6 = (~(Dwoov6 & Ssxnv6));
assign T9rov6 = (Jbrov6 & Qbrov6);
assign Qbrov6 = (~(X91ov6 & Ik48v6));
assign Jbrov6 = (~(Ea1ov6 & Wps7v6));
assign F9rov6 = (Xbrov6 & Ecrov6);
assign Ecrov6 = (Lcrov6 & Scrov6);
assign Scrov6 = (~(Nb1ov6 & Bk48v6));
assign Lcrov6 = (~(Byc7z6[11] & Ub1ov6));
assign Xbrov6 = (Zcrov6 & Gdrov6);
assign Gdrov6 = (~(Pc1ov6 & Zrynv6));
assign Zcrov6 = (~(Zec7z6[11] & Wc1ov6));
assign Vmj8v6 = (Vs9ov6 ? Qwddt6 : A4a7z6);
assign Omj8v6 = (!Ndrov6);
assign Ndrov6 = (N3onv6 ? Udrov6 : K397z6);
assign Udrov6 = (~(Qwddt6 & Berov6));
assign Berov6 = (~(Zhbdt6 & Ierov6));
assign Hmj8v6 = (~(Perov6 & Werov6));
assign Werov6 = (~(Snvnv6 & Ovbdt6));
assign Perov6 = (~(M5e7z6[1] & Dcnov6));
assign Amj8v6 = (~(Dfrov6 & Kfrov6));
assign Kfrov6 = (Rfrov6 & Yfrov6);
assign Yfrov6 = (Fgrov6 & Mgrov6);
assign Mgrov6 = (~(Bvoov6 & Dqs7v6));
assign Fgrov6 = (Tgrov6 & Ahrov6);
assign Ahrov6 = (~(Byc7z6[26] & Wvoov6));
assign Tgrov6 = (~(Dwoov6 & Hxxnv6));
assign Rfrov6 = (Hhrov6 & Ohrov6);
assign Ohrov6 = (~(X91ov6 & Uj48v6));
assign Hhrov6 = (~(Ea1ov6 & Kqs7v6));
assign Dfrov6 = (Vhrov6 & Cirov6);
assign Cirov6 = (Jirov6 & Qirov6);
assign Qirov6 = (~(Nb1ov6 & Nj48v6));
assign Jirov6 = (~(Byc7z6[10] & Ub1ov6));
assign Vhrov6 = (Xirov6 & Ejrov6);
assign Ejrov6 = (~(Pc1ov6 & Owynv6));
assign Xirov6 = (~(Zec7z6[10] & Wc1ov6));
assign Tlj8v6 = (~(Ljrov6 & Sjrov6));
assign Sjrov6 = (Zjrov6 & Gkrov6);
assign Gkrov6 = (Nkrov6 & Ukrov6);
assign Ukrov6 = (~(Bvoov6 & Rqs7v6));
assign Nkrov6 = (Blrov6 & Ilrov6);
assign Ilrov6 = (~(Byc7z6[25] & Wvoov6));
assign Blrov6 = (~(Dwoov6 & W1ynv6));
assign Zjrov6 = (Plrov6 & Wlrov6);
assign Wlrov6 = (~(X91ov6 & Gj48v6));
assign Plrov6 = (~(Ea1ov6 & Yqs7v6));
assign Ljrov6 = (Dmrov6 & Kmrov6);
assign Kmrov6 = (Rmrov6 & Ymrov6);
assign Ymrov6 = (~(Nb1ov6 & Zi48v6));
assign Rmrov6 = (~(Byc7z6[9] & Ub1ov6));
assign Dmrov6 = (Fnrov6 & Mnrov6);
assign Mnrov6 = (~(Pc1ov6 & D1znv6));
assign Fnrov6 = (~(Zec7z6[9] & Wc1ov6));
assign Mlj8v6 = (~(Tnrov6 & Aorov6));
assign Aorov6 = (Horov6 & Oorov6);
assign Oorov6 = (Vorov6 & Cprov6);
assign Cprov6 = (~(Bvoov6 & Frs7v6));
assign Vorov6 = (Jprov6 & Qprov6);
assign Qprov6 = (~(Byc7z6[24] & Wvoov6));
assign Jprov6 = (~(Dwoov6 & P9xnv6));
assign Horov6 = (Xprov6 & Eqrov6);
assign Eqrov6 = (~(X91ov6 & Si48v6));
assign Xprov6 = (~(Ea1ov6 & Mrs7v6));
assign Tnrov6 = (Lqrov6 & Sqrov6);
assign Sqrov6 = (Zqrov6 & Grrov6);
assign Grrov6 = (~(Nb1ov6 & Li48v6));
assign Zqrov6 = (~(Byc7z6[8] & Ub1ov6));
assign Lqrov6 = (Nrrov6 & Urrov6);
assign Urrov6 = (~(Pc1ov6 & S5znv6));
assign Nrrov6 = (~(Zec7z6[8] & Wc1ov6));
assign Flj8v6 = (~(Bsrov6 & Isrov6));
assign Isrov6 = (~(Uobdt6 & Dcnov6));
assign Ykj8v6 = (~(Psrov6 & Wsrov6));
assign Wsrov6 = (Dtrov6 & Ktrov6);
assign Ktrov6 = (Rtrov6 & Ytrov6);
assign Ytrov6 = (~(Bvoov6 & Trs7v6));
assign Rtrov6 = (Furov6 & Murov6);
assign Murov6 = (~(Byc7z6[23] & Wvoov6));
assign Furov6 = (~(Dwoov6 & Maynv6));
assign Dtrov6 = (Turov6 & Avrov6);
assign Avrov6 = (~(X91ov6 & Ei48v6));
assign Turov6 = (~(Ea1ov6 & Ass7v6));
assign Psrov6 = (Hvrov6 & Ovrov6);
assign Ovrov6 = (Vvrov6 & Cwrov6);
assign Cwrov6 = (~(Nb1ov6 & Xh48v6));
assign Vvrov6 = (~(Byc7z6[7] & Ub1ov6));
assign Hvrov6 = (Jwrov6 & Qwrov6);
assign Qwrov6 = (~(Pc1ov6 & N1xnv6));
assign Jwrov6 = (~(Zec7z6[7] & Wc1ov6));
assign Rkj8v6 = (~(Xwrov6 & Exrov6));
assign Exrov6 = (Lxrov6 & Sxrov6);
assign Lxrov6 = (~(Zxrov6 & Zec7z6[7]));
assign Xwrov6 = (Gyrov6 & Nyrov6);
assign Nyrov6 = (~(Uyrov6 & Zec7z6[9]));
assign Gyrov6 = (~(Ide7z6[1] & Vs9ov6));
assign Kkj8v6 = (~(Bzrov6 & Izrov6));
assign Izrov6 = (Pzrov6 & Sxrov6);
assign Pzrov6 = (~(Zxrov6 & Zec7z6[8]));
assign Bzrov6 = (Wzrov6 & D0sov6);
assign D0sov6 = (~(Uyrov6 & Zec7z6[10]));
assign Wzrov6 = (~(Ide7z6[2] & Vs9ov6));
assign Dkj8v6 = (~(K0sov6 & R0sov6));
assign R0sov6 = (Y0sov6 & Sxrov6);
assign Sxrov6 = (~(F1sov6 & M1sov6));
assign M1sov6 = (T1sov6 & A2sov6);
assign F1sov6 = (N3onv6 & H2sov6);
assign Y0sov6 = (~(Zxrov6 & Zec7z6[9]));
assign K0sov6 = (O2sov6 & V2sov6);
assign V2sov6 = (~(Uyrov6 & Zec7z6[11]));
assign O2sov6 = (~(Ide7z6[3] & Vs9ov6));
assign Wjj8v6 = (~(C3sov6 & J3sov6));
assign J3sov6 = (~(K7e7z6[0] & Dcnov6));
assign C3sov6 = (Q3sov6 & X3sov6);
assign Q3sov6 = (~(E4sov6 & L4sov6));
assign E4sov6 = (N3onv6 & Zec7z6[30]);
assign Pjj8v6 = (~(X3sov6 & S4sov6));
assign S4sov6 = (~(K7e7z6[1] & Dcnov6));
assign X3sov6 = (~(Z4sov6 & G5sov6));
assign Z4sov6 = (N3onv6 & Zec7z6[7]);
assign Ijj8v6 = (~(N5sov6 & U5sov6));
assign U5sov6 = (B6sov6 & I6sov6);
assign I6sov6 = (P6sov6 & W6sov6);
assign W6sov6 = (~(Bvoov6 & Hss7v6));
assign P6sov6 = (D7sov6 & K7sov6);
assign K7sov6 = (~(Byc7z6[22] & Wvoov6));
assign D7sov6 = (~(Dwoov6 & Bfynv6));
assign B6sov6 = (R7sov6 & Y7sov6);
assign Y7sov6 = (~(X91ov6 & Qh48v6));
assign R7sov6 = (~(Ea1ov6 & Oss7v6));
assign N5sov6 = (F8sov6 & M8sov6);
assign M8sov6 = (T8sov6 & A9sov6);
assign A9sov6 = (~(Nb1ov6 & Jh48v6));
assign T8sov6 = (~(Byc7z6[6] & Ub1ov6));
assign F8sov6 = (H9sov6 & O9sov6);
assign O9sov6 = (~(Pc1ov6 & Eexnv6));
assign H9sov6 = (~(Zec7z6[6] & Wc1ov6));
assign Bjj8v6 = (~(V9sov6 & Casov6));
assign Casov6 = (Jasov6 & Qasov6);
assign Qasov6 = (~(Zxrov6 & Zec7z6[6]));
assign Zxrov6 = (~(H2sov6 | Vs9ov6));
assign Jasov6 = (~(Uyrov6 & Zec7z6[8]));
assign Uyrov6 = (~(Vs9ov6 | T1sov6));
assign V9sov6 = (Xasov6 & Ebsov6);
assign Ebsov6 = (~(Ide7z6[0] & Vs9ov6));
assign Xasov6 = (~(Yxd7z6[0] & Zec7z6[11]));
assign Uij8v6 = (~(Lbsov6 & Sbsov6));
assign Sbsov6 = (~(I5cdt6 & Dcnov6));
assign Lbsov6 = (~(Zbsov6 & N3onv6));
assign Nij8v6 = (~(Gcsov6 & Ncsov6));
assign Ncsov6 = (Ucsov6 & Bdsov6);
assign Bdsov6 = (Idsov6 & Pdsov6);
assign Pdsov6 = (~(Bvoov6 & Vss7v6));
assign Idsov6 = (Wdsov6 & Desov6);
assign Desov6 = (~(Byc7z6[21] & Wvoov6));
assign Wdsov6 = (~(Dwoov6 & Qjynv6));
assign Ucsov6 = (Kesov6 & Resov6);
assign Resov6 = (~(X91ov6 & Ch48v6));
assign Kesov6 = (~(Ea1ov6 & Cts7v6));
assign Gcsov6 = (Yesov6 & Ffsov6);
assign Ffsov6 = (Mfsov6 & Tfsov6);
assign Tfsov6 = (~(Nb1ov6 & Vg48v6));
assign Mfsov6 = (~(Byc7z6[5] & Ub1ov6));
assign Yesov6 = (Agsov6 & Hgsov6);
assign Hgsov6 = (~(Pc1ov6 & Tixnv6));
assign Agsov6 = (~(Zec7z6[5] & Wc1ov6));
assign Gij8v6 = (~(Ogsov6 & Vgsov6));
assign Vgsov6 = (~(Chsov6 & Jhsov6));
assign Chsov6 = (Snvnv6 & Zec7z6[0]);
assign Ogsov6 = (~(I9e7z6[1] & Dcnov6));
assign Zhj8v6 = (~(Qhsov6 & Xhsov6));
assign Xhsov6 = (Eisov6 & Lisov6);
assign Lisov6 = (Sisov6 & Zisov6);
assign Zisov6 = (~(Bvoov6 & Jts7v6));
assign Sisov6 = (Gjsov6 & Njsov6);
assign Njsov6 = (~(Byc7z6[20] & Wvoov6));
assign Gjsov6 = (~(Dwoov6 & Foynv6));
assign Eisov6 = (Ujsov6 & Bksov6);
assign Bksov6 = (~(X91ov6 & Og48v6));
assign Ujsov6 = (~(Ea1ov6 & Qts7v6));
assign Qhsov6 = (Iksov6 & Pksov6);
assign Pksov6 = (Wksov6 & Dlsov6);
assign Dlsov6 = (~(Nb1ov6 & Hg48v6));
assign Wksov6 = (~(Byc7z6[4] & Ub1ov6));
assign Iksov6 = (Klsov6 & Rlsov6);
assign Rlsov6 = (~(Pc1ov6 & Inxnv6));
assign Klsov6 = (~(Zec7z6[4] & Wc1ov6));
assign Shj8v6 = (~(Ylsov6 & Fmsov6));
assign Fmsov6 = (~(Mmsov6 & Tmsov6));
assign Mmsov6 = (Ansov6 & Snvnv6);
assign Ylsov6 = (~(M5e7z6[0] & Dcnov6));
assign Lhj8v6 = (~(Hnsov6 & Onsov6));
assign Onsov6 = (~(Snvnv6 & Vnsov6));
assign Vnsov6 = (~(Cosov6 & Josov6));
assign Josov6 = (Qosov6 & Xosov6);
assign Qosov6 = (Epsov6 & Lpsov6);
assign Cosov6 = (Spsov6 & Zpsov6);
assign Spsov6 = (Gqsov6 & Nqsov6);
assign Nqsov6 = (Qtnov6 | O7onv6);
assign O7onv6 = (Uqsov6 & Brsov6);
assign Brsov6 = (Irsov6 & Prsov6);
assign Uqsov6 = (Wrsov6 & Dssov6);
assign Gqsov6 = (~(Tmsov6 & Kssov6));
assign Hnsov6 = (~(Lwfdt6 & Vs9ov6));
assign Ehj8v6 = (~(Rssov6 & Yssov6));
assign Yssov6 = (~(Ftsov6 & Mtsov6));
assign Ftsov6 = (Snvnv6 & Uqd7z6[20]);
assign Rssov6 = (~(M3e7z6[1] & Dcnov6));
assign Xgj8v6 = (~(Ttsov6 & Ausov6));
assign Ausov6 = (~(Husov6 & Mtsov6));
assign Husov6 = (Snvnv6 & E9onv6);
assign Ttsov6 = (~(M3e7z6[0] & Dcnov6));
assign Qgj8v6 = (~(Ousov6 & Vusov6));
assign Vusov6 = (~(Cvsov6 & Jhsov6));
assign Cvsov6 = (Snvnv6 & Zec7z6[4]);
assign Ousov6 = (~(I9e7z6[0] & Dcnov6));
assign Jgj8v6 = (~(Jvsov6 & Qvsov6));
assign Qvsov6 = (Xvsov6 & Ewsov6);
assign Ewsov6 = (Lwsov6 & Swsov6);
assign Swsov6 = (~(Bvoov6 & Xts7v6));
assign Lwsov6 = (Zwsov6 & Gxsov6);
assign Gxsov6 = (~(Byc7z6[19] & Wvoov6));
assign Zwsov6 = (~(Dwoov6 & Usynv6));
assign Xvsov6 = (Nxsov6 & Uxsov6);
assign Uxsov6 = (~(X91ov6 & Ag48v6));
assign Nxsov6 = (~(Ea1ov6 & Eus7v6));
assign Jvsov6 = (Bysov6 & Iysov6);
assign Iysov6 = (Pysov6 & Wysov6);
assign Wysov6 = (~(Nb1ov6 & Tf48v6));
assign Pysov6 = (~(Byc7z6[3] & Ub1ov6));
assign Bysov6 = (Dzsov6 & Kzsov6);
assign Kzsov6 = (~(Pc1ov6 & Xrxnv6));
assign Dzsov6 = (~(Zec7z6[3] & Wc1ov6));
assign Cgj8v6 = (~(Rzsov6 & Yzsov6));
assign Yzsov6 = (F0tov6 & M0tov6);
assign M0tov6 = (T0tov6 & A1tov6);
assign A1tov6 = (~(Bvoov6 & Lus7v6));
assign T0tov6 = (H1tov6 & O1tov6);
assign O1tov6 = (~(Byc7z6[18] & Wvoov6));
assign H1tov6 = (~(Dwoov6 & Jxynv6));
assign F0tov6 = (V1tov6 & C2tov6);
assign C2tov6 = (~(X91ov6 & Mf48v6));
assign V1tov6 = (~(Ea1ov6 & Sus7v6));
assign Rzsov6 = (J2tov6 & Q2tov6);
assign Q2tov6 = (X2tov6 & E3tov6);
assign E3tov6 = (~(Nb1ov6 & Ff48v6));
assign X2tov6 = (~(Byc7z6[2] & Ub1ov6));
assign J2tov6 = (L3tov6 & S3tov6);
assign S3tov6 = (~(Pc1ov6 & Mwxnv6));
assign L3tov6 = (~(Zec7z6[2] & Wc1ov6));
assign Vfj8v6 = (~(Z3tov6 & G4tov6));
assign G4tov6 = (N4tov6 & U4tov6);
assign U4tov6 = (B5tov6 & I5tov6);
assign I5tov6 = (~(Bvoov6 & Zus7v6));
assign Bvoov6 = (~(P5tov6 | W5tov6));
assign P5tov6 = (K6tov6 ? C3mnv6 : D6tov6);
assign B5tov6 = (R6tov6 & Y6tov6);
assign Y6tov6 = (~(Byc7z6[17] & Wvoov6));
assign Wvoov6 = (~(F7tov6 | Hpqov6));
assign R6tov6 = (~(Dwoov6 & Y1znv6));
assign Dwoov6 = (~(F7tov6 | Opqov6));
assign F7tov6 = (!A81ov6);
assign A81ov6 = (~(M7tov6 | W5tov6));
assign M7tov6 = (K6tov6 ? K0mnv6 : T7tov6);
assign N4tov6 = (A8tov6 & H8tov6);
assign H8tov6 = (~(X91ov6 & Ye48v6));
assign X91ov6 = (O8tov6 & V8tov6);
assign O8tov6 = (K6tov6 ? W6mnv6 : Bfd7z6[0]);
assign A8tov6 = (~(Ea1ov6 & Gvs7v6));
assign Ea1ov6 = (~(C9tov6 | W5tov6));
assign C9tov6 = (K6tov6 ? S4mnv6 : J9tov6);
assign Z3tov6 = (Q9tov6 & X9tov6);
assign X9tov6 = (Eatov6 & Latov6);
assign Latov6 = (~(Nb1ov6 & Re48v6));
assign Nb1ov6 = (~(Satov6 | W5tov6));
assign W5tov6 = (!V8tov6);
assign V8tov6 = (Zatov6 & Gbtov6);
assign Satov6 = (K6tov6 ? X3mnv6 : Nbtov6);
assign Eatov6 = (~(Byc7z6[1] & Ub1ov6));
assign Ub1ov6 = (Ubtov6 & Zatov6);
assign Ubtov6 = (Bctov6 & Opqov6);
assign Q9tov6 = (Ictov6 & Pctov6);
assign Pctov6 = (~(Pc1ov6 & B1ynv6));
assign Pc1ov6 = (Wctov6 & Hpqov6);
assign Wctov6 = (Zatov6 & Bctov6);
assign Bctov6 = (!Gbtov6);
assign Gbtov6 = (~(Ddtov6 | Mao7v6));
assign Ddtov6 = (K6tov6 ? M1mnv6 : Bfd7z6[4]);
assign Zatov6 = (!Wc1ov6);
assign Ictov6 = (~(Zec7z6[1] & Wc1ov6));
assign Wc1ov6 = (~(Kdtov6 & Rdtov6));
assign Kdtov6 = (~(Ydtov6 & M8mnv6));
assign Ydtov6 = (Ij1ov6 & Fetov6);
assign Ofj8v6 = (~(Metov6 & Tetov6));
assign Tetov6 = (~(Aftov6 & Hftov6));
assign Metov6 = (~(Ibe7z6[0] & Dcnov6));
assign Hfj8v6 = (~(Oftov6 & Vftov6));
assign Vftov6 = (~(Cgtov6 & Aftov6));
assign Cgtov6 = (Ovbdt6 & Jgtov6);
assign Oftov6 = (~(Ibe7z6[1] & Dcnov6));
assign Afj8v6 = (~(Qgtov6 & Xgtov6));
assign Xgtov6 = (~(Ehtov6 & Aftov6));
assign Qgtov6 = (~(Ibe7z6[2] & Dcnov6));
assign Tej8v6 = (~(Lhtov6 & Shtov6));
assign Shtov6 = (~(Zhtov6 & Aftov6));
assign Aftov6 = (Gitov6 & Nitov6);
assign Lhtov6 = (~(Ibe7z6[3] & Dcnov6));
assign Mej8v6 = (~(Uitov6 & Bjtov6));
assign Bjtov6 = (~(Nitov6 & Ijtov6));
assign Nitov6 = (Pjtov6 & Wjtov6);
assign Wjtov6 = (Dktov6 & Uqd7z6[20]);
assign Dktov6 = (Kktov6 & Rktov6);
assign Pjtov6 = (Tmsov6 & Snvnv6);
assign Uitov6 = (~(Ibe7z6[4] & Dcnov6));
assign Fej8v6 = (~(Yktov6 & Fltov6));
assign Fltov6 = (~(N3onv6 & Mltov6));
assign Mltov6 = (~(Tltov6 & Amtov6));
assign Yktov6 = (Hmtov6 | Sb77z6);
assign Ydj8v6 = (~(Omtov6 & Vmtov6));
assign Vmtov6 = (Vs9ov6 | Cntov6);
assign Omtov6 = (~(I0c7z6[1] & Dcnov6));
assign Rdj8v6 = (~(Jntov6 & Mmehw6));
assign Mmehw6 = (Vs9ov6 | Tmehw6);
assign Jntov6 = (~(I0c7z6[0] & Dcnov6));
assign Kdj8v6 = (Shmov6 ? Edh7z6[0] : Wbhnv6);
assign Ddj8v6 = (Uimov6 ? Gsb7z6[0] : Wbhnv6);
assign Wcj8v6 = (Shmov6 ? Edh7z6[1] : Anehw6);
assign Pcj8v6 = (Uimov6 ? Gsb7z6[1] : Anehw6);
assign Icj8v6 = (~(Hnehw6 & Onehw6));
assign Onehw6 = (~(N3onv6 & Vnehw6));
assign Vnehw6 = (~(Coehw6 & Joehw6));
assign Joehw6 = (Qoehw6 & Xoehw6);
assign Xoehw6 = (Epehw6 & Lpehw6);
assign Lpehw6 = (~(Spehw6 & Zpehw6));
assign Spehw6 = (~(Gqehw6 & Nqehw6));
assign Epehw6 = (Uqehw6 | Zec7z6[7]);
assign Qoehw6 = (Brehw6 & Irehw6);
assign Irehw6 = (~(Prehw6 & Qtnov6));
assign Brehw6 = (Wrehw6 | Dsehw6);
assign Coehw6 = (Ksehw6 & Rsehw6);
assign Rsehw6 = (Ysehw6 & Ftehw6);
assign Ftehw6 = (~(Mtehw6 & Ttehw6));
assign Ysehw6 = (~(Auehw6 & Zec7z6[8]));
assign Ksehw6 = (Huehw6 & Ouehw6);
assign Ouehw6 = (~(Vuehw6 & Cvehw6));
assign Hnehw6 = (~(Mrbdt6 & Dcnov6));
assign Bcj8v6 = (Shmov6 ? Vt2et6 : Mrbdt6);
assign Ubj8v6 = (~(Jvehw6 & Qvehw6));
assign Qvehw6 = (~(T3cdt6 & Dcnov6));
assign Jvehw6 = (Vs9ov6 | Xvehw6);
assign Nbj8v6 = (~(Ewehw6 & Lwehw6));
assign Lwehw6 = (~(Swehw6 & Snvnv6));
assign Swehw6 = (~(Tmehw6 | Zwehw6));
assign Tmehw6 = (Gxehw6 & Nxehw6);
assign Nxehw6 = (Uxehw6 & Byehw6);
assign Byehw6 = (Iyehw6 & Wrehw6);
assign Iyehw6 = (Pyehw6 & Wyehw6);
assign Uxehw6 = (Dzehw6 & Kzehw6);
assign Kzehw6 = (~(Uqd7z6[20] & Rzehw6));
assign Rzehw6 = (~(Yzehw6 & F0fhw6));
assign Dzehw6 = (~(M0fhw6 & Zec7z6[26]));
assign Gxehw6 = (T0fhw6 & A1fhw6);
assign A1fhw6 = (H1fhw6 & O1fhw6);
assign O1fhw6 = (~(Vuehw6 & V1fhw6));
assign H1fhw6 = (C2fhw6 & J2fhw6);
assign J2fhw6 = (~(Mtehw6 & Fcinv6));
assign C2fhw6 = (T6onv6 | Q2fhw6);
assign T0fhw6 = (Huehw6 & X2fhw6);
assign X2fhw6 = (~(E3fhw6 & Auehw6));
assign Huehw6 = (L3fhw6 & S3fhw6);
assign S3fhw6 = (~(Vuehw6 & Z3fhw6));
assign L3fhw6 = (G4fhw6 & N4fhw6);
assign G4fhw6 = (~(U4fhw6 & B5fhw6));
assign B5fhw6 = (I5fhw6 & Gginv6);
assign U4fhw6 = (P5fhw6 & V1fhw6);
assign Ewehw6 = (~(W5fhw6 & Tfh7z6[0]));
assign Gbj8v6 = (~(D6fhw6 & K6fhw6));
assign K6fhw6 = (~(R6fhw6 & Snvnv6));
assign R6fhw6 = (~(Cntov6 | Zwehw6));
assign Cntov6 = (Y6fhw6 & F7fhw6);
assign F7fhw6 = (M7fhw6 & T7fhw6);
assign T7fhw6 = (A8fhw6 & H8fhw6);
assign H8fhw6 = (O8fhw6 & Amtov6);
assign A8fhw6 = (~(Zbsov6 | V8fhw6));
assign M7fhw6 = (C9fhw6 & J9fhw6);
assign J9fhw6 = (Q9fhw6 & X9fhw6);
assign C9fhw6 = (Eafhw6 & Lafhw6);
assign Lafhw6 = (~(Safhw6 & P5fhw6));
assign Safhw6 = (Zafhw6 & Gbfhw6);
assign Eafhw6 = (~(Auehw6 & Nbfhw6));
assign Y6fhw6 = (Ubfhw6 & Bcfhw6);
assign Bcfhw6 = (Icfhw6 & Pcfhw6);
assign Pcfhw6 = (Wcfhw6 & Ddfhw6);
assign Ddfhw6 = (~(Vuehw6 & Kdfhw6));
assign Wcfhw6 = (~(Rdfhw6 & Ydfhw6));
assign Icfhw6 = (Fefhw6 & Mefhw6);
assign Ubfhw6 = (Tefhw6 & Affhw6);
assign Affhw6 = (M0fhw6 ? Offhw6 : Hffhw6);
assign Tefhw6 = (Vffhw6 & Cgfhw6);
assign D6fhw6 = (~(Tfh7z6[1] & W5fhw6));
assign Zaj8v6 = (~(Jgfhw6 & Qgfhw6));
assign Qgfhw6 = (~(Pbadt6 & Vs9ov6));
assign Saj8v6 = (Ehfhw6 ? Xgfhw6 : P4c7z6[0]);
assign Laj8v6 = (Lhfhw6 ? E8h7z6[0] : P4c7z6[0]);
assign Eaj8v6 = (Ehfhw6 ? Shfhw6 : Lvg7z6[3]);
assign X9j8v6 = (Ehfhw6 ? Zhfhw6 : Lvg7z6[2]);
assign Q9j8v6 = (Ehfhw6 ? Gifhw6 : Lvg7z6[1]);
assign J9j8v6 = (Ehfhw6 ? Nifhw6 : Lvg7z6[0]);
assign C9j8v6 = (Ehfhw6 ? Uifhw6 : P4c7z6[3]);
assign V8j8v6 = (Lhfhw6 ? E8h7z6[3] : P4c7z6[3]);
assign O8j8v6 = (Ehfhw6 ? Bjfhw6 : P4c7z6[2]);
assign H8j8v6 = (Lhfhw6 ? E8h7z6[2] : P4c7z6[2]);
assign A8j8v6 = (Ehfhw6 ? Ijfhw6 : P4c7z6[1]);
assign T7j8v6 = (Lhfhw6 ? E8h7z6[1] : P4c7z6[1]);
assign M7j8v6 = (!Pjfhw6);
assign Pjfhw6 = (Kkfhw6 ? Dkfhw6 : Wjfhw6);
assign Dkfhw6 = (Rkfhw6 & Ykfhw6);
assign Ykfhw6 = (~(Flfhw6 & Mlfhw6));
assign Mlfhw6 = (~(Tlfhw6 & Amfhw6));
assign Tlfhw6 = (Hmfhw6 & Omfhw6);
assign Hmfhw6 = (~(Vmfhw6 & Cnfhw6));
assign Cnfhw6 = (Xnfhw6 ? Qnfhw6 : Jnfhw6);
assign Qnfhw6 = (~(Eofhw6 & Lofhw6));
assign Jnfhw6 = (Sofhw6 ? Zec7z6[27] : Zec7z6[25]);
assign Vmfhw6 = (Zofhw6 & Gpfhw6);
assign Gpfhw6 = (~(Npfhw6 & Upfhw6));
assign Upfhw6 = (!Bqfhw6);
assign Flfhw6 = (Wqfhw6 ? Pqfhw6 : Iqfhw6);
assign Pqfhw6 = (Amfhw6 ? Krfhw6 : Drfhw6);
assign Amfhw6 = (!Rrfhw6);
assign Krfhw6 = (Yrfhw6 & Fsfhw6);
assign Fsfhw6 = (~(Msfhw6 & Npfhw6));
assign Yrfhw6 = (Xnfhw6 ? Atfhw6 : Tsfhw6);
assign Atfhw6 = (~(Eofhw6 & Htfhw6));
assign Tsfhw6 = (Sofhw6 ? Vtfhw6 : Otfhw6);
assign Drfhw6 = (Cufhw6 & Jufhw6);
assign Jufhw6 = (~(Qufhw6 & Npfhw6));
assign Cufhw6 = (Xnfhw6 ? Evfhw6 : Xufhw6);
assign Evfhw6 = (~(Lvfhw6 & Eofhw6));
assign Xufhw6 = (Sofhw6 ? Zvfhw6 : Svfhw6);
assign Iqfhw6 = (~(Gwfhw6 & Nwfhw6));
assign Nwfhw6 = (Xnfhw6 ? Bxfhw6 : Uwfhw6);
assign Bxfhw6 = (~(Eofhw6 & Ixfhw6));
assign Uwfhw6 = (~(Pxfhw6 & Sofhw6));
assign Gwfhw6 = (Wxfhw6 & Rrfhw6);
assign Wxfhw6 = (~(Npfhw6 & Dyfhw6));
assign Rkfhw6 = (~(Kyfhw6 & Ryfhw6));
assign Kyfhw6 = (~(Yyfhw6 | Qtnov6));
assign F7j8v6 = (Jgfhw6 ? Ecc7z6[14] : Fzfhw6);
assign Y6j8v6 = (Jgfhw6 ? Ecc7z6[13] : Mzfhw6);
assign R6j8v6 = (Dcnov6 ? Ozbdt6 : Bi9ov6);
assign K6j8v6 = (!Tzfhw6);
assign Tzfhw6 = (Kkfhw6 ? H0ghw6 : A0ghw6);
assign H0ghw6 = (~(O0ghw6 & V0ghw6));
assign V0ghw6 = (C1ghw6 & J1ghw6);
assign C1ghw6 = (Q1ghw6 & Lofhw6);
assign O0ghw6 = (Zec7z6[25] & Auehw6);
assign D6j8v6 = (!X1ghw6);
assign X1ghw6 = (Kkfhw6 ? E2ghw6 : V5jnv6);
assign E2ghw6 = (L2ghw6 & S2ghw6);
assign S2ghw6 = (Z2ghw6 & G3ghw6);
assign Z2ghw6 = (~(N3ghw6 | U3ghw6));
assign L2ghw6 = (B4ghw6 & I4ghw6);
assign V5jnv6 = (!Ecc7z6[11]);
assign W5j8v6 = (~(P4ghw6 & W4ghw6));
assign W4ghw6 = (~(P58et6 & Zs4ov6));
assign P5j8v6 = (~(D5ghw6 & Xr4ov6));
assign D5ghw6 = (K5ghw6 & R5ghw6);
assign R5ghw6 = (~(Bmo8v6 & Ss4ov6));
assign K5ghw6 = (~(Oyh7z6[30] & Zs4ov6));
assign I5j8v6 = (~(Y5ghw6 & Xr4ov6));
assign Y5ghw6 = (F6ghw6 & M6ghw6);
assign M6ghw6 = (~(Zio8v6 & Ss4ov6));
assign F6ghw6 = (~(Oyh7z6[29] & Zs4ov6));
assign B5j8v6 = (~(T6ghw6 & Xr4ov6));
assign T6ghw6 = (A7ghw6 & H7ghw6);
assign H7ghw6 = (~(Xfo8v6 & Ss4ov6));
assign A7ghw6 = (~(Oyh7z6[28] & Zs4ov6));
assign U4j8v6 = (~(O7ghw6 & Xr4ov6));
assign O7ghw6 = (V7ghw6 & C8ghw6);
assign C8ghw6 = (~(Vco8v6 & Ss4ov6));
assign V7ghw6 = (~(Oyh7z6[27] & Zs4ov6));
assign N4j8v6 = (~(J8ghw6 & Xr4ov6));
assign J8ghw6 = (Q8ghw6 & X8ghw6);
assign X8ghw6 = (~(T9o8v6 & Ss4ov6));
assign Q8ghw6 = (~(Oyh7z6[26] & Zs4ov6));
assign G4j8v6 = (~(E9ghw6 & Xr4ov6));
assign E9ghw6 = (L9ghw6 & S9ghw6);
assign S9ghw6 = (~(R6o8v6 & Ss4ov6));
assign L9ghw6 = (~(Oyh7z6[25] & Zs4ov6));
assign Z3j8v6 = (~(Z9ghw6 & Xr4ov6));
assign Z9ghw6 = (Gaghw6 & Naghw6);
assign Naghw6 = (~(P3o8v6 & Ss4ov6));
assign Gaghw6 = (~(Oyh7z6[24] & Zs4ov6));
assign S3j8v6 = (~(Uaghw6 & Xr4ov6));
assign Uaghw6 = (Bbghw6 & Ibghw6);
assign Ibghw6 = (~(N0o8v6 & Ss4ov6));
assign Bbghw6 = (~(Oyh7z6[23] & Zs4ov6));
assign L3j8v6 = (~(Pbghw6 & Xr4ov6));
assign Pbghw6 = (Wbghw6 & Dcghw6);
assign Dcghw6 = (~(Lxn8v6 & Ss4ov6));
assign Wbghw6 = (~(Oyh7z6[22] & Zs4ov6));
assign E3j8v6 = (~(Kcghw6 & Xr4ov6));
assign Kcghw6 = (Rcghw6 & Ycghw6);
assign Ycghw6 = (~(Jun8v6 & Ss4ov6));
assign Rcghw6 = (~(Oyh7z6[21] & Zs4ov6));
assign X2j8v6 = (~(Fdghw6 & Xr4ov6));
assign Fdghw6 = (Mdghw6 & Tdghw6);
assign Tdghw6 = (~(Hrn8v6 & Ss4ov6));
assign Mdghw6 = (~(Oyh7z6[20] & Zs4ov6));
assign Q2j8v6 = (~(Aeghw6 & Xr4ov6));
assign Aeghw6 = (Heghw6 & Oeghw6);
assign Oeghw6 = (~(Fon8v6 & Ss4ov6));
assign Heghw6 = (~(Oyh7z6[19] & Zs4ov6));
assign J2j8v6 = (~(Veghw6 & Xr4ov6));
assign Veghw6 = (Cfghw6 & Jfghw6);
assign Jfghw6 = (~(Dln8v6 & Ss4ov6));
assign Cfghw6 = (~(Oyh7z6[18] & Zs4ov6));
assign C2j8v6 = (~(Qfghw6 & Xr4ov6));
assign Qfghw6 = (Xfghw6 & Egghw6);
assign Egghw6 = (~(Bin8v6 & Ss4ov6));
assign Xfghw6 = (~(Oyh7z6[17] & Zs4ov6));
assign V1j8v6 = (~(Lgghw6 & Xr4ov6));
assign Lgghw6 = (Sgghw6 & Zgghw6);
assign Zgghw6 = (~(Zen8v6 & Ss4ov6));
assign Sgghw6 = (~(Oyh7z6[16] & Zs4ov6));
assign O1j8v6 = (~(Ghghw6 & Xr4ov6));
assign Ghghw6 = (Nhghw6 & Uhghw6);
assign Uhghw6 = (~(Xbn8v6 & Ss4ov6));
assign Nhghw6 = (~(Oyh7z6[15] & Zs4ov6));
assign H1j8v6 = (~(Bighw6 & Xr4ov6));
assign Bighw6 = (Iighw6 & Pighw6);
assign Pighw6 = (~(V8n8v6 & Ss4ov6));
assign Iighw6 = (~(Oyh7z6[14] & Zs4ov6));
assign A1j8v6 = (~(Wighw6 & Xr4ov6));
assign Wighw6 = (Djghw6 & Kjghw6);
assign Kjghw6 = (~(T5n8v6 & Ss4ov6));
assign Djghw6 = (~(Oyh7z6[13] & Zs4ov6));
assign T0j8v6 = (~(Rjghw6 & Xr4ov6));
assign Xr4ov6 = (Fkghw6 ? P4ghw6 : Yjghw6);
assign Rjghw6 = (Mkghw6 & Tkghw6);
assign Tkghw6 = (~(R2n8v6 & Ss4ov6));
assign Mkghw6 = (~(Oyh7z6[12] & Zs4ov6));
assign M0j8v6 = (~(Alghw6 & Hlghw6));
assign Hlghw6 = (~(Oyh7z6[11] & Zs4ov6));
assign Alghw6 = (Olghw6 ? P4ghw6 : Yjghw6);
assign Olghw6 = (Vlghw6 & Cmghw6);
assign Cmghw6 = (~(Pzm8v6 & Jmghw6));
assign Vlghw6 = (Qmghw6 & Fkghw6);
assign Fkghw6 = (~(G4i7z6[9] & Xmghw6));
assign Qmghw6 = (Enghw6 | Lnghw6);
assign F0j8v6 = (~(Snghw6 & Znghw6));
assign Znghw6 = (~(Oyh7z6[10] & Zs4ov6));
assign Snghw6 = (Goghw6 ? P4ghw6 : Yjghw6);
assign Goghw6 = (Noghw6 & Uoghw6);
assign Uoghw6 = (~(Nwm8v6 & Jmghw6));
assign Noghw6 = (Bpghw6 & Ipghw6);
assign Ipghw6 = (Enghw6 | Ppghw6);
assign Bpghw6 = (~(G4i7z6[8] & Xmghw6));
assign Yzi8v6 = (~(Wpghw6 & Dqghw6));
assign Dqghw6 = (~(Oyh7z6[9] & Zs4ov6));
assign Wpghw6 = (Kqghw6 ? P4ghw6 : Yjghw6);
assign Kqghw6 = (Rqghw6 & Yqghw6);
assign Yqghw6 = (~(Mtm8v6 & Jmghw6));
assign Rqghw6 = (Frghw6 & Mrghw6);
assign Mrghw6 = (Enghw6 | Trghw6);
assign Frghw6 = (~(G4i7z6[7] & Xmghw6));
assign Rzi8v6 = (~(Asghw6 & Hsghw6));
assign Hsghw6 = (~(Oyh7z6[8] & Zs4ov6));
assign Asghw6 = (Osghw6 ? P4ghw6 : Yjghw6);
assign Osghw6 = (Vsghw6 & Ctghw6);
assign Ctghw6 = (~(Lqm8v6 & Jmghw6));
assign Vsghw6 = (Jtghw6 & Qtghw6);
assign Qtghw6 = (Enghw6 | Xtghw6);
assign Jtghw6 = (~(G4i7z6[6] & Xmghw6));
assign Kzi8v6 = (~(Eughw6 & Lughw6));
assign Lughw6 = (~(Oyh7z6[7] & Zs4ov6));
assign Eughw6 = (Sughw6 ? P4ghw6 : Yjghw6);
assign Sughw6 = (Zughw6 & Gvghw6);
assign Gvghw6 = (Nvghw6 & Uvghw6);
assign Uvghw6 = (~(Bwghw6 & Q1h7z6[5]));
assign Nvghw6 = (~(Knm8v6 & Jmghw6));
assign Zughw6 = (Iwghw6 & Pwghw6);
assign Pwghw6 = (~(Wwghw6 & Dxghw6));
assign Iwghw6 = (~(G4i7z6[5] & Xmghw6));
assign Dzi8v6 = (~(Kxghw6 & Rxghw6));
assign Rxghw6 = (~(Oyh7z6[6] & Zs4ov6));
assign Kxghw6 = (Yxghw6 ? P4ghw6 : Yjghw6);
assign Yxghw6 = (Fyghw6 & Myghw6);
assign Myghw6 = (Tyghw6 & Azghw6);
assign Azghw6 = (~(G4i7z6[4] & Xmghw6));
assign Tyghw6 = (Hzghw6 & Qsaov6);
assign Hzghw6 = (~(Jkm8v6 & Jmghw6));
assign Fyghw6 = (Ozghw6 & Vzghw6);
assign Vzghw6 = (~(Wwghw6 & C0hhw6));
assign Ozghw6 = (~(Bwghw6 & Q1h7z6[4]));
assign Bwghw6 = (J0hhw6 & Q0hhw6);
assign Wyi8v6 = (~(X0hhw6 & E1hhw6));
assign E1hhw6 = (~(Oyh7z6[5] & Zs4ov6));
assign X0hhw6 = (L1hhw6 ? P4ghw6 : Yjghw6);
assign L1hhw6 = (S1hhw6 & Z1hhw6);
assign Z1hhw6 = (G2hhw6 & N2hhw6);
assign N2hhw6 = (~(G4i7z6[3] & Xmghw6));
assign G2hhw6 = (U2hhw6 & B3hhw6);
assign U2hhw6 = (~(J0hhw6 & I3hhw6));
assign I3hhw6 = (~(P3hhw6 & W3hhw6));
assign W3hhw6 = (~(Q0hhw6 & Q1h7z6[3]));
assign P3hhw6 = (~(Nzg7z6[3] & D4hhw6));
assign S1hhw6 = (K4hhw6 & R4hhw6);
assign R4hhw6 = (Enghw6 | Y4hhw6);
assign K4hhw6 = (F5hhw6 & M5hhw6);
assign M5hhw6 = (~(T5hhw6 & A6hhw6));
assign F5hhw6 = (~(Ihm8v6 & Jmghw6));
assign Pyi8v6 = (~(H6hhw6 & O6hhw6));
assign O6hhw6 = (~(Oyh7z6[4] & Zs4ov6));
assign H6hhw6 = (V6hhw6 ? P4ghw6 : Yjghw6);
assign V6hhw6 = (C7hhw6 & J7hhw6);
assign J7hhw6 = (Q7hhw6 & X7hhw6);
assign X7hhw6 = (~(G4i7z6[2] & Xmghw6));
assign Q7hhw6 = (E8hhw6 & L8hhw6);
assign E8hhw6 = (~(J0hhw6 & S8hhw6));
assign S8hhw6 = (~(Z8hhw6 & G9hhw6));
assign Z8hhw6 = (N9hhw6 & U9hhw6);
assign U9hhw6 = (~(Nzg7z6[2] & D4hhw6));
assign N9hhw6 = (~(Q0hhw6 & Q1h7z6[2]));
assign J0hhw6 = (~(Bahhw6 | Tnzdt6));
assign C7hhw6 = (Iahhw6 & Pahhw6);
assign Pahhw6 = (~(Wwghw6 & Wahhw6));
assign Iahhw6 = (Dbhhw6 & Kbhhw6);
assign Kbhhw6 = (~(T5hhw6 & Rbhhw6));
assign Dbhhw6 = (~(Hem8v6 & Jmghw6));
assign Iyi8v6 = (~(Ybhhw6 & Fchhw6));
assign Fchhw6 = (~(Oyh7z6[3] & Zs4ov6));
assign Ybhhw6 = (Mchhw6 ? P4ghw6 : Yjghw6);
assign Mchhw6 = (Tchhw6 & Adhhw6);
assign Adhhw6 = (Hdhhw6 & Odhhw6);
assign Odhhw6 = (Enghw6 | Vdhhw6);
assign Hdhhw6 = (~(Cehhw6 & T5hhw6));
assign Tchhw6 = (Jehhw6 & Qehhw6);
assign Qehhw6 = (~(Xehhw6 & Efhhw6));
assign Efhhw6 = (~(Lfhhw6 & Sfhhw6));
assign Sfhhw6 = (Zfhhw6 & Gghhw6);
assign Gghhw6 = (Nghhw6 & Ughhw6);
assign Ughhw6 = (~(Hir8v6 & Bhhhw6));
assign Bhhhw6 = (~(Ihhhw6 & Phhhw6));
assign Phhhw6 = (~(Whhhw6 & Dihhw6));
assign Whhhw6 = (~(Kihhw6 | Xumov6));
assign Ihhhw6 = (Rihhw6 | Yihhw6);
assign Nghhw6 = (Fjhhw6 & L8hhw6);
assign Fjhhw6 = (~(Mjhhw6 & Tjhhw6));
assign Tjhhw6 = (~(Akhhw6 & Hkhhw6));
assign Akhhw6 = (Okhhw6 & Vkhhw6);
assign Okhhw6 = (~(Clhhw6 & Aga7z6));
assign Mjhhw6 = (G4i7z6[1] | Jlhhw6);
assign Zfhhw6 = (Qlhhw6 & Xlhhw6);
assign Xlhhw6 = (~(Emhhw6 & Clhhw6));
assign Qlhhw6 = (Hkhhw6 | Iga7z6);
assign Lfhhw6 = (Lmhhw6 & Smhhw6);
assign Smhhw6 = (Zmhhw6 & Gnhhw6);
assign Gnhhw6 = (~(Nzg7z6[1] & D4hhw6));
assign Zmhhw6 = (~(Q0hhw6 & Q1h7z6[1]));
assign Jehhw6 = (~(Gbm8v6 & Jmghw6));
assign Byi8v6 = (~(Nnhhw6 & Unhhw6));
assign Unhhw6 = (~(Oyh7z6[2] & Zs4ov6));
assign Nnhhw6 = (Bohhw6 ? P4ghw6 : Yjghw6);
assign Bohhw6 = (Iohhw6 & Pohhw6);
assign Pohhw6 = (Wohhw6 & Dphhw6);
assign Dphhw6 = (~(Wwghw6 & Kphhw6));
assign Wohhw6 = (~(T5hhw6 & Rphhw6));
assign T5hhw6 = (Yphhw6 & Fqhhw6);
assign Yphhw6 = (Mqhhw6 & Bahhw6);
assign Iohhw6 = (Tqhhw6 & Arhhw6);
assign Arhhw6 = (~(Xehhw6 & Hrhhw6));
assign Hrhhw6 = (~(Orhhw6 & Vrhhw6));
assign Vrhhw6 = (Cshhw6 & Jshhw6);
assign Jshhw6 = (~(Clhhw6 & Lxydt6));
assign Cshhw6 = (Qshhw6 & Xshhw6);
assign Xshhw6 = (~(Ethhw6 & Qg2nv6));
assign Ethhw6 = (~(Lthhw6 & Sthhw6));
assign Sthhw6 = (~(Nzg7z6[0] & D4hhw6));
assign Lthhw6 = (~(Q0hhw6 & Q1h7z6[0]));
assign Qshhw6 = (~(G4i7z6[0] & Xmghw6));
assign Xmghw6 = (~(Zthhw6 | Jlhhw6));
assign Jlhhw6 = (Guhhw6 & Nuhhw6);
assign Nuhhw6 = (~(U6i7z6[1] & Uebdt6));
assign Guhhw6 = (~(U6i7z6[0] & Tnzdt6));
assign Zthhw6 = (Uuhhw6 & Bvhhw6);
assign Bvhhw6 = (Hkhhw6 | Bfo7v6);
assign Uuhhw6 = (Ivhhw6 & Vkhhw6);
assign Ivhhw6 = (~(Clhhw6 & Pvhhw6));
assign Orhhw6 = (Wvhhw6 & Jzaov6);
assign Tqhhw6 = (~(F8m8v6 & Jmghw6));
assign Uxi8v6 = (~(Dwhhw6 & Kwhhw6));
assign Kwhhw6 = (Rwhhw6 ? Yjghw6 : P4ghw6);
assign Rwhhw6 = (Wwghw6 & Ywhhw6);
assign Wwghw6 = (!Enghw6);
assign Dwhhw6 = (Fxhhw6 & Mxhhw6);
assign Mxhhw6 = (~(Txhhw6 & Gvo8v6));
assign Txhhw6 = (Ss4ov6 & Ayhhw6);
assign Ss4ov6 = (Hyhhw6 & Jmghw6);
assign Fxhhw6 = (~(Oyh7z6[1] & Zs4ov6));
assign Nxi8v6 = (~(Oyhhw6 & Vyhhw6));
assign Vyhhw6 = (~(Oyh7z6[0] & Zs4ov6));
assign Oyhhw6 = (Czhhw6 ? P4ghw6 : Yjghw6);
assign Czhhw6 = (Jzhhw6 & Qzhhw6);
assign Qzhhw6 = (Enghw6 | Xzhhw6);
assign Enghw6 = (~(E0ihw6 & L0ihw6));
assign L0ihw6 = (~(Xehhw6 | Xvehw6));
assign Xehhw6 = (!Bahhw6);
assign E0ihw6 = (Fqhhw6 & S0ihw6);
assign Fqhhw6 = (!Z0ihw6);
assign Jzhhw6 = (~(G1ihw6 & Fso8v6));
assign Fso8v6 = (~(Pmknv6 | O7c7z6[7]));
assign O7c7z6[7] = (Uqd7z6[20] & N1ihw6);
assign N1ihw6 = (~(U1ihw6 & B2ihw6));
assign B2ihw6 = (~(I2ihw6 & P2ihw6));
assign I2ihw6 = (N3onv6 & Auehw6);
assign Pmknv6 = (W2ihw6 & D3ihw6);
assign D3ihw6 = (~(K3ihw6 & E7jnv6));
assign K3ihw6 = (~(Q5knv6 | R3ihw6));
assign Q5knv6 = (~(Y3ihw6 | F4ihw6));
assign W2ihw6 = (N8jnv6 | Tefov6);
assign Tefov6 = (M4ihw6 & T4ihw6);
assign T4ihw6 = (A5ihw6 & H5ihw6);
assign H5ihw6 = (O5ihw6 & V5ihw6);
assign V5ihw6 = (C6ihw6 & J6ihw6);
assign J6ihw6 = (~(Pic7z6[0] & U32ov6));
assign C6ihw6 = (~(vis_r12_o[0] & W42ov6));
assign O5ihw6 = (Q6ihw6 & X6ihw6);
assign X6ihw6 = (~(vis_r11_o[0] & F62ov6));
assign Q6ihw6 = (~(vis_r10_o[0] & M62ov6));
assign A5ihw6 = (E7ihw6 & L7ihw6);
assign L7ihw6 = (~(vis_r7_o[0] & L92ov6));
assign E7ihw6 = (S7ihw6 & Z7ihw6);
assign Z7ihw6 = (~(vis_r9_o[0] & H72ov6));
assign S7ihw6 = (~(vis_r8_o[0] & O72ov6));
assign M4ihw6 = (G8ihw6 & N8ihw6);
assign N8ihw6 = (U8ihw6 & B9ihw6);
assign B9ihw6 = (I9ihw6 & P9ihw6);
assign P9ihw6 = (~(vis_r6_o[0] & S92ov6));
assign I9ihw6 = (~(vis_r5_o[0] & Na2ov6));
assign U8ihw6 = (W9ihw6 & Daihw6);
assign Daihw6 = (~(vis_r4_o[0] & Ua2ov6));
assign W9ihw6 = (~(vis_r3_o[0] & Dc2ov6));
assign G8ihw6 = (Kaihw6 & Raihw6);
assign Raihw6 = (~(vis_r0_o[0] & Md2ov6));
assign Kaihw6 = (Yaihw6 & Fbihw6);
assign Fbihw6 = (~(vis_r2_o[0] & Kc2ov6));
assign Yaihw6 = (~(vis_r1_o[0] & Fd2ov6));
assign N8jnv6 = (E7jnv6 | Mbihw6);
assign E7jnv6 = (Tbihw6 & Acihw6);
assign Acihw6 = (Hcihw6 & Ocihw6);
assign Ocihw6 = (~(Vcihw6 ^ F4ihw6));
assign Tbihw6 = (Cdihw6 & Jdihw6);
assign Jdihw6 = (~(Qdihw6 ^ Xdihw6));
assign Cdihw6 = (Eeihw6 & Leihw6);
assign Leihw6 = (~(Seihw6 ^ Zeihw6));
assign Eeihw6 = (~(Gfihw6 ^ Nfihw6));
assign G1ihw6 = (Jmghw6 & Ayhhw6);
assign Ayhhw6 = (!O7c7z6[8]);
assign O7c7z6[8] = (Ufihw6 & Bgihw6);
assign Bgihw6 = (Uqd7z6[21] & Auehw6);
assign Ufihw6 = (P2ihw6 & N3onv6);
assign Jmghw6 = (Igihw6 & Bahhw6);
assign Bahhw6 = (~(Pgihw6 & Wgihw6));
assign Wgihw6 = (Dhihw6 & Khihw6);
assign Khihw6 = (~(Rhihw6 & Qg2nv6));
assign Dhihw6 = (Yhihw6 & Fiihw6);
assign Yhihw6 = (~(Miihw6 & Lxydt6));
assign Miihw6 = (~(Hkhhw6 & Tiihw6));
assign Tiihw6 = (Ajihw6 | Hjihw6);
assign Pgihw6 = (Ojihw6 & Vjihw6);
assign Ojihw6 = (~(Ckihw6 & Jkihw6));
assign Igihw6 = (~(U1ihw6 & Qkihw6));
assign Qkihw6 = (~(Yqvnv6 & Xvehw6));
assign P4ghw6 = (Zs4ov6 | Xkihw6);
assign Yjghw6 = (~(Xkihw6 & Hyhhw6));
assign Xkihw6 = (Elihw6 & Llihw6);
assign Llihw6 = (Slihw6 & Zlihw6);
assign Zlihw6 = (~(Gmihw6 & Zwehw6));
assign Gmihw6 = (Tnzdt6 & Nmihw6);
assign Nmihw6 = (~(Umihw6 & Bnihw6));
assign Bnihw6 = (Inihw6 & Pnihw6);
assign Pnihw6 = (~(Bhoov6 & Dwb7z6[3]));
assign Inihw6 = (~(Wnihw6 | Doihw6));
assign Umihw6 = (Koihw6 & Roihw6);
assign Roihw6 = (Dwb7z6[5] ? Fpihw6 : Yoihw6);
assign Fpihw6 = (~(Ytlnv6 & Mpihw6));
assign Yoihw6 = (Tpihw6 & Mpihw6);
assign Tpihw6 = (~(Dioov6 & Aqihw6));
assign Koihw6 = (Hqihw6 & Oqihw6);
assign Oqihw6 = (~(Nvvnv6 & Bwvnv6));
assign Hqihw6 = (~(Vqihw6 & Gvvnv6));
assign Slihw6 = (Crihw6 & Qsaov6);
assign Crihw6 = (~(Jrihw6 & Qrihw6));
assign Qrihw6 = (~(Xrihw6 | N3ghw6));
assign N3ghw6 = (Ryfhw6 & Zec7z6[7]);
assign Xrihw6 = (U3ghw6 | Esihw6);
assign U3ghw6 = (Lsihw6 & Ssihw6);
assign Ssihw6 = (~(Zsihw6 & Auehw6));
assign Zsihw6 = (Gtihw6 & Xeinv6);
assign Gtihw6 = (~(Rktov6 & Ntihw6));
assign Ntihw6 = (~(Utihw6 & Buihw6));
assign Jrihw6 = (Iuihw6 & B4ghw6);
assign Iuihw6 = (I4ghw6 & G3ghw6);
assign Elihw6 = (Puihw6 & Wuihw6);
assign Wuihw6 = (~(Q0hhw6 & Ecc7z6[11]));
assign Puihw6 = (L8hhw6 | Dwb7z6[5]);
assign Gxi8v6 = (Jgfhw6 ? Ecc7z6[10] : Z0ihw6);
assign Z0ihw6 = (~(Dvihw6 & B4ghw6));
assign B4ghw6 = (Kvihw6 & Rvihw6);
assign Rvihw6 = (~(Zofhw6 & Zec7z6[7]));
assign Kvihw6 = (Yvihw6 & O8fhw6);
assign Dvihw6 = (Fwihw6 & Mwihw6);
assign Mwihw6 = (~(Twihw6 & Axihw6));
assign Twihw6 = (~(Hxihw6 | Zec7z6[26]));
assign Fwihw6 = (~(Ryfhw6 & Bainv6));
assign Zwi8v6 = (Jgfhw6 ? Ecc7z6[9] : Oxihw6);
assign Swi8v6 = (Lhfhw6 ? Whxdt6 : Vxihw6);
assign Lwi8v6 = (Jgfhw6 ? Ecc7z6[6] : Cyihw6);
assign Jgfhw6 = (!Kkfhw6);
assign Ewi8v6 = (~(Jyihw6 & Qyihw6));
assign Qyihw6 = (~(Bh2et6 & Lhfhw6));
assign Xvi8v6 = (~(Xyihw6 & Ezihw6));
assign Ezihw6 = (~(Zdxdt6 & Lzihw6));
assign Lzihw6 = (Ypinv6 | Bqmov6);
assign Xyihw6 = (Eg9ov6 | B3wnv6);
assign Eg9ov6 = (~(Szihw6 & Msmov6));
assign Szihw6 = (Zzihw6 & Bi9ov6);
assign Qvi8v6 = (~(G0jhw6 & N0jhw6));
assign N0jhw6 = (~(U0jhw6 & R3h7z6[0]));
assign Jvi8v6 = (B1jhw6 | I1jhw6);
assign I1jhw6 = (Thbet6 & P1jhw6);
assign Cvi8v6 = (Kkfhw6 ? Mqhhw6 : Ecc7z6[5]);
assign Vui8v6 = (Kkfhw6 ? Yqvnv6 : Ecc7z6[3]);
assign Oui8v6 = (~(W1jhw6 & D2jhw6));
assign D2jhw6 = (~(K2jhw6 & Ubhdt6));
assign Hui8v6 = (Ehfhw6 ? Nfihw6 : Pxg7z6[3]);
assign Aui8v6 = (Ehfhw6 ? Xdihw6 : Pxg7z6[2]);
assign Tti8v6 = (Ehfhw6 ? F4ihw6 : Pxg7z6[1]);
assign Mti8v6 = (Ehfhw6 ? Zeihw6 : Pxg7z6[0]);
assign Fti8v6 = (Uicdt6 ? Y2jhw6 : R2jhw6);
assign Y2jhw6 = (F3jhw6 & M3jhw6);
assign M3jhw6 = (~(T3jhw6 & A4jhw6));
assign F3jhw6 = (Ga3nv6 & X6xnv6);
assign R2jhw6 = (H4jhw6 & Cgc7z6[1]);
assign H4jhw6 = (O4jhw6 & V4jhw6);
assign Ysi8v6 = (Oe2et6 ? Ga3nv6 : Dqnov6);
assign Ksi8v6 = (Udkov6 ? C5jhw6 : Bsgdt6);
assign Dsi8v6 = (Udkov6 ? J5jhw6 : Mpe7z6[4]);
assign Wri8v6 = (Udkov6 ? Q5jhw6 : Mpe7z6[3]);
assign Pri8v6 = (Udkov6 ? X5jhw6 : Mpe7z6[2]);
assign Iri8v6 = (Udkov6 ? E6jhw6 : Xpgdt6);
assign Bri8v6 = (Qf2ov6 ? L6jhw6 : Pne7z6[1]);
assign Uqi8v6 = (Qf2ov6 ? S6jhw6 : Pne7z6[0]);
assign S6jhw6 = (!Bsgdt6);
assign Nqi8v6 = (Z6jhw6 ? D5f7z6[2] : Dknnv6);
assign Gqi8v6 = (Z6jhw6 ? D5f7z6[4] : Pjnnv6);
assign Zpi8v6 = (Z6jhw6 ? D5f7z6[5] : Bjnnv6);
assign Spi8v6 = (Z6jhw6 ? D5f7z6[0] : Rknnv6);
assign Lpi8v6 = (~(G7jhw6 & N7jhw6));
assign N7jhw6 = (U7jhw6 & B8jhw6);
assign B8jhw6 = (~(Okpdt6 & U8bov6));
assign U7jhw6 = (I8jhw6 & P8jhw6);
assign P8jhw6 = (~(Bymdt6 & P9bov6));
assign I8jhw6 = (~(W9bov6 & Onf7z6[28]));
assign G7jhw6 = (W8jhw6 & D9jhw6);
assign D9jhw6 = (~(L0g7z6[28] & Rabov6));
assign W8jhw6 = (K9jhw6 & R9jhw6);
assign R9jhw6 = (~(Vzkdt6 & Mbbov6));
assign K9jhw6 = (~(L0g7z6[12] & Gcmnv6));
assign Epi8v6 = (~(Y9jhw6 & Fajhw6));
assign Fajhw6 = (Majhw6 & Tajhw6);
assign Tajhw6 = (~(Mnpdt6 & U8bov6));
assign Majhw6 = (Abjhw6 & Hbjhw6);
assign Hbjhw6 = (~(A1ndt6 & P9bov6));
assign Abjhw6 = (~(W9bov6 & Onf7z6[27]));
assign Y9jhw6 = (Objhw6 & Vbjhw6);
assign Vbjhw6 = (~(L0g7z6[27] & Rabov6));
assign Objhw6 = (Ccjhw6 & Jcjhw6);
assign Jcjhw6 = (~(Y1ldt6 & Mbbov6));
assign Ccjhw6 = (~(L0g7z6[11] & Gcmnv6));
assign Xoi8v6 = (~(Qcjhw6 & Xcjhw6));
assign Xcjhw6 = (Edjhw6 & Ldjhw6);
assign Ldjhw6 = (~(Kqpdt6 & U8bov6));
assign Edjhw6 = (Sdjhw6 & Zdjhw6);
assign Zdjhw6 = (~(Z3ndt6 & P9bov6));
assign Sdjhw6 = (~(W9bov6 & Onf7z6[26]));
assign Qcjhw6 = (Gejhw6 & Nejhw6);
assign Nejhw6 = (~(L0g7z6[26] & Rabov6));
assign Gejhw6 = (Uejhw6 & Bfjhw6);
assign Bfjhw6 = (~(B4ldt6 & Mbbov6));
assign Uejhw6 = (~(L0g7z6[10] & Gcmnv6));
assign Qoi8v6 = (~(Ifjhw6 & Pfjhw6));
assign Pfjhw6 = (Wfjhw6 & Dgjhw6);
assign Dgjhw6 = (~(Itpdt6 & U8bov6));
assign Wfjhw6 = (Kgjhw6 & Rgjhw6);
assign Rgjhw6 = (~(Y6ndt6 & P9bov6));
assign Kgjhw6 = (~(W9bov6 & Onf7z6[25]));
assign Ifjhw6 = (Ygjhw6 & Fhjhw6);
assign Fhjhw6 = (~(L0g7z6[25] & Rabov6));
assign Ygjhw6 = (Mhjhw6 & Thjhw6);
assign Thjhw6 = (~(E6ldt6 & Mbbov6));
assign Mhjhw6 = (~(L0g7z6[9] & Gcmnv6));
assign Joi8v6 = (~(Aijhw6 & Hijhw6));
assign Hijhw6 = (Oijhw6 & Vijhw6);
assign Vijhw6 = (~(Gwpdt6 & U8bov6));
assign Oijhw6 = (Cjjhw6 & Jjjhw6);
assign Jjjhw6 = (~(X9ndt6 & P9bov6));
assign Cjjhw6 = (~(W9bov6 & Onf7z6[24]));
assign Aijhw6 = (Qjjhw6 & Xjjhw6);
assign Xjjhw6 = (~(L0g7z6[24] & Rabov6));
assign Qjjhw6 = (Ekjhw6 & Lkjhw6);
assign Lkjhw6 = (~(H8ldt6 & Mbbov6));
assign Ekjhw6 = (~(L0g7z6[8] & Gcmnv6));
assign Coi8v6 = (~(Skjhw6 & Zkjhw6));
assign Zkjhw6 = (Gljhw6 & Nljhw6);
assign Nljhw6 = (~(Ezpdt6 & U8bov6));
assign Gljhw6 = (Uljhw6 & Bmjhw6);
assign Bmjhw6 = (~(Wcndt6 & P9bov6));
assign Uljhw6 = (~(W9bov6 & Onf7z6[23]));
assign Skjhw6 = (Imjhw6 & Pmjhw6);
assign Pmjhw6 = (~(L0g7z6[23] & Rabov6));
assign Imjhw6 = (Wmjhw6 & Dnjhw6);
assign Dnjhw6 = (~(Kaldt6 & Mbbov6));
assign Wmjhw6 = (~(L0g7z6[7] & Gcmnv6));
assign Vni8v6 = (~(Knjhw6 & Rnjhw6));
assign Rnjhw6 = (Ynjhw6 & Fojhw6);
assign Fojhw6 = (~(C2qdt6 & U8bov6));
assign Ynjhw6 = (Mojhw6 & Tojhw6);
assign Tojhw6 = (~(Vfndt6 & P9bov6));
assign Mojhw6 = (~(W9bov6 & Onf7z6[22]));
assign Knjhw6 = (Apjhw6 & Hpjhw6);
assign Hpjhw6 = (~(L0g7z6[22] & Rabov6));
assign Apjhw6 = (Opjhw6 & Vpjhw6);
assign Vpjhw6 = (~(Ncldt6 & Mbbov6));
assign Opjhw6 = (~(L0g7z6[6] & Gcmnv6));
assign Oni8v6 = (~(Cqjhw6 & Jqjhw6));
assign Jqjhw6 = (Qqjhw6 & Xqjhw6);
assign Xqjhw6 = (~(A5qdt6 & U8bov6));
assign Qqjhw6 = (Erjhw6 & Lrjhw6);
assign Lrjhw6 = (~(Uindt6 & P9bov6));
assign Erjhw6 = (~(W9bov6 & Onf7z6[21]));
assign Cqjhw6 = (Srjhw6 & Zrjhw6);
assign Zrjhw6 = (~(L0g7z6[21] & Rabov6));
assign Srjhw6 = (Gsjhw6 & Nsjhw6);
assign Nsjhw6 = (~(Qeldt6 & Mbbov6));
assign Gsjhw6 = (~(L0g7z6[5] & Gcmnv6));
assign Hni8v6 = (~(Usjhw6 & Btjhw6));
assign Btjhw6 = (Itjhw6 & Ptjhw6);
assign Ptjhw6 = (~(Y7qdt6 & U8bov6));
assign Itjhw6 = (Wtjhw6 & Dujhw6);
assign Dujhw6 = (~(Tlndt6 & P9bov6));
assign Wtjhw6 = (~(W9bov6 & Onf7z6[20]));
assign Usjhw6 = (Kujhw6 & Rujhw6);
assign Rujhw6 = (~(L0g7z6[20] & Rabov6));
assign Kujhw6 = (Yujhw6 & Fvjhw6);
assign Fvjhw6 = (~(Tgldt6 & Mbbov6));
assign Yujhw6 = (~(L0g7z6[4] & Gcmnv6));
assign Ani8v6 = (~(Mvjhw6 & Tvjhw6));
assign Tvjhw6 = (Awjhw6 & Hwjhw6);
assign Hwjhw6 = (~(Waqdt6 & U8bov6));
assign Awjhw6 = (Owjhw6 & Vwjhw6);
assign Vwjhw6 = (~(Sondt6 & P9bov6));
assign Owjhw6 = (~(W9bov6 & Onf7z6[19]));
assign Mvjhw6 = (Cxjhw6 & Jxjhw6);
assign Jxjhw6 = (~(L0g7z6[19] & Rabov6));
assign Cxjhw6 = (Qxjhw6 & Xxjhw6);
assign Xxjhw6 = (~(Wildt6 & Mbbov6));
assign Qxjhw6 = (~(L0g7z6[3] & Gcmnv6));
assign Tmi8v6 = (~(Eyjhw6 & Lyjhw6));
assign Lyjhw6 = (Syjhw6 & Zyjhw6);
assign Zyjhw6 = (~(Udqdt6 & U8bov6));
assign Syjhw6 = (Gzjhw6 & Nzjhw6);
assign Nzjhw6 = (~(Rrndt6 & P9bov6));
assign Gzjhw6 = (~(W9bov6 & Onf7z6[18]));
assign Eyjhw6 = (Uzjhw6 & B0khw6);
assign B0khw6 = (~(L0g7z6[18] & Rabov6));
assign Uzjhw6 = (I0khw6 & P0khw6);
assign P0khw6 = (~(Zkldt6 & Mbbov6));
assign I0khw6 = (~(L0g7z6[2] & Gcmnv6));
assign Mmi8v6 = (~(W0khw6 & D1khw6));
assign D1khw6 = (K1khw6 & R1khw6);
assign R1khw6 = (~(Sgqdt6 & U8bov6));
assign K1khw6 = (Y1khw6 & F2khw6);
assign F2khw6 = (~(Qundt6 & P9bov6));
assign Y1khw6 = (~(W9bov6 & Onf7z6[17]));
assign W0khw6 = (M2khw6 & T2khw6);
assign T2khw6 = (~(L0g7z6[17] & Rabov6));
assign M2khw6 = (A3khw6 & H3khw6);
assign H3khw6 = (~(Cnldt6 & Mbbov6));
assign A3khw6 = (~(L0g7z6[1] & Gcmnv6));
assign Fmi8v6 = (~(O3khw6 & V3khw6));
assign V3khw6 = (C4khw6 & J4khw6);
assign J4khw6 = (~(Qjqdt6 & U8bov6));
assign C4khw6 = (Q4khw6 & X4khw6);
assign X4khw6 = (~(Pxndt6 & P9bov6));
assign Q4khw6 = (~(W9bov6 & Onf7z6[16]));
assign O3khw6 = (E5khw6 & L5khw6);
assign L5khw6 = (~(L0g7z6[16] & Rabov6));
assign E5khw6 = (S5khw6 & Z5khw6);
assign Z5khw6 = (~(Fpldt6 & Mbbov6));
assign S5khw6 = (~(L0g7z6[0] & Gcmnv6));
assign Yli8v6 = (~(G6khw6 & N6khw6));
assign N6khw6 = (U6khw6 & B7khw6);
assign B7khw6 = (~(Omqdt6 & U8bov6));
assign U6khw6 = (I7khw6 & P7khw6);
assign P7khw6 = (~(O0odt6 & P9bov6));
assign I7khw6 = (~(Onf7z6[15] & Ohkov6));
assign G6khw6 = (W7khw6 & D8khw6);
assign D8khw6 = (~(Irldt6 & Mbbov6));
assign W7khw6 = (~(L0g7z6[15] & Rabov6));
assign Rli8v6 = (~(K8khw6 & R8khw6));
assign R8khw6 = (Y8khw6 & F9khw6);
assign F9khw6 = (~(Mpqdt6 & U8bov6));
assign Y8khw6 = (M9khw6 & T9khw6);
assign T9khw6 = (~(N3odt6 & P9bov6));
assign M9khw6 = (~(Onf7z6[14] & Ohkov6));
assign K8khw6 = (Aakhw6 & Hakhw6);
assign Hakhw6 = (~(Ltldt6 & Mbbov6));
assign Aakhw6 = (~(L0g7z6[14] & Rabov6));
assign Kli8v6 = (~(Oakhw6 & Vakhw6));
assign Vakhw6 = (Cbkhw6 & Jbkhw6);
assign Jbkhw6 = (~(Ksqdt6 & U8bov6));
assign Cbkhw6 = (Qbkhw6 & Xbkhw6);
assign Xbkhw6 = (~(M6odt6 & P9bov6));
assign Qbkhw6 = (~(Onf7z6[13] & Ohkov6));
assign Oakhw6 = (Eckhw6 & Lckhw6);
assign Lckhw6 = (~(Ovldt6 & Mbbov6));
assign Eckhw6 = (~(L0g7z6[13] & Rabov6));
assign Dli8v6 = (~(Sckhw6 & Zckhw6));
assign Zckhw6 = (Gdkhw6 & Ndkhw6);
assign Ndkhw6 = (~(Ivqdt6 & U8bov6));
assign Gdkhw6 = (Udkhw6 & Bekhw6);
assign Bekhw6 = (~(L9odt6 & P9bov6));
assign Udkhw6 = (~(Onf7z6[12] & Ohkov6));
assign Sckhw6 = (Iekhw6 & Pekhw6);
assign Pekhw6 = (~(Rxldt6 & Mbbov6));
assign Iekhw6 = (~(L0g7z6[12] & Rabov6));
assign Wki8v6 = (~(Wekhw6 & Dfkhw6));
assign Dfkhw6 = (Kfkhw6 & Rfkhw6);
assign Rfkhw6 = (~(Gyqdt6 & U8bov6));
assign Kfkhw6 = (Yfkhw6 & Fgkhw6);
assign Fgkhw6 = (~(Kcodt6 & P9bov6));
assign Yfkhw6 = (~(Onf7z6[11] & Ohkov6));
assign Wekhw6 = (Mgkhw6 & Tgkhw6);
assign Tgkhw6 = (~(Uzldt6 & Mbbov6));
assign Mgkhw6 = (~(L0g7z6[11] & Rabov6));
assign Pki8v6 = (~(Ahkhw6 & Hhkhw6));
assign Hhkhw6 = (Ohkhw6 & Vhkhw6);
assign Vhkhw6 = (~(E1rdt6 & U8bov6));
assign Ohkhw6 = (Cikhw6 & Jikhw6);
assign Jikhw6 = (~(Jfodt6 & P9bov6));
assign Cikhw6 = (~(Onf7z6[10] & Ohkov6));
assign Ahkhw6 = (Qikhw6 & Xikhw6);
assign Xikhw6 = (~(X1mdt6 & Mbbov6));
assign Qikhw6 = (~(L0g7z6[10] & Rabov6));
assign Iki8v6 = (~(Ejkhw6 & Ljkhw6));
assign Ljkhw6 = (Sjkhw6 & Zjkhw6);
assign Zjkhw6 = (~(C4rdt6 & U8bov6));
assign Sjkhw6 = (Gkkhw6 & Nkkhw6);
assign Nkkhw6 = (~(Iiodt6 & P9bov6));
assign Gkkhw6 = (~(Onf7z6[9] & Ohkov6));
assign Ejkhw6 = (Ukkhw6 & Blkhw6);
assign Blkhw6 = (~(A4mdt6 & Mbbov6));
assign Ukkhw6 = (~(L0g7z6[9] & Rabov6));
assign Bki8v6 = (~(Ilkhw6 & Plkhw6));
assign Plkhw6 = (Wlkhw6 & Dmkhw6);
assign Dmkhw6 = (~(A7rdt6 & U8bov6));
assign Wlkhw6 = (Kmkhw6 & Rmkhw6);
assign Rmkhw6 = (~(Hlodt6 & P9bov6));
assign Kmkhw6 = (~(Onf7z6[8] & Ohkov6));
assign Ilkhw6 = (Ymkhw6 & Fnkhw6);
assign Fnkhw6 = (~(D6mdt6 & Mbbov6));
assign Ymkhw6 = (~(L0g7z6[8] & Rabov6));
assign Uji8v6 = (~(Mnkhw6 & Tnkhw6));
assign Tnkhw6 = (Aokhw6 & Hokhw6);
assign Hokhw6 = (~(Y9rdt6 & U8bov6));
assign Aokhw6 = (Ookhw6 & Vokhw6);
assign Vokhw6 = (~(Goodt6 & P9bov6));
assign Ookhw6 = (~(Onf7z6[7] & Ohkov6));
assign Mnkhw6 = (Cpkhw6 & Jpkhw6);
assign Jpkhw6 = (~(G8mdt6 & Mbbov6));
assign Cpkhw6 = (~(L0g7z6[7] & Rabov6));
assign Nji8v6 = (~(Qpkhw6 & Xpkhw6));
assign Xpkhw6 = (Eqkhw6 & Lqkhw6);
assign Lqkhw6 = (~(Wcrdt6 & U8bov6));
assign Eqkhw6 = (Sqkhw6 & Zqkhw6);
assign Zqkhw6 = (~(Frodt6 & P9bov6));
assign Sqkhw6 = (~(Onf7z6[6] & Ohkov6));
assign Qpkhw6 = (Grkhw6 & Nrkhw6);
assign Nrkhw6 = (~(Jamdt6 & Mbbov6));
assign Grkhw6 = (~(L0g7z6[6] & Rabov6));
assign Gji8v6 = (~(Urkhw6 & Bskhw6));
assign Bskhw6 = (Iskhw6 & Pskhw6);
assign Pskhw6 = (~(Ufrdt6 & U8bov6));
assign Iskhw6 = (Wskhw6 & Dtkhw6);
assign Dtkhw6 = (~(Euodt6 & P9bov6));
assign Wskhw6 = (~(Onf7z6[5] & Ohkov6));
assign Urkhw6 = (Ktkhw6 & Rtkhw6);
assign Rtkhw6 = (~(Mcmdt6 & Mbbov6));
assign Ktkhw6 = (~(L0g7z6[5] & Rabov6));
assign Zii8v6 = (~(Ytkhw6 & Fukhw6));
assign Fukhw6 = (Mukhw6 & Tukhw6);
assign Tukhw6 = (~(Sirdt6 & U8bov6));
assign Mukhw6 = (Avkhw6 & Hvkhw6);
assign Hvkhw6 = (~(Dxodt6 & P9bov6));
assign Avkhw6 = (~(Onf7z6[4] & Ohkov6));
assign Ytkhw6 = (Ovkhw6 & Vvkhw6);
assign Vvkhw6 = (~(Pemdt6 & Mbbov6));
assign Ovkhw6 = (~(L0g7z6[4] & Rabov6));
assign Sii8v6 = (~(Cwkhw6 & Jwkhw6));
assign Jwkhw6 = (Qwkhw6 & Xwkhw6);
assign Xwkhw6 = (~(Qlrdt6 & U8bov6));
assign Qwkhw6 = (Exkhw6 & Lxkhw6);
assign Lxkhw6 = (~(C0pdt6 & P9bov6));
assign Exkhw6 = (~(Onf7z6[3] & Ohkov6));
assign Cwkhw6 = (Sxkhw6 & Zxkhw6);
assign Zxkhw6 = (~(Sgmdt6 & Mbbov6));
assign Sxkhw6 = (~(L0g7z6[3] & Rabov6));
assign Lii8v6 = (~(Gykhw6 & Nykhw6));
assign Nykhw6 = (Uykhw6 & Bzkhw6);
assign Bzkhw6 = (~(Oordt6 & U8bov6));
assign Uykhw6 = (Izkhw6 & Pzkhw6);
assign Pzkhw6 = (~(A3pdt6 & P9bov6));
assign Izkhw6 = (~(Onf7z6[2] & Ohkov6));
assign Gykhw6 = (Wzkhw6 & D0lhw6);
assign D0lhw6 = (~(Vimdt6 & Mbbov6));
assign Wzkhw6 = (~(L0g7z6[2] & Rabov6));
assign Eii8v6 = (~(K0lhw6 & R0lhw6));
assign R0lhw6 = (Y0lhw6 & F1lhw6);
assign F1lhw6 = (~(Mrrdt6 & U8bov6));
assign U8bov6 = (M1lhw6 & T1lhw6);
assign Y0lhw6 = (A2lhw6 & H2lhw6);
assign H2lhw6 = (~(Y5pdt6 & P9bov6));
assign P9bov6 = (M1lhw6 & O2lhw6);
assign O2lhw6 = (!T1lhw6);
assign A2lhw6 = (~(Onf7z6[1] & Ohkov6));
assign Ohkov6 = (Gcmnv6 | W9bov6);
assign W9bov6 = (V2lhw6 & C3lhw6);
assign C3lhw6 = (~(M1lhw6 | Rabov6));
assign V2lhw6 = (~(Mbbov6 | Gcmnv6));
assign K0lhw6 = (J3lhw6 & Q3lhw6);
assign Q3lhw6 = (~(Ykmdt6 & Mbbov6));
assign Mbbov6 = (~(X3lhw6 & E4lhw6));
assign J3lhw6 = (~(L0g7z6[1] & Rabov6));
assign Xhi8v6 = (Ehfhw6 ? L4lhw6 : Ntg7z6[3]);
assign Qhi8v6 = (Efhov6 ? L4lhw6 : Oac7z6[3]);
assign Jhi8v6 = (Ehfhw6 ? S4lhw6 : Ntg7z6[2]);
assign Chi8v6 = (Efhov6 ? S4lhw6 : Oac7z6[2]);
assign Efhov6 = (!K2jhw6);
assign Vgi8v6 = (Ehfhw6 ? Xehov6 : Ntg7z6[1]);
assign Ogi8v6 = (~(Z4lhw6 & G5lhw6));
assign G5lhw6 = (~(Z8c7z6[0] & Vs9ov6));
assign Z4lhw6 = (N5lhw6 & U5lhw6);
assign U5lhw6 = (~(B6lhw6 & I6lhw6));
assign N5lhw6 = (~(P6lhw6 & Nifhw6));
assign Hgi8v6 = (~(W6lhw6 & D7lhw6));
assign D7lhw6 = (~(Z8c7z6[1] & Vs9ov6));
assign W6lhw6 = (K7lhw6 & R7lhw6);
assign R7lhw6 = (~(B6lhw6 & Xehov6));
assign K7lhw6 = (~(P6lhw6 & Gifhw6));
assign Agi8v6 = (~(Y7lhw6 & F8lhw6));
assign F8lhw6 = (~(Z8c7z6[2] & Vs9ov6));
assign Y7lhw6 = (M8lhw6 & T8lhw6);
assign T8lhw6 = (~(B6lhw6 & S4lhw6));
assign M8lhw6 = (~(P6lhw6 & Zhfhw6));
assign Tfi8v6 = (~(A9lhw6 & H9lhw6));
assign H9lhw6 = (~(Z8c7z6[3] & Vs9ov6));
assign A9lhw6 = (O9lhw6 & V9lhw6);
assign V9lhw6 = (~(B6lhw6 & L4lhw6));
assign B6lhw6 = (~(Vs9ov6 | P6lhw6));
assign O9lhw6 = (~(P6lhw6 & Shfhw6));
assign Mfi8v6 = (Ehfhw6 ? I6lhw6 : Ntg7z6[0]);
assign Ehfhw6 = (Kkfhw6 & Calhw6);
assign Kkfhw6 = (Snvnv6 & Jalhw6);
assign Jalhw6 = (Qalhw6 | Fzfhw6);
assign Ffi8v6 = (~(Xalhw6 & Eblhw6));
assign Eblhw6 = (~(O5h7z6[0] & Lhfhw6));
assign Xalhw6 = (Lblhw6 & Sblhw6);
assign Sblhw6 = (~(Zblhw6 & Lvg7z6[0]));
assign Lblhw6 = (Jyihw6 | Gclhw6);
assign Yei8v6 = (~(Nclhw6 & Uclhw6));
assign Uclhw6 = (~(O5h7z6[1] & Lhfhw6));
assign Nclhw6 = (Bdlhw6 & Idlhw6);
assign Idlhw6 = (~(Zblhw6 & Lvg7z6[1]));
assign Bdlhw6 = (Jyihw6 | Pdlhw6);
assign Rei8v6 = (~(Wdlhw6 & Delhw6));
assign Delhw6 = (~(O5h7z6[2] & Lhfhw6));
assign Wdlhw6 = (Kelhw6 & Relhw6);
assign Relhw6 = (~(Zblhw6 & Lvg7z6[2]));
assign Kelhw6 = (Jyihw6 | Yelhw6);
assign Kei8v6 = (~(Fflhw6 & Mflhw6));
assign Mflhw6 = (~(O5h7z6[3] & Lhfhw6));
assign Fflhw6 = (Tflhw6 & Aglhw6);
assign Aglhw6 = (~(Zblhw6 & Lvg7z6[3]));
assign Zblhw6 = (~(Lhfhw6 | Zzihw6));
assign Lhfhw6 = (!Hglhw6);
assign Tflhw6 = (Jyihw6 | Oglhw6);
assign Jyihw6 = (~(Hglhw6 & Zzihw6));
assign Hglhw6 = (Gr2et6 & Vglhw6);
assign Dei8v6 = (K2jhw6 ? Oac7z6[0] : I6lhw6);
assign K2jhw6 = (W1jhw6 & Chlhw6);
assign Chlhw6 = (~(Ubhdt6 & Jhlhw6));
assign Jhlhw6 = (~(Qhlhw6 & Dcnov6));
assign Qhlhw6 = (~(Xhlhw6 & Ixfov6));
assign W1jhw6 = (~(N3onv6 & Eilhw6));
assign Wdi8v6 = (Trnov6 & Lilhw6);
assign Lilhw6 = (Silhw6 | Zilhw6);
assign Pdi8v6 = (~(Gjlhw6 & Njlhw6));
assign Njlhw6 = (~(Ujlhw6 & Frnov6));
assign Frnov6 = (Bklhw6 & C0wnv6);
assign Ujlhw6 = (Qyddt6 & Mrnov6);
assign Gjlhw6 = (~(Trnov6 & Iklhw6));
assign Iklhw6 = (~(Pklhw6 & Wklhw6));
assign Wklhw6 = (~(Vsnov6 & Ovbdt6));
assign Pklhw6 = (~(Jtnov6 & Zec7z6[4]));
assign Idi8v6 = (Pyeov6 ? Dllhw6 : R7fet6);
assign Dllhw6 = (!Lunov6);
assign Bdi8v6 = (Kllhw6 & Rllhw6);
assign Rllhw6 = (Yllhw6 & Fmlhw6);
assign Fmlhw6 = (Mmlhw6 & Tmlhw6);
assign Tmlhw6 = (Anlhw6 & Hnlhw6);
assign Hnlhw6 = (Onlhw6 & Vnlhw6);
assign Anlhw6 = (W4onv6 & Hffhw6);
assign Mmlhw6 = (~(Colhw6 | Mtsov6));
assign Mtsov6 = (Jolhw6 & Qolhw6);
assign Colhw6 = (Jhsov6 | Xolhw6);
assign Yllhw6 = (Eplhw6 & Lplhw6);
assign Lplhw6 = (Splhw6 & F0fhw6);
assign Splhw6 = (Zplhw6 & Calhw6);
assign Calhw6 = (!Fzfhw6);
assign Fzfhw6 = (Gqlhw6 & Nqlhw6);
assign Eplhw6 = (Uqlhw6 & I4ghw6);
assign Uqlhw6 = (Brlhw6 & Irlhw6);
assign Irlhw6 = (~(Prlhw6 & Zec7z6[10]));
assign Prlhw6 = (Wrlhw6 & Dslhw6);
assign Wrlhw6 = (~(Zec7z6[9] & Zec7z6[8]));
assign Kllhw6 = (Kslhw6 & Rslhw6);
assign Rslhw6 = (Yslhw6 & Ftlhw6);
assign Ftlhw6 = (Mtlhw6 & Ttlhw6);
assign Ttlhw6 = (Aulhw6 & Hulhw6);
assign Mtlhw6 = (Oulhw6 & Vulhw6);
assign Yslhw6 = (Cvlhw6 & Jvlhw6);
assign Cvlhw6 = (Qvlhw6 & Xvlhw6);
assign Kslhw6 = (Ewlhw6 & Lwlhw6);
assign Lwlhw6 = (~(Swlhw6 | Zwlhw6));
assign Swlhw6 = (Gxlhw6 | Nxlhw6);
assign Ewlhw6 = (Uxlhw6 & Bylhw6);
assign Uxlhw6 = (Iylhw6 & Trnov6);
assign Uci8v6 = (~(Pylhw6 & Wylhw6));
assign Wylhw6 = (~(Bfd7z6[0] & M8mnv6));
assign Pylhw6 = (Dzlhw6 & Kzlhw6);
assign Kzlhw6 = (~(Rzlhw6 & W6mnv6));
assign W6mnv6 = (~(Yzlhw6 & F0mhw6));
assign F0mhw6 = (M0mhw6 & Iwnov6);
assign M0mhw6 = (~(T0mhw6 & A1mhw6));
assign T0mhw6 = (H1mhw6 ? Bfd7z6[4] : Bfd7z6[5]);
assign Yzlhw6 = (O1mhw6 & V1mhw6);
assign V1mhw6 = (~(F8mnv6 & Kboov6));
assign O1mhw6 = (C2mhw6 | Pdc7z6[1]);
assign Dzlhw6 = (~(F8mnv6 & U5mnv6));
assign Nci8v6 = (~(J2mhw6 & Q2mhw6));
assign Q2mhw6 = (K0mnv6 | D7mnv6);
assign K0mnv6 = (~(X2mhw6 & A1mhw6));
assign X2mhw6 = (H1mhw6 ? Bfd7z6[3] : Bfd7z6[4]);
assign J2mhw6 = (~(M8mnv6 & Bfd7z6[5]));
assign Gci8v6 = (~(E3mhw6 & L3mhw6));
assign L3mhw6 = (~(M1mnv6 & Rzlhw6));
assign M1mnv6 = (S3mhw6 & A1mhw6);
assign S3mhw6 = (H1mhw6 ? Bfd7z6[2] : Bfd7z6[3]);
assign E3mhw6 = (~(Bfd7z6[4] & M8mnv6));
assign Zbi8v6 = (~(Z3mhw6 & G4mhw6));
assign G4mhw6 = (C3mnv6 | D7mnv6);
assign C3mnv6 = (~(N4mhw6 & A1mhw6));
assign N4mhw6 = (H1mhw6 ? Bfd7z6[1] : Bfd7z6[2]);
assign Z3mhw6 = (~(M8mnv6 & Bfd7z6[3]));
assign Sbi8v6 = (~(U4mhw6 & B5mhw6));
assign B5mhw6 = (X3mnv6 | D7mnv6);
assign X3mnv6 = (~(I5mhw6 & A1mhw6));
assign I5mhw6 = (H1mhw6 ? Bfd7z6[0] : Bfd7z6[1]);
assign U4mhw6 = (~(Bfd7z6[2] & M8mnv6));
assign Lbi8v6 = (~(P5mhw6 & W5mhw6));
assign W5mhw6 = (~(M8mnv6 & Bfd7z6[1]));
assign P5mhw6 = (D6mhw6 & K6mhw6);
assign K6mhw6 = (D7mnv6 | S4mnv6);
assign S4mnv6 = (R6mhw6 & Y6mhw6);
assign Y6mhw6 = (~(Pdc7z6[1] & F7mhw6));
assign R6mhw6 = (M7mhw6 & T7mhw6);
assign T7mhw6 = (~(A8mhw6 & A1mhw6));
assign A8mhw6 = (H1mhw6 ? Bfd7z6[5] : Bfd7z6[0]);
assign H1mhw6 = (~(H8mhw6 | Tao7v6));
assign H8mhw6 = (!Yiaov6);
assign M7mhw6 = (~(Kboov6 & B6mnv6));
assign D7mnv6 = (!Rzlhw6);
assign Rzlhw6 = (~(U5mnv6 | M8mnv6));
assign M8mnv6 = (D61ov6 & O8mhw6);
assign O8mhw6 = (~(K6tov6 & V8mhw6));
assign V8mhw6 = (~(C9mhw6 & Pacdt6));
assign C9mhw6 = (C2mhw6 & Iwnov6);
assign K6tov6 = (~(J9mhw6 & C2mhw6));
assign C2mhw6 = (!F7mhw6);
assign F7mhw6 = (~(Q9mhw6 & Z8oov6));
assign Q9mhw6 = (~(X9mhw6 & Iwnov6));
assign J9mhw6 = (Eamhw6 & Iwnov6);
assign Iwnov6 = (~(X9mhw6 & A4jhw6));
assign Eamhw6 = (~(N3onv6 & A1mhw6));
assign A1mhw6 = (!Lamhw6);
assign D6mhw6 = (~(U5mnv6 & B6mnv6));
assign B6mnv6 = (!F8mnv6);
assign F8mnv6 = (Samhw6 & Zamhw6);
assign Zamhw6 = (Qdcdt6 ? Nbmhw6 : Gbmhw6);
assign Nbmhw6 = (~(Lp0ov6 & E3c7z6[1]));
assign Gbmhw6 = (~(Ubmhw6 & Bcmhw6));
assign Bcmhw6 = (Icmhw6 & Pcmhw6);
assign Icmhw6 = (Wkd7z6[1] | Jamnv6);
assign Ubmhw6 = (Lp0ov6 & Wcmhw6);
assign Wcmhw6 = (Vnd7z6[1] | Ddmhw6);
assign Samhw6 = (Lp0ov6 ? Rdmhw6 : Kdmhw6);
assign Lp0ov6 = (Af1ov6 & Gpmov6);
assign Rdmhw6 = (~(Pic7z6[1] & Ir0ov6));
assign U5mnv6 = (~(Lamhw6 | D61ov6));
assign Lamhw6 = (Cgc7z6[3] ? Cgc7z6[1] : Ydmhw6);
assign Ebi8v6 = (~(Femhw6 & Memhw6));
assign Memhw6 = (~(Riaov6 & Lpc7z6[0]));
assign Xai8v6 = (~(Temhw6 & Afmhw6));
assign Afmhw6 = (~(Hfmhw6 & Snvnv6));
assign Hfmhw6 = (~(Ofmhw6 | Pacdt6));
assign Temhw6 = (~(Vfmhw6 & Efcdt6));
assign Vfmhw6 = (Qv0ov6 & X6xnv6);
assign Qai8v6 = (~(Brlhw6 | Cgmhw6));
assign Cgmhw6 = (!Trnov6);
assign Brlhw6 = (~(Jgmhw6 & Qgmhw6));
assign Qgmhw6 = (Zec7z6[12] & Zec7z6[8]);
assign Jgmhw6 = (Z3fhw6 & Xgmhw6);
assign Cai8v6 = (Ehmhw6 & Trnov6);
assign Ehmhw6 = (Lhmhw6 & Dslhw6);
assign Dslhw6 = (Shmhw6 | Zhmhw6);
assign Lhmhw6 = (Gbfhw6 | Gimhw6);
assign Gimhw6 = (~(Painv6 | Zec7z6[8]));
assign O9i8v6 = (Nimhw6 & Uimhw6);
assign Uimhw6 = (Tuddt6 | Bjmhw6);
assign Bjmhw6 = (Ffadt6 & Lamov6);
assign Lamov6 = (Tnzdt6 | Etinv6);
assign Nimhw6 = (Samov6 & Ijmhw6);
assign Samov6 = (~(Dj9ov6 & O5a7z6));
assign H9i8v6 = (~(Pjmhw6 | V9i8v6));
assign Pjmhw6 = (Vs9ov6 & Wjmhw6);
assign Wjmhw6 = (~(Dkmhw6 & Oaadt6));
assign Dkmhw6 = (Wpvnv6 & Kkmhw6);
assign Wpvnv6 = (~(Rkmhw6 & Ykmhw6));
assign Ykmhw6 = (Flmhw6 & Q0wnv6);
assign Flmhw6 = (~(Dj9ov6 | S1wnv6));
assign Rkmhw6 = (C9mov6 & Mlmhw6);
assign T8i8v6 = (!Tlmhw6);
assign Tlmhw6 = (Ammhw6 ? Xzhhw6 : J6jnv6);
assign M8i8v6 = (~(Hmmhw6 & Ommhw6));
assign Ommhw6 = (Vmmhw6 & Cnmhw6);
assign Cnmhw6 = (~(Jnmhw6 & Uqd7z6[20]));
assign Vmmhw6 = (Qnmhw6 & Xnmhw6);
assign Qnmhw6 = (~(Eomhw6 & Lomhw6));
assign Hmmhw6 = (Somhw6 & Zomhw6);
assign Zomhw6 = (~(V1c7z6[31] & Gpmhw6));
assign Somhw6 = (Npmhw6 & Upmhw6);
assign Upmhw6 = (~(Bqmhw6 & Zec7z6[3]));
assign F8i8v6 = (~(Iqmhw6 & Pqmhw6));
assign Pqmhw6 = (Wqmhw6 & Drmhw6);
assign Drmhw6 = (~(Jnmhw6 & Uqd7z6[19]));
assign Wqmhw6 = (Krmhw6 & Xnmhw6);
assign Krmhw6 = (~(Rrmhw6 & Eomhw6));
assign Iqmhw6 = (Yrmhw6 & Fsmhw6);
assign Fsmhw6 = (~(V1c7z6[30] & Gpmhw6));
assign Yrmhw6 = (Msmhw6 & Tsmhw6);
assign Tsmhw6 = (~(Bqmhw6 & Zec7z6[2]));
assign Y7i8v6 = (~(Atmhw6 & Htmhw6));
assign Htmhw6 = (Otmhw6 & Vtmhw6);
assign Vtmhw6 = (~(Jnmhw6 & Uqd7z6[18]));
assign Otmhw6 = (Cumhw6 & Xnmhw6);
assign Cumhw6 = (~(Jumhw6 & Eomhw6));
assign Atmhw6 = (Qumhw6 & Xumhw6);
assign Xumhw6 = (~(V1c7z6[29] & Gpmhw6));
assign Qumhw6 = (Evmhw6 & Lvmhw6);
assign Lvmhw6 = (~(Bqmhw6 & Zec7z6[1]));
assign R7i8v6 = (~(Svmhw6 & Zvmhw6));
assign Zvmhw6 = (Gwmhw6 & Nwmhw6);
assign Nwmhw6 = (~(Jnmhw6 & Uqd7z6[17]));
assign Gwmhw6 = (Uwmhw6 & Xnmhw6);
assign Uwmhw6 = (~(Bxmhw6 & Eomhw6));
assign Svmhw6 = (Ixmhw6 & Pxmhw6);
assign Pxmhw6 = (~(V1c7z6[28] & Gpmhw6));
assign Ixmhw6 = (Wxmhw6 & Dymhw6);
assign Dymhw6 = (~(Bqmhw6 & Zec7z6[0]));
assign K7i8v6 = (~(Kymhw6 & Rymhw6));
assign Rymhw6 = (Yymhw6 & Fzmhw6);
assign Fzmhw6 = (~(Bqmhw6 & Zec7z6[10]));
assign Yymhw6 = (Mzmhw6 & Xnmhw6);
assign Mzmhw6 = (~(Jnmhw6 & Ovbdt6));
assign Jnmhw6 = (Ammhw6 & Tzmhw6);
assign Tzmhw6 = (~(A0nhw6 & Uqehw6));
assign A0nhw6 = (H0nhw6 & O0nhw6);
assign H0nhw6 = (~(V0nhw6 & E3fhw6));
assign Kymhw6 = (C1nhw6 & J1nhw6);
assign J1nhw6 = (~(V1c7z6[27] & Gpmhw6));
assign C1nhw6 = (Q1nhw6 & X1nhw6);
assign X1nhw6 = (~(Eomhw6 & E2nhw6));
assign Q1nhw6 = (~(L2nhw6 & Uqd7z6[19]));
assign D7i8v6 = (~(S2nhw6 & Z2nhw6));
assign Z2nhw6 = (G3nhw6 & N3nhw6);
assign N3nhw6 = (~(Eomhw6 & U3nhw6));
assign G3nhw6 = (B4nhw6 & Xnmhw6);
assign B4nhw6 = (~(Bqmhw6 & Zec7z6[30]));
assign S2nhw6 = (I4nhw6 & P4nhw6);
assign P4nhw6 = (~(L2nhw6 & Uqd7z6[18]));
assign I4nhw6 = (~(V1c7z6[26] & Gpmhw6));
assign W6i8v6 = (~(W4nhw6 & D5nhw6));
assign D5nhw6 = (K5nhw6 & R5nhw6);
assign R5nhw6 = (~(Eomhw6 & Y5nhw6));
assign K5nhw6 = (F6nhw6 & Xnmhw6);
assign F6nhw6 = (~(Bqmhw6 & M6nhw6));
assign W4nhw6 = (T6nhw6 & A7nhw6);
assign A7nhw6 = (~(L2nhw6 & Uqd7z6[17]));
assign T6nhw6 = (~(V1c7z6[25] & Gpmhw6));
assign P6i8v6 = (~(H7nhw6 & O7nhw6));
assign O7nhw6 = (V7nhw6 & C8nhw6);
assign C8nhw6 = (~(Eomhw6 & J8nhw6));
assign V7nhw6 = (Q8nhw6 & Xnmhw6);
assign Xnmhw6 = (~(X8nhw6 & E9nhw6));
assign E9nhw6 = (~(L9nhw6 & S9nhw6));
assign Q8nhw6 = (~(Bqmhw6 & Z9nhw6));
assign H7nhw6 = (Ganhw6 & Nanhw6);
assign Nanhw6 = (~(L2nhw6 & Ovbdt6));
assign Ganhw6 = (~(V1c7z6[24] & Gpmhw6));
assign I6i8v6 = (~(Uanhw6 & Bbnhw6));
assign Bbnhw6 = (Ibnhw6 & Pbnhw6);
assign Pbnhw6 = (~(Wbnhw6 & Lomhw6));
assign Ibnhw6 = (Dcnhw6 & Kcnhw6);
assign Dcnhw6 = (~(Rcnhw6 & Ycnhw6));
assign Rcnhw6 = (M6nhw6 ^ Painv6);
assign Uanhw6 = (Fdnhw6 & Mdnhw6);
assign Mdnhw6 = (~(V1c7z6[23] & Gpmhw6));
assign Fdnhw6 = (Tdnhw6 & Aenhw6);
assign Aenhw6 = (~(Eomhw6 & Q1s8v6));
assign Tdnhw6 = (~(Henhw6 & Oenhw6));
assign B6i8v6 = (~(Venhw6 & Cfnhw6));
assign Cfnhw6 = (Jfnhw6 & Qfnhw6);
assign Qfnhw6 = (~(Ycnhw6 & Msnnv6));
assign Msnnv6 = (Zec7z6[10] ^ Offhw6);
assign Jfnhw6 = (Xfnhw6 & Kcnhw6);
assign Xfnhw6 = (~(Wbnhw6 & Rrmhw6));
assign Venhw6 = (Egnhw6 & Lgnhw6);
assign Lgnhw6 = (~(V1c7z6[22] & Gpmhw6));
assign Egnhw6 = (Sgnhw6 & Zgnhw6);
assign Zgnhw6 = (~(Eomhw6 & Ryr8v6));
assign Sgnhw6 = (~(Uqd7z6[22] & Henhw6));
assign U5i8v6 = (~(Ghnhw6 & Nhnhw6));
assign Nhnhw6 = (Uhnhw6 & Binhw6);
assign Binhw6 = (~(Ycnhw6 & Zec7z6[9]));
assign Uhnhw6 = (Iinhw6 & Kcnhw6);
assign Iinhw6 = (~(Wbnhw6 & Jumhw6));
assign Ghnhw6 = (Pinhw6 & Winhw6);
assign Winhw6 = (~(V1c7z6[21] & Gpmhw6));
assign Pinhw6 = (Djnhw6 & Kjnhw6);
assign Kjnhw6 = (~(Eomhw6 & Svr8v6));
assign Djnhw6 = (~(Uqd7z6[21] & Henhw6));
assign N5i8v6 = (~(Rjnhw6 & Yjnhw6));
assign Yjnhw6 = (Fknhw6 & Mknhw6);
assign Mknhw6 = (~(Ycnhw6 & Zec7z6[8]));
assign Fknhw6 = (Tknhw6 & Kcnhw6);
assign Kcnhw6 = (~(X8nhw6 & Alnhw6));
assign Alnhw6 = (~(Hlnhw6 & Olnhw6));
assign Hlnhw6 = (Pxnnv6 & H2sov6);
assign X8nhw6 = (Ammhw6 & Vlnhw6);
assign Vlnhw6 = (~(Olnhw6 & Painv6));
assign Tknhw6 = (~(Wbnhw6 & Bxmhw6));
assign Rjnhw6 = (Cmnhw6 & Jmnhw6);
assign Jmnhw6 = (~(V1c7z6[20] & Gpmhw6));
assign Cmnhw6 = (Qmnhw6 & Xmnhw6);
assign Xmnhw6 = (~(Eomhw6 & Tsr8v6));
assign Qmnhw6 = (~(Uqd7z6[20] & Henhw6));
assign G5i8v6 = (~(Ennhw6 & Lnnhw6));
assign Lnnhw6 = (Snnhw6 & Znnhw6);
assign Znnhw6 = (~(Ycnhw6 & Zec7z6[7]));
assign Snnhw6 = (Gonhw6 & Nonhw6);
assign Gonhw6 = (~(Eomhw6 & Uonhw6));
assign Ennhw6 = (~(Bpnhw6 | Ipnhw6));
assign Ipnhw6 = (Ammhw6 ? Ppnhw6 : V1c7z6[19]);
assign Ppnhw6 = (Wpnhw6 & Zec7z6[27]);
assign Bpnhw6 = (~(Dqnhw6 & Kqnhw6));
assign Kqnhw6 = (~(Uqd7z6[19] & Henhw6));
assign Dqnhw6 = (~(Wbnhw6 & E2nhw6));
assign Z4i8v6 = (~(Rqnhw6 & Yqnhw6));
assign Yqnhw6 = (Frnhw6 & Mrnhw6);
assign Mrnhw6 = (~(Ycnhw6 & Zec7z6[6]));
assign Ycnhw6 = (Ammhw6 & L4sov6);
assign Frnhw6 = (Trnhw6 & Nonhw6);
assign Trnhw6 = (~(Eomhw6 & Asnhw6));
assign Rqnhw6 = (~(Hsnhw6 | Osnhw6));
assign Osnhw6 = (Ammhw6 ? Vsnhw6 : V1c7z6[18]);
assign Vsnhw6 = (Wpnhw6 & M6nhw6);
assign Hsnhw6 = (~(Ctnhw6 & Jtnhw6));
assign Jtnhw6 = (~(Uqd7z6[18] & Henhw6));
assign Ctnhw6 = (~(Wbnhw6 & U3nhw6));
assign S4i8v6 = (~(Qtnhw6 & Xtnhw6));
assign Xtnhw6 = (Eunhw6 & Lunhw6);
assign Lunhw6 = (~(Uqd7z6[17] & Henhw6));
assign Eunhw6 = (Sunhw6 & Nonhw6);
assign Sunhw6 = (~(Eomhw6 & Zunhw6));
assign Eomhw6 = (Gvnhw6 & Ammhw6);
assign Gvnhw6 = (Nvnhw6 & Painv6);
assign Qtnhw6 = (~(Uvnhw6 | Bwnhw6));
assign Bwnhw6 = (Wbnhw6 & Y5nhw6);
assign Uvnhw6 = (Ammhw6 ? Iwnhw6 : V1c7z6[17]);
assign Iwnhw6 = (~(Zpehw6 | S9nhw6));
assign L4i8v6 = (~(Pwnhw6 & Wwnhw6));
assign Wwnhw6 = (Dxnhw6 & Nonhw6);
assign Dxnhw6 = (~(Ovbdt6 & Henhw6));
assign Henhw6 = (Bqmhw6 | Kxnhw6);
assign Kxnhw6 = (Rxnhw6 & Ammhw6);
assign Rxnhw6 = (~(Yxnhw6 | Kfa7z6));
assign Bqmhw6 = (Fynhw6 & Ammhw6);
assign Fynhw6 = (Mynhw6 & Zec7z6[7]);
assign Pwnhw6 = (~(Tynhw6 | Aznhw6));
assign Aznhw6 = (Wbnhw6 & J8nhw6);
assign Tynhw6 = (Ammhw6 ? Hznhw6 : V1c7z6[16]);
assign Hznhw6 = (~(Qtnov6 | S9nhw6));
assign E4i8v6 = (~(Oznhw6 & Vznhw6));
assign Vznhw6 = (C0ohw6 & Npmhw6);
assign Npmhw6 = (~(L2nhw6 & Oenhw6));
assign C0ohw6 = (J0ohw6 & Nonhw6);
assign J0ohw6 = (~(Q0ohw6 & Lomhw6));
assign Oznhw6 = (X0ohw6 & E1ohw6);
assign E1ohw6 = (Gpmhw6 ? S1ohw6 : L1ohw6);
assign X0ohw6 = (Z1ohw6 & G2ohw6);
assign G2ohw6 = (N2ohw6 | U2ohw6);
assign Z1ohw6 = (~(Wbnhw6 & Q1s8v6));
assign X3i8v6 = (~(B3ohw6 & I3ohw6));
assign I3ohw6 = (P3ohw6 & Msmhw6);
assign Msmhw6 = (~(L2nhw6 & Uqd7z6[22]));
assign P3ohw6 = (W3ohw6 & Nonhw6);
assign W3ohw6 = (~(Q0ohw6 & Rrmhw6));
assign Rrmhw6 = (D4ohw6 & K4ohw6);
assign B3ohw6 = (~(R4ohw6 | Y4ohw6));
assign Y4ohw6 = (Ammhw6 ? Dyfhw6 : V1c7z6[14]);
assign R4ohw6 = (~(F5ohw6 & M5ohw6));
assign M5ohw6 = (N2ohw6 | T5ohw6);
assign F5ohw6 = (~(Wbnhw6 & Ryr8v6));
assign Q3i8v6 = (~(A6ohw6 & H6ohw6));
assign H6ohw6 = (O6ohw6 & Evmhw6);
assign Evmhw6 = (~(L2nhw6 & Uqd7z6[21]));
assign O6ohw6 = (V6ohw6 & Nonhw6);
assign V6ohw6 = (~(Q0ohw6 & Jumhw6));
assign Jumhw6 = (C7ohw6 & Bat8v6);
assign Q0ohw6 = (Ammhw6 & J7ohw6);
assign A6ohw6 = (Q7ohw6 & X7ohw6);
assign X7ohw6 = (~(V1c7z6[13] & Gpmhw6));
assign Q7ohw6 = (E8ohw6 & L8ohw6);
assign L8ohw6 = (N2ohw6 | S8ohw6);
assign E8ohw6 = (~(Wbnhw6 & Svr8v6));
assign J3i8v6 = (~(Z8ohw6 & G9ohw6));
assign G9ohw6 = (N9ohw6 & U9ohw6);
assign U9ohw6 = (N2ohw6 | Baohw6);
assign N2ohw6 = (~(Ammhw6 & Iaohw6));
assign Iaohw6 = (~(S9nhw6 & Paohw6));
assign N9ohw6 = (Wxmhw6 & Nonhw6);
assign Nonhw6 = (~(Ammhw6 & Waohw6));
assign Waohw6 = (~(Olnhw6 & Pxnnv6));
assign Wxmhw6 = (~(L2nhw6 & Uqd7z6[20]));
assign L2nhw6 = (Ammhw6 & Dbohw6);
assign Z8ohw6 = (~(Kbohw6 | Rbohw6));
assign Rbohw6 = (Wbnhw6 & Tsr8v6);
assign Wbnhw6 = (Ammhw6 & Ybohw6);
assign Kbohw6 = (Ammhw6 ? Fcohw6 : V1c7z6[12]);
assign Fcohw6 = (~(Mcohw6 & Tcohw6));
assign Tcohw6 = (O0nhw6 | Adohw6);
assign Mcohw6 = (~(Hdohw6 | Ixfhw6));
assign Hdohw6 = (Bxmhw6 & J7ohw6);
assign Bxmhw6 = (~(M6nhw6 | Odohw6));
assign C3i8v6 = (!Vdohw6);
assign Vdohw6 = (Ammhw6 ? Lnghw6 : Ceohw6);
assign Lnghw6 = (Jeohw6 & Qeohw6);
assign Qeohw6 = (Xeohw6 & Efohw6);
assign Efohw6 = (L9nhw6 & Lfohw6);
assign Lfohw6 = (~(Ybohw6 & Uonhw6));
assign L9nhw6 = (Olnhw6 & Pxnnv6);
assign Pxnnv6 = (Sfohw6 | Painv6);
assign Xeohw6 = (Zfohw6 & Ggohw6);
assign Ggohw6 = (~(Zec7z6[27] & Ngohw6));
assign Zfohw6 = (~(J7ohw6 & E2nhw6));
assign E2nhw6 = (!Ugohw6);
assign Ugohw6 = (Oenhw6 ? Ihohw6 : Bhohw6);
assign Ihohw6 = (Phohw6 & Whohw6);
assign Whohw6 = (~(Diohw6 & Uqd7z6[22]));
assign Phohw6 = (~(D4ohw6 & Uqd7z6[20]));
assign Bhohw6 = (Kiohw6 & Riohw6);
assign Riohw6 = (~(Diohw6 & Uqd7z6[21]));
assign Kiohw6 = (~(Yiohw6 & Kfa7z6));
assign Yiohw6 = (~(Bat8v6 & Fjohw6));
assign Jeohw6 = (Mjohw6 & Tjohw6);
assign Tjohw6 = (Akohw6 & Hkohw6);
assign Hkohw6 = (~(Dbohw6 & Uqd7z6[19]));
assign Akohw6 = (~(Zec7z6[10] & Okohw6));
assign Mjohw6 = (Vkohw6 & Clohw6);
assign Clohw6 = (O0nhw6 | Bat8v6);
assign Vkohw6 = (Jlohw6 | S9nhw6);
assign V2i8v6 = (!Qlohw6);
assign Qlohw6 = (Ammhw6 ? Ppghw6 : Xlohw6);
assign Ppghw6 = (Emohw6 & Lmohw6);
assign Lmohw6 = (Smohw6 & Zmohw6);
assign Zmohw6 = (Gnohw6 & Nnohw6);
assign Nnohw6 = (~(Zec7z6[26] & Ngohw6));
assign Gnohw6 = (Unohw6 & Olnhw6);
assign Unohw6 = (~(Asnhw6 & Ybohw6));
assign Smohw6 = (Boohw6 & Ioohw6);
assign Ioohw6 = (~(J7ohw6 & U3nhw6));
assign U3nhw6 = (Poohw6 | Woohw6);
assign Woohw6 = (Oenhw6 ? Kpohw6 : Dpohw6);
assign Kpohw6 = (Uqd7z6[19] & Kfa7z6);
assign Poohw6 = (~(Rpohw6 & Ypohw6));
assign Ypohw6 = (~(Diohw6 & Fqohw6));
assign Rpohw6 = (~(Mqohw6 & K4ohw6));
assign Boohw6 = (~(Dbohw6 & Uqd7z6[18]));
assign Emohw6 = (Tqohw6 & Arohw6);
assign Arohw6 = (Hrohw6 & Orohw6);
assign Orohw6 = (~(Zec7z6[30] & Okohw6));
assign Hrohw6 = (O0nhw6 | Kfa7z6);
assign Tqohw6 = (Dynnv6 & Vrohw6);
assign Vrohw6 = (Buihw6 | S9nhw6);
assign Dynnv6 = (~(Csohw6 & Zec7z6[9]));
assign O2i8v6 = (!Jsohw6);
assign Jsohw6 = (Ammhw6 ? Trghw6 : Qsohw6);
assign Trghw6 = (Xsohw6 & Etohw6);
assign Etohw6 = (Ltohw6 & Stohw6);
assign Stohw6 = (Ztohw6 & Guohw6);
assign Guohw6 = (~(Nuohw6 & Oenhw6));
assign Ztohw6 = (Uuohw6 & Olnhw6);
assign Olnhw6 = (T1sov6 | Xeinv6);
assign Uuohw6 = (Xeinv6 | Bvohw6);
assign Ltohw6 = (Ivohw6 & Pvohw6);
assign Pvohw6 = (~(Zec7z6[25] & Ngohw6));
assign Ivohw6 = (~(Zunhw6 & Ybohw6));
assign Ybohw6 = (Nvnhw6 & Adohw6);
assign Xsohw6 = (Wvohw6 & Dwohw6);
assign Dwohw6 = (Kwohw6 & Rwohw6);
assign Rwohw6 = (~(Okohw6 & M6nhw6));
assign Kwohw6 = (Ywohw6 & Fxohw6);
assign Fxohw6 = (~(J7ohw6 & Y5nhw6));
assign Y5nhw6 = (~(Mxohw6 & Txohw6));
assign Txohw6 = (~(C7ohw6 & M6nhw6));
assign C7ohw6 = (Oenhw6 ? Hyohw6 : Ayohw6);
assign Hyohw6 = (Uqd7z6[22] & Kfa7z6);
assign Ayohw6 = (~(Kfa7z6 & Dsehw6));
assign Mxohw6 = (Sfa7z6 ? Vyohw6 : Oyohw6);
assign Oyohw6 = (!Dpohw6);
assign Dpohw6 = (~(Czohw6 & Jzohw6));
assign Jzohw6 = (~(Diohw6 & Uqd7z6[20]));
assign Czohw6 = (~(D4ohw6 & Uqd7z6[18]));
assign Ywohw6 = (~(Dbohw6 & Uqd7z6[17]));
assign Wvohw6 = (Mlnnv6 & Qzohw6);
assign Qzohw6 = (Lofhw6 | S9nhw6);
assign Mlnnv6 = (~(Csohw6 & Zec7z6[8]));
assign H2i8v6 = (!Xzohw6);
assign Xzohw6 = (Ammhw6 ? Xtghw6 : E0phw6);
assign Xtghw6 = (L0phw6 & S0phw6);
assign S0phw6 = (Z0phw6 & G1phw6);
assign G1phw6 = (N1phw6 & U1phw6);
assign U1phw6 = (~(Uqd7z6[22] & Nuohw6));
assign Nuohw6 = (~(B2phw6 & O0nhw6));
assign N1phw6 = (~(Zec7z6[24] & Ngohw6));
assign Ngohw6 = (Zofhw6 | I2phw6);
assign Z0phw6 = (P2phw6 & W2phw6);
assign W2phw6 = (~(J7ohw6 & J8nhw6));
assign J8nhw6 = (~(D3phw6 & K3phw6));
assign K3phw6 = (Oenhw6 ? Vyohw6 : R3phw6);
assign Vyohw6 = (Y3phw6 & F4phw6);
assign F4phw6 = (~(Diohw6 & Uqd7z6[19]));
assign Y3phw6 = (~(D4ohw6 & Uqd7z6[17]));
assign R3phw6 = (~(Diohw6 & Uqd7z6[18]));
assign Diohw6 = (~(M6nhw6 | Kfa7z6));
assign D3phw6 = (M4phw6 & T4phw6);
assign T4phw6 = (~(Lomhw6 & Ovbdt6));
assign Lomhw6 = (D4ohw6 & Sfa7z6);
assign M4phw6 = (Odohw6 | Bat8v6);
assign Odohw6 = (~(A5phw6 | Fqohw6));
assign A5phw6 = (Z9nhw6 ? K4ohw6 : H5phw6);
assign H5phw6 = (Uqd7z6[20] & Sfa7z6);
assign P2phw6 = (~(Dbohw6 & Ovbdt6));
assign Dbohw6 = (~(Yxnhw6 | Bat8v6));
assign L0phw6 = (O5phw6 & V5phw6);
assign V5phw6 = (C6phw6 & J6phw6);
assign J6phw6 = (~(Okohw6 & Z9nhw6));
assign C6phw6 = (~(Zec7z6[6] & Zwlhw6));
assign O5phw6 = (Q6phw6 & X6phw6);
assign X6phw6 = (S9nhw6 | Sfa7z6);
assign Q6phw6 = (Xeinv6 | E7phw6);
assign A2i8v6 = (Gpmhw6 ? V1c7z6[7] : Dxghw6);
assign T1i8v6 = (Gpmhw6 ? V1c7z6[6] : C0hhw6);
assign M1i8v6 = (!L7phw6);
assign L7phw6 = (Ammhw6 ? Y4hhw6 : S7phw6);
assign F1i8v6 = (Gpmhw6 ? V1c7z6[4] : Wahhw6);
assign Y0i8v6 = (!Z7phw6);
assign Z7phw6 = (Ammhw6 ? Vdhhw6 : G8phw6);
assign R0i8v6 = (Gpmhw6 ? V1c7z6[2] : Kphhw6);
assign K0i8v6 = (Gpmhw6 ? V1c7z6[1] : Ywhhw6);
assign Gpmhw6 = (!Ammhw6);
assign Ammhw6 = (~(Z2onv6 | N8phw6));
assign N8phw6 = (U8phw6 & B9phw6);
assign B9phw6 = (I9phw6 & P9phw6);
assign P9phw6 = (W9phw6 & Kkmhw6);
assign I9phw6 = (Daphw6 & Kaphw6);
assign U8phw6 = (Raphw6 & Yaphw6);
assign Yaphw6 = (~(Fbphw6 | Mbphw6));
assign Raphw6 = (Tbphw6 & Xvehw6);
assign D0i8v6 = (Hcphw6 ? Wfxdt6 : Acphw6);
assign Hcphw6 = (Nnaov6 & Ocphw6);
assign Ocphw6 = (~(Vcphw6 & Cdphw6));
assign Cdphw6 = (Jdphw6 & Qdphw6);
assign Qdphw6 = (~(Cehhw6 | Xdphw6));
assign Jdphw6 = (Cwlnv6 & Gr2et6);
assign Vcphw6 = (~(Eephw6 | A6hhw6));
assign Eephw6 = (Rphhw6 | Rbhhw6);
assign Nnaov6 = (!W4nov6);
assign W4nov6 = (~(Lephw6 & Sephw6));
assign Sephw6 = (Zephw6 & Gfphw6);
assign Gfphw6 = (Nfphw6 & Ufphw6);
assign Nfphw6 = (~(Clhhw6 & Jc2et6));
assign Jc2et6 = (~(Vrinv6 & Kwinv6));
assign Kwinv6 = (Ypinv6 | Bfo7v6);
assign Zephw6 = (Bgphw6 & Igphw6);
assign Igphw6 = (~(Gr2et6 & Pgphw6));
assign Pgphw6 = (~(Wgphw6 & Dhphw6));
assign Dhphw6 = (Khphw6 & Rhphw6);
assign Khphw6 = (Jsaov6 & Srknv6);
assign Wgphw6 = (Yhphw6 & Jzaov6);
assign Jzaov6 = (Fiphw6 & Miphw6);
assign Miphw6 = (~(Tiphw6 & Fxaov6));
assign Fiphw6 = (Ajphw6 & Hjphw6);
assign Yhphw6 = (Ojphw6 & Vjphw6);
assign Vjphw6 = (~(Ckphw6 & Vqihw6));
assign Bgphw6 = (~(Jkphw6 & O5a7z6));
assign Jkphw6 = (Qkphw6 & Xkphw6);
assign Xkphw6 = (~(Txaov6 & Elphw6));
assign Qkphw6 = (~(Xdphw6 & Qtvnv6));
assign Lephw6 = (Llphw6 & Slphw6);
assign Slphw6 = (~(Zlphw6 & Gmphw6));
assign Zlphw6 = (Nmphw6 & Qtvnv6);
assign Nmphw6 = (~(Umphw6 & Bnphw6));
assign Bnphw6 = (Inphw6 | Iga7z6);
assign Umphw6 = (Txaov6 | Uebdt6);
assign Txaov6 = (Pnphw6 & Wnphw6);
assign Wnphw6 = (~(Dophw6 & Fulnv6));
assign Pnphw6 = (~(Kophw6 & Dioov6));
assign Llphw6 = (Rophw6 & Yophw6);
assign Yophw6 = (~(Lyknv6 & C0ydt6));
assign Rophw6 = (~(Fpphw6 & Msmov6));
assign Acphw6 = (~(Mpphw6 & Tpphw6));
assign Tpphw6 = (~(Aqphw6 & Hqphw6));
assign Hqphw6 = (Oqphw6 & Vqphw6);
assign Vqphw6 = (~(Crphw6 | Cehhw6));
assign Crphw6 = (Mqhhw6 | S1wnv6);
assign Oqphw6 = (Jrphw6 & Ldo7v6);
assign Jrphw6 = (Pbadt6 & Rphhw6);
assign Aqphw6 = (Qrphw6 & Xrphw6);
assign Xrphw6 = (Esphw6 & Ecc7z6[5]);
assign Esphw6 = (Tlmov6 & Lsphw6);
assign Qrphw6 = (~(Rbhhw6 | A6hhw6));
assign Mpphw6 = (~(Ssphw6 & Cwlnv6));
assign Ssphw6 = (Msmov6 & Yioov6);
assign Wzh8v6 = (!Zsphw6);
assign Zsphw6 = (Vfmov6 ? Hjihw6 : Sj77z6);
assign Pzh8v6 = (Gtphw6 ? Q1h7z6[0] : Rphhw6);
assign Izh8v6 = (Gtphw6 ? Q1h7z6[1] : Cehhw6);
assign Bzh8v6 = (Gtphw6 ? Q1h7z6[2] : Rbhhw6);
assign Uyh8v6 = (Gtphw6 ? Q1h7z6[3] : A6hhw6);
assign Nyh8v6 = (Q1h7z6[4] & Gtphw6);
assign Gyh8v6 = (Q1h7z6[5] & Gtphw6);
assign Gtphw6 = (!Iwvnv6);
assign Zxh8v6 = (Utphw6 ? Gg7et6 : Ntphw6);
assign Utphw6 = (Buphw6 & Iuphw6);
assign Iuphw6 = (~(Wmknv6 & Gr2et6));
assign Wmknv6 = (Gg7et6 & Puphw6);
assign Buphw6 = (~(Wuphw6 & Dvphw6));
assign Dvphw6 = (Kvphw6 & Vxihw6);
assign Kvphw6 = (Rvphw6 & Ntphw6);
assign Rvphw6 = (~(Yvphw6 & Fwphw6));
assign Yvphw6 = (~(Etinv6 & Iga7z6));
assign Wuphw6 = (Ecc7z6[11] & Mwphw6);
assign Ntphw6 = (~(Twphw6 & Fwphw6));
assign Fwphw6 = (~(Axphw6 & Hxphw6));
assign Hxphw6 = (Oxphw6 & Vxphw6);
assign Oxphw6 = (Bfo7v6 & Hjihw6);
assign Axphw6 = (O5a7z6 & Tnzdt6);
assign Sxh8v6 = (Uimov6 ? Ozadt6 : Cyphw6);
assign Lxh8v6 = (~(Jyphw6 & Qyphw6));
assign Qyphw6 = (~(Xyphw6 & Ezphw6));
assign Xyphw6 = (Lzphw6 & Szphw6);
assign Jyphw6 = (~(Dkm7z6[1] & Zzphw6));
assign Exh8v6 = (N0qhw6 ? S7n7z6[0] : G0qhw6);
assign G0qhw6 = (~(U0qhw6 & B1qhw6));
assign B1qhw6 = (~(Wbhnv6 & Fbqnv6));
assign U0qhw6 = (~(Uclov6 & Hub7z6[0]));
assign Xwh8v6 = (N0qhw6 ? S7n7z6[1] : I1qhw6);
assign I1qhw6 = (~(P1qhw6 & W1qhw6));
assign W1qhw6 = (~(Fbqnv6 & Anehw6));
assign P1qhw6 = (~(Uclov6 & Hub7z6[1]));
assign Qwh8v6 = (~(D2qhw6 & K2qhw6));
assign K2qhw6 = (~(R2qhw6 & Cyphw6));
assign D2qhw6 = (~(E1uet6 & Y2qhw6));
assign Jwh8v6 = (~(F3qhw6 & M3qhw6));
assign M3qhw6 = (~(T3qhw6 & A4qhw6));
assign F3qhw6 = (~(H4qhw6 & Znn7z6[1]));
assign Cwh8v6 = (V4qhw6 ? O4qhw6 : Ppzet6);
assign V4qhw6 = (Kr97z6 & C5qhw6);
assign C5qhw6 = (~(O4qhw6 & J5qhw6));
assign J5qhw6 = (~(Q5qhw6 & X5qhw6));
assign X5qhw6 = (~(E6qhw6 | L6qhw6));
assign Q5qhw6 = (Ee47v6 & Dbymz6[1]);
assign Vvh8v6 = (Z6qhw6 ? S6qhw6 : Io47v6);
assign S6qhw6 = (!Cewnv6);
assign Ovh8v6 = (~(G7qhw6 & N7qhw6));
assign N7qhw6 = (~(S067v6 & U7qhw6));
assign U7qhw6 = (~(L5ymz6[8] & B8qhw6));
assign G7qhw6 = (W8qhw6 ? P8qhw6 : I8qhw6);
assign I8qhw6 = (~(D9qhw6 & K9qhw6));
assign D9qhw6 = (~(R9qhw6 | Y9qhw6));
assign Y9qhw6 = (Kh47v6 & Gj47v6);
assign Hvh8v6 = (~(Faqhw6 & Maqhw6));
assign Maqhw6 = (Taqhw6 & Abqhw6);
assign Abqhw6 = (~(Krxmz6[31] & Hbqhw6));
assign Taqhw6 = (~(Obqhw6 & Ii47v6));
assign Faqhw6 = (Vbqhw6 & Ccqhw6);
assign Ccqhw6 = (~(Jcqhw6 & Coxmz6[31]));
assign Vbqhw6 = (Edqhw6 ? Xcqhw6 : Qcqhw6);
assign Xcqhw6 = (!Cxxmz6[31]);
assign Qcqhw6 = (Ldqhw6 | Sdqhw6);
assign Avh8v6 = (Zdqhw6 ? Omxmz6[31] : Cxxmz6[31]);
assign Tuh8v6 = (~(Geqhw6 & Neqhw6));
assign Neqhw6 = (~(Dbymz6[0] & Ueqhw6));
assign Ueqhw6 = (~(Adwnv6 & Bfqhw6));
assign Bfqhw6 = (~(Ifqhw6 & Qewnv6));
assign Ifqhw6 = (Jewnv6 & Cewnv6);
assign Cewnv6 = (~(Pfqhw6 & Wfqhw6));
assign Wfqhw6 = (Dgqhw6 & Kgqhw6);
assign Dgqhw6 = (Rgqhw6 & Ygqhw6);
assign Pfqhw6 = (Oeo7z6[0] & Fhqhw6);
assign Fhqhw6 = (~(Mhqhw6 & Thqhw6));
assign Thqhw6 = (~(Fvzet6 | Tszet6));
assign Mhqhw6 = (Gco7z6[6] & Aiqhw6);
assign Jewnv6 = (Viqhw6 ? Oiqhw6 : Hiqhw6);
assign Oiqhw6 = (~(Cjqhw6 & Jjqhw6));
assign Hiqhw6 = (~(Qjqhw6 & Xjqhw6));
assign Geqhw6 = (~(Adwnv6 & Ekqhw6));
assign Adwnv6 = (Kr97z6 & Lkqhw6);
assign Lkqhw6 = (~(Skqhw6 & Zkqhw6));
assign Zkqhw6 = (~(Dbymz6[0] & Glqhw6));
assign Skqhw6 = (~(Ekqhw6 ^ Nlqhw6));
assign Nlqhw6 = (~(Dbymz6[0] | Ye47v6));
assign Muh8v6 = (Bmqhw6 ? F5o7z6[2] : Ulqhw6);
assign Fuh8v6 = (Bmqhw6 ? F5o7z6[3] : Imqhw6);
assign Yth8v6 = (Bmqhw6 ? F5o7z6[4] : Pmqhw6);
assign Rth8v6 = (Bmqhw6 ? F5o7z6[5] : Wmqhw6);
assign Kth8v6 = (Bmqhw6 ? F5o7z6[6] : Dnqhw6);
assign Dth8v6 = (Bmqhw6 ? F5o7z6[7] : Knqhw6);
assign Wsh8v6 = (Rnqhw6 ? Cb77z6 : Gco7z6[6]);
assign Psh8v6 = (~(Ynqhw6 & Foqhw6));
assign Foqhw6 = (Moqhw6 & Toqhw6);
assign Toqhw6 = (~(Tfxmz6[1] & Zfwnv6));
assign Moqhw6 = (~(Njxmz6[1] & Ggwnv6));
assign Ynqhw6 = (Apqhw6 & Hpqhw6);
assign Hpqhw6 = (~(Ul67v6 & Bhwnv6));
assign Apqhw6 = (~(Hnxmz6[1] & Ihwnv6));
assign Ish8v6 = (~(Opqhw6 & Vpqhw6));
assign Vpqhw6 = (Cqqhw6 & Jqqhw6);
assign Jqqhw6 = (~(Tfxmz6[2] & Zfwnv6));
assign Cqqhw6 = (~(Njxmz6[2] & Ggwnv6));
assign Opqhw6 = (Qqqhw6 & Xqqhw6);
assign Xqqhw6 = (~(Uk67v6 & Bhwnv6));
assign Qqqhw6 = (~(Hnxmz6[2] & Ihwnv6));
assign Bsh8v6 = (~(Erqhw6 & Lrqhw6));
assign Lrqhw6 = (Srqhw6 & Zrqhw6);
assign Zrqhw6 = (~(Tfxmz6[3] & Zfwnv6));
assign Srqhw6 = (~(Njxmz6[3] & Ggwnv6));
assign Erqhw6 = (Gsqhw6 & Nsqhw6);
assign Nsqhw6 = (~(Uj67v6 & Bhwnv6));
assign Gsqhw6 = (~(Hnxmz6[3] & Ihwnv6));
assign Urh8v6 = (~(Usqhw6 & Btqhw6));
assign Btqhw6 = (Itqhw6 & Ptqhw6);
assign Ptqhw6 = (~(Tfxmz6[4] & Zfwnv6));
assign Itqhw6 = (~(Njxmz6[4] & Ggwnv6));
assign Usqhw6 = (Wtqhw6 & Duqhw6);
assign Duqhw6 = (~(Ui67v6 & Bhwnv6));
assign Wtqhw6 = (~(Hnxmz6[4] & Ihwnv6));
assign Nrh8v6 = (~(Kuqhw6 & Ruqhw6));
assign Ruqhw6 = (Yuqhw6 & Fvqhw6);
assign Fvqhw6 = (~(Tfxmz6[5] & Zfwnv6));
assign Yuqhw6 = (~(Njxmz6[5] & Ggwnv6));
assign Kuqhw6 = (Mvqhw6 & Tvqhw6);
assign Tvqhw6 = (~(Uh67v6 & Bhwnv6));
assign Mvqhw6 = (~(Hnxmz6[5] & Ihwnv6));
assign Grh8v6 = (~(Awqhw6 & Hwqhw6));
assign Hwqhw6 = (Owqhw6 & Vwqhw6);
assign Vwqhw6 = (~(Tfxmz6[6] & Zfwnv6));
assign Owqhw6 = (~(Njxmz6[6] & Ggwnv6));
assign Awqhw6 = (Cxqhw6 & Jxqhw6);
assign Jxqhw6 = (~(Ug67v6 & Bhwnv6));
assign Cxqhw6 = (~(Hnxmz6[6] & Ihwnv6));
assign Zqh8v6 = (~(Qxqhw6 & Xxqhw6));
assign Xxqhw6 = (Eyqhw6 & Lyqhw6);
assign Lyqhw6 = (~(Tfxmz6[7] & Zfwnv6));
assign Eyqhw6 = (~(Njxmz6[7] & Ggwnv6));
assign Qxqhw6 = (Syqhw6 & Zyqhw6);
assign Zyqhw6 = (~(Uf67v6 & Bhwnv6));
assign Syqhw6 = (~(Hnxmz6[7] & Ihwnv6));
assign Sqh8v6 = (~(Gzqhw6 & Nzqhw6));
assign Nzqhw6 = (Uzqhw6 & B0rhw6);
assign B0rhw6 = (~(Tfxmz6[8] & Zfwnv6));
assign Uzqhw6 = (~(Njxmz6[8] & Ggwnv6));
assign Gzqhw6 = (I0rhw6 & P0rhw6);
assign P0rhw6 = (~(Ue67v6 & Bhwnv6));
assign I0rhw6 = (~(Hnxmz6[8] & Ihwnv6));
assign Lqh8v6 = (~(W0rhw6 & D1rhw6));
assign D1rhw6 = (K1rhw6 & R1rhw6);
assign R1rhw6 = (~(Tfxmz6[9] & Zfwnv6));
assign K1rhw6 = (~(Njxmz6[9] & Ggwnv6));
assign W0rhw6 = (Y1rhw6 & F2rhw6);
assign F2rhw6 = (~(Ud67v6 & Bhwnv6));
assign Y1rhw6 = (~(Hnxmz6[9] & Ihwnv6));
assign Eqh8v6 = (~(M2rhw6 & T2rhw6));
assign T2rhw6 = (A3rhw6 & H3rhw6);
assign H3rhw6 = (~(Tfxmz6[10] & Zfwnv6));
assign A3rhw6 = (~(Njxmz6[10] & Ggwnv6));
assign M2rhw6 = (O3rhw6 & V3rhw6);
assign V3rhw6 = (~(Uc67v6 & Bhwnv6));
assign O3rhw6 = (~(Hnxmz6[10] & Ihwnv6));
assign Xph8v6 = (~(C4rhw6 & J4rhw6));
assign J4rhw6 = (Q4rhw6 & X4rhw6);
assign X4rhw6 = (~(Tfxmz6[0] & Zfwnv6));
assign Zfwnv6 = (E5rhw6 & JTAGNSW);
assign E5rhw6 = (L5rhw6 & E6qhw6);
assign Q4rhw6 = (~(Njxmz6[0] & Ggwnv6));
assign Ggwnv6 = (S5rhw6 & L5rhw6);
assign S5rhw6 = (Dz1nv6 & E6qhw6);
assign C4rhw6 = (Z5rhw6 & G6rhw6);
assign G6rhw6 = (~(Um67v6 & Bhwnv6));
assign Bhwnv6 = (N6rhw6 & U6rhw6);
assign N6rhw6 = (Dbymz6[0] & L5rhw6);
assign Z5rhw6 = (~(Hnxmz6[0] & Ihwnv6));
assign Ihwnv6 = (!L5rhw6);
assign L5rhw6 = (~(B7rhw6 & I7rhw6));
assign I7rhw6 = (~(Z6qhw6 & P7rhw6));
assign P7rhw6 = (U6rhw6 | Ee47v6);
assign U6rhw6 = (Qewnv6 & W7rhw6);
assign W7rhw6 = (~(D8rhw6 & K8rhw6));
assign K8rhw6 = (~(Qjqhw6 & Cjqhw6));
assign D8rhw6 = (Viqhw6 ? Cjqhw6 : Qjqhw6);
assign Cjqhw6 = (!Xjqhw6);
assign Qewnv6 = (~(R8rhw6 | Ee47v6));
assign R8rhw6 = (Y8rhw6 & F9rhw6);
assign F9rhw6 = (M9rhw6 & T9rhw6);
assign T9rhw6 = (~(Aarhw6 | Hnxmz6[7]));
assign Aarhw6 = (Hnxmz6[8] | Hnxmz6[9]);
assign M9rhw6 = (~(Harhw6 | Hnxmz6[4]));
assign Harhw6 = (Hnxmz6[5] | Hnxmz6[6]);
assign Y8rhw6 = (Oarhw6 & Varhw6);
assign Varhw6 = (~(Cbrhw6 | Hnxmz6[1]));
assign Cbrhw6 = (Hnxmz6[2] | Hnxmz6[3]);
assign Oarhw6 = (~(Jbrhw6 | Hnxmz6[0]));
assign Jbrhw6 = (Hnxmz6[10] | Hnxmz6[11]);
assign B7rhw6 = (~(Qbrhw6 & Xbrhw6));
assign Xbrhw6 = (E6qhw6 & Ekqhw6);
assign Qbrhw6 = (Ye47v6 & Kr97z6);
assign Qph8v6 = (~(Ecrhw6 & Lcrhw6));
assign Lcrhw6 = (~(Cxxmz6[23] & Scrhw6));
assign Ecrhw6 = (Zcrhw6 & Gdrhw6);
assign Gdrhw6 = (~(Ndrhw6 & Njxmz6[11]));
assign Zcrhw6 = (~(Udrhw6 & Hnxmz6[11]));
assign Jph8v6 = (Berhw6 & Ierhw6);
assign Ierhw6 = (Perhw6 & Werhw6);
assign Berhw6 = (Dfrhw6 & Lc57v6);
assign Cph8v6 = (~(Kfrhw6 & Rfrhw6));
assign Rfrhw6 = (~(R957v6 & Yfrhw6));
assign Voh8v6 = (~(Fgrhw6 & Mgrhw6));
assign Mgrhw6 = (~(Tgrhw6 & Io47v6));
assign Fgrhw6 = (Ahrhw6 & Hhrhw6);
assign Ahrhw6 = (~(H557v6 & Ohrhw6));
assign Ooh8v6 = (~(Vhrhw6 & Cirhw6));
assign Cirhw6 = (Jirhw6 & Qirhw6);
assign Qirhw6 = (Xirhw6 & Ejrhw6);
assign Xirhw6 = (~(Ovxmz6[1] & Ljrhw6));
assign Jirhw6 = (Sjrhw6 & Zjrhw6);
assign Zjrhw6 = (~(Coxmz6[1] & Gkrhw6));
assign Sjrhw6 = (~(Nkrhw6 & Cxxmz6[2]));
assign Vhrhw6 = (Ukrhw6 & Blrhw6);
assign Blrhw6 = (~(Cxxmz6[1] & Edqhw6));
assign Ukrhw6 = (Ilrhw6 & Plrhw6);
assign Plrhw6 = (~(Krxmz6[1] & Hbqhw6));
assign Ilrhw6 = (~(V357v6 & Obqhw6));
assign Hoh8v6 = (~(Wlrhw6 & Dmrhw6));
assign Dmrhw6 = (Kmrhw6 & Rmrhw6);
assign Rmrhw6 = (~(Krxmz6[2] & Hbqhw6));
assign Kmrhw6 = (Ymrhw6 & Ejrhw6);
assign Ymrhw6 = (~(Cxxmz6[3] & Nkrhw6));
assign Wlrhw6 = (Fnrhw6 & Mnrhw6);
assign Mnrhw6 = (~(Coxmz6[2] & Jcqhw6));
assign Fnrhw6 = (Tnrhw6 & Aorhw6);
assign Aorhw6 = (~(Blxmz6[0] & Obqhw6));
assign Tnrhw6 = (~(Cxxmz6[2] & Edqhw6));
assign Aoh8v6 = (~(Horhw6 & Oorhw6));
assign Oorhw6 = (Vorhw6 & Cprhw6);
assign Cprhw6 = (~(Blxmz6[1] & Obqhw6));
assign Vorhw6 = (Jprhw6 & Qprhw6);
assign Qprhw6 = (~(Cxxmz6[4] & Nkrhw6));
assign Jprhw6 = (~(Krxmz6[3] & Hbqhw6));
assign Horhw6 = (Xprhw6 & Eqrhw6);
assign Eqrhw6 = (~(Cxxmz6[3] & Edqhw6));
assign Xprhw6 = (~(Coxmz6[3] & Jcqhw6));
assign Tnh8v6 = (~(Lqrhw6 & Sqrhw6));
assign Sqrhw6 = (Zqrhw6 & Grrhw6);
assign Grrhw6 = (~(Krxmz6[4] & Hbqhw6));
assign Zqrhw6 = (Nrrhw6 & Ejrhw6);
assign Nrrhw6 = (~(Cxxmz6[5] & Nkrhw6));
assign Lqrhw6 = (Urrhw6 & Bsrhw6);
assign Bsrhw6 = (~(Coxmz6[4] & Jcqhw6));
assign Urrhw6 = (Isrhw6 & Psrhw6);
assign Psrhw6 = (~(S657v6 & Obqhw6));
assign Isrhw6 = (~(Cxxmz6[4] & Edqhw6));
assign Mnh8v6 = (~(Wsrhw6 & Dtrhw6));
assign Dtrhw6 = (Ktrhw6 & Rtrhw6);
assign Rtrhw6 = (~(Krxmz6[5] & Hbqhw6));
assign Ktrhw6 = (Ytrhw6 & Ejrhw6);
assign Ytrhw6 = (~(Cxxmz6[6] & Nkrhw6));
assign Wsrhw6 = (Furhw6 & Murhw6);
assign Murhw6 = (~(Coxmz6[5] & Jcqhw6));
assign Furhw6 = (Turhw6 & Avrhw6);
assign Avrhw6 = (~(H557v6 & Obqhw6));
assign Turhw6 = (~(Cxxmz6[5] & Edqhw6));
assign Fnh8v6 = (~(Hvrhw6 & Ovrhw6));
assign Ovrhw6 = (Vvrhw6 & Cwrhw6);
assign Cwrhw6 = (Ejrhw6 & Jwrhw6);
assign Jwrhw6 = (!Ljrhw6);
assign Vvrhw6 = (Qwrhw6 & Xwrhw6);
assign Xwrhw6 = (~(Yt47v6 & Exrhw6));
assign Qwrhw6 = (~(Coxmz6[6] & Gkrhw6));
assign Hvrhw6 = (Lxrhw6 & Sxrhw6);
assign Sxrhw6 = (~(Cxxmz6[6] & Edqhw6));
assign Lxrhw6 = (Zxrhw6 & Gyrhw6);
assign Gyrhw6 = (~(Cxxmz6[7] & Nkrhw6));
assign Zxrhw6 = (~(Krxmz6[6] & Hbqhw6));
assign Ymh8v6 = (~(Nyrhw6 & Uyrhw6));
assign Uyrhw6 = (Bzrhw6 & Izrhw6);
assign Izrhw6 = (~(Ud57v6 & Obqhw6));
assign Bzrhw6 = (Pzrhw6 & Wzrhw6);
assign Wzrhw6 = (~(Cxxmz6[8] & Nkrhw6));
assign Pzrhw6 = (~(Krxmz6[7] & Hbqhw6));
assign Nyrhw6 = (D0shw6 & K0shw6);
assign K0shw6 = (~(Cxxmz6[7] & Edqhw6));
assign D0shw6 = (~(Coxmz6[7] & Jcqhw6));
assign Rmh8v6 = (~(R0shw6 & Y0shw6));
assign Y0shw6 = (F1shw6 & M1shw6);
assign M1shw6 = (~(Krxmz6[8] & Hbqhw6));
assign F1shw6 = (T1shw6 & A2shw6);
assign A2shw6 = (~(Fuxmz6[0] & Ljrhw6));
assign T1shw6 = (~(Cxxmz6[9] & Nkrhw6));
assign R0shw6 = (H2shw6 & O2shw6);
assign O2shw6 = (~(Coxmz6[8] & Jcqhw6));
assign H2shw6 = (V2shw6 & C3shw6);
assign C3shw6 = (~(Ikxmz6[0] & Obqhw6));
assign V2shw6 = (~(Cxxmz6[8] & Edqhw6));
assign Kmh8v6 = (~(J3shw6 & Q3shw6));
assign Q3shw6 = (X3shw6 & E4shw6);
assign E4shw6 = (~(Krxmz6[9] & Hbqhw6));
assign X3shw6 = (L4shw6 & S4shw6);
assign S4shw6 = (~(Fuxmz6[1] & Ljrhw6));
assign L4shw6 = (~(Cxxmz6[10] & Nkrhw6));
assign J3shw6 = (Z4shw6 & G5shw6);
assign G5shw6 = (~(Coxmz6[9] & Jcqhw6));
assign Z4shw6 = (N5shw6 & U5shw6);
assign U5shw6 = (~(Ikxmz6[1] & Obqhw6));
assign N5shw6 = (~(Cxxmz6[9] & Edqhw6));
assign Dmh8v6 = (~(B6shw6 & I6shw6));
assign I6shw6 = (P6shw6 & W6shw6);
assign W6shw6 = (~(Krxmz6[10] & Hbqhw6));
assign P6shw6 = (D7shw6 & Ejrhw6);
assign D7shw6 = (~(Cxxmz6[11] & Nkrhw6));
assign B6shw6 = (K7shw6 & R7shw6);
assign R7shw6 = (~(Coxmz6[10] & Jcqhw6));
assign K7shw6 = (Y7shw6 & F8shw6);
assign F8shw6 = (~(Ikxmz6[2] & Obqhw6));
assign Y7shw6 = (~(Cxxmz6[10] & Edqhw6));
assign Wlh8v6 = (~(M8shw6 & T8shw6));
assign T8shw6 = (A9shw6 & H9shw6);
assign H9shw6 = (~(Ikxmz6[3] & Obqhw6));
assign A9shw6 = (O9shw6 & V9shw6);
assign V9shw6 = (~(Cxxmz6[12] & Nkrhw6));
assign O9shw6 = (~(Krxmz6[11] & Hbqhw6));
assign M8shw6 = (Cashw6 & Jashw6);
assign Jashw6 = (~(Cxxmz6[11] & Edqhw6));
assign Cashw6 = (~(Coxmz6[11] & Jcqhw6));
assign Plh8v6 = (~(Qashw6 & Xashw6));
assign Xashw6 = (Ebshw6 & Lbshw6);
assign Lbshw6 = (~(Krxmz6[12] & Hbqhw6));
assign Ebshw6 = (Sbshw6 & Ejrhw6);
assign Sbshw6 = (~(Cxxmz6[13] & Nkrhw6));
assign Qashw6 = (Zbshw6 & Gcshw6);
assign Gcshw6 = (~(Coxmz6[12] & Jcqhw6));
assign Zbshw6 = (Ncshw6 & Ucshw6);
assign Ucshw6 = (~(Njxmz6[0] & Obqhw6));
assign Ncshw6 = (~(Cxxmz6[12] & Edqhw6));
assign Ilh8v6 = (~(Bdshw6 & Idshw6));
assign Idshw6 = (Pdshw6 & Wdshw6);
assign Wdshw6 = (~(Njxmz6[1] & Obqhw6));
assign Pdshw6 = (Deshw6 & Keshw6);
assign Keshw6 = (~(Cxxmz6[14] & Nkrhw6));
assign Deshw6 = (~(Krxmz6[13] & Hbqhw6));
assign Bdshw6 = (Reshw6 & Yeshw6);
assign Yeshw6 = (~(Cxxmz6[13] & Edqhw6));
assign Reshw6 = (~(Coxmz6[13] & Jcqhw6));
assign Blh8v6 = (~(Ffshw6 & Mfshw6));
assign Mfshw6 = (Tfshw6 & Agshw6);
assign Agshw6 = (~(Njxmz6[2] & Obqhw6));
assign Tfshw6 = (Hgshw6 & Ogshw6);
assign Ogshw6 = (~(Cxxmz6[15] & Nkrhw6));
assign Hgshw6 = (~(Krxmz6[14] & Hbqhw6));
assign Ffshw6 = (Vgshw6 & Chshw6);
assign Chshw6 = (~(Cxxmz6[14] & Edqhw6));
assign Vgshw6 = (~(Coxmz6[14] & Jcqhw6));
assign Ukh8v6 = (~(Jhshw6 & Qhshw6));
assign Qhshw6 = (Xhshw6 & Eishw6);
assign Eishw6 = (~(Njxmz6[3] & Obqhw6));
assign Xhshw6 = (Lishw6 & Sishw6);
assign Sishw6 = (~(Cxxmz6[16] & Nkrhw6));
assign Lishw6 = (~(Krxmz6[15] & Hbqhw6));
assign Jhshw6 = (Zishw6 & Gjshw6);
assign Gjshw6 = (~(Cxxmz6[15] & Edqhw6));
assign Zishw6 = (~(Coxmz6[15] & Jcqhw6));
assign Nkh8v6 = (~(Njshw6 & Ujshw6));
assign Ujshw6 = (Bkshw6 & Ikshw6);
assign Ikshw6 = (~(Njxmz6[4] & Obqhw6));
assign Bkshw6 = (Pkshw6 & Wkshw6);
assign Wkshw6 = (~(Cxxmz6[17] & Nkrhw6));
assign Pkshw6 = (~(Krxmz6[16] & Hbqhw6));
assign Njshw6 = (Dlshw6 & Klshw6);
assign Klshw6 = (~(Cxxmz6[16] & Edqhw6));
assign Dlshw6 = (~(Coxmz6[16] & Jcqhw6));
assign Gkh8v6 = (~(Rlshw6 & Ylshw6));
assign Ylshw6 = (Fmshw6 & Mmshw6);
assign Mmshw6 = (~(Njxmz6[5] & Obqhw6));
assign Fmshw6 = (Tmshw6 & Anshw6);
assign Anshw6 = (~(Cxxmz6[18] & Nkrhw6));
assign Tmshw6 = (~(Krxmz6[17] & Hbqhw6));
assign Rlshw6 = (Hnshw6 & Onshw6);
assign Onshw6 = (~(Cxxmz6[17] & Edqhw6));
assign Hnshw6 = (~(Coxmz6[17] & Jcqhw6));
assign Zjh8v6 = (~(Vnshw6 & Coshw6));
assign Coshw6 = (Joshw6 & Qoshw6);
assign Qoshw6 = (~(Njxmz6[6] & Obqhw6));
assign Joshw6 = (Xoshw6 & Epshw6);
assign Epshw6 = (~(Cxxmz6[19] & Nkrhw6));
assign Xoshw6 = (~(Krxmz6[18] & Hbqhw6));
assign Vnshw6 = (Lpshw6 & Spshw6);
assign Spshw6 = (~(Cxxmz6[18] & Edqhw6));
assign Lpshw6 = (~(Coxmz6[18] & Jcqhw6));
assign Sjh8v6 = (~(Zpshw6 & Gqshw6));
assign Gqshw6 = (Nqshw6 & Uqshw6);
assign Uqshw6 = (~(Njxmz6[7] & Obqhw6));
assign Nqshw6 = (Brshw6 & Irshw6);
assign Irshw6 = (~(Cxxmz6[20] & Nkrhw6));
assign Brshw6 = (~(Krxmz6[19] & Hbqhw6));
assign Zpshw6 = (Prshw6 & Wrshw6);
assign Wrshw6 = (~(Cxxmz6[19] & Edqhw6));
assign Prshw6 = (~(Coxmz6[19] & Jcqhw6));
assign Ljh8v6 = (~(Dsshw6 & Ksshw6));
assign Ksshw6 = (Rsshw6 & Ysshw6);
assign Ysshw6 = (~(Njxmz6[8] & Obqhw6));
assign Rsshw6 = (Ftshw6 & Mtshw6);
assign Mtshw6 = (~(Cxxmz6[21] & Nkrhw6));
assign Ftshw6 = (~(Krxmz6[20] & Hbqhw6));
assign Dsshw6 = (Ttshw6 & Aushw6);
assign Aushw6 = (~(Cxxmz6[20] & Edqhw6));
assign Ttshw6 = (~(Coxmz6[20] & Jcqhw6));
assign Ejh8v6 = (~(Hushw6 & Oushw6));
assign Oushw6 = (Vushw6 & Cvshw6);
assign Cvshw6 = (~(Krxmz6[21] & Hbqhw6));
assign Vushw6 = (Jvshw6 & Ejrhw6);
assign Jvshw6 = (~(Cxxmz6[22] & Nkrhw6));
assign Hushw6 = (Qvshw6 & Xvshw6);
assign Xvshw6 = (~(Coxmz6[21] & Jcqhw6));
assign Qvshw6 = (Ewshw6 & Lwshw6);
assign Lwshw6 = (~(Njxmz6[9] & Obqhw6));
assign Ewshw6 = (~(Cxxmz6[21] & Edqhw6));
assign Xih8v6 = (~(Swshw6 & Zwshw6));
assign Zwshw6 = (Gxshw6 & Nxshw6);
assign Nxshw6 = (~(Njxmz6[10] & Obqhw6));
assign Gxshw6 = (Uxshw6 & Byshw6);
assign Byshw6 = (~(Nkrhw6 & Cxxmz6[23]));
assign Uxshw6 = (~(Krxmz6[22] & Hbqhw6));
assign Swshw6 = (Iyshw6 & Pyshw6);
assign Pyshw6 = (~(Cxxmz6[22] & Edqhw6));
assign Iyshw6 = (~(Coxmz6[22] & Jcqhw6));
assign Qih8v6 = (~(Wyshw6 & Dzshw6));
assign Dzshw6 = (Kzshw6 & Rzshw6);
assign Rzshw6 = (~(Krxmz6[23] & Hbqhw6));
assign Kzshw6 = (Yzshw6 & Ejrhw6);
assign Yzshw6 = (~(Cxxmz6[24] & Nkrhw6));
assign Wyshw6 = (F0thw6 & M0thw6);
assign M0thw6 = (~(Coxmz6[23] & Jcqhw6));
assign F0thw6 = (T0thw6 & A1thw6);
assign A1thw6 = (~(Obqhw6 & Njxmz6[11]));
assign T0thw6 = (~(Cxxmz6[23] & Edqhw6));
assign Jih8v6 = (~(H1thw6 & O1thw6));
assign O1thw6 = (V1thw6 & C2thw6);
assign C2thw6 = (~(Krxmz6[24] & Hbqhw6));
assign V1thw6 = (J2thw6 & Ejrhw6);
assign J2thw6 = (~(Cxxmz6[25] & Nkrhw6));
assign H1thw6 = (Q2thw6 & X2thw6);
assign X2thw6 = (~(Cxxmz6[24] & Edqhw6));
assign Q2thw6 = (~(Coxmz6[24] & Jcqhw6));
assign Cih8v6 = (~(E3thw6 & L3thw6));
assign L3thw6 = (S3thw6 & Z3thw6);
assign Z3thw6 = (~(Krxmz6[25] & Hbqhw6));
assign S3thw6 = (G4thw6 & Ejrhw6);
assign G4thw6 = (~(Cxxmz6[26] & Nkrhw6));
assign E3thw6 = (N4thw6 & U4thw6);
assign U4thw6 = (~(Cxxmz6[25] & Edqhw6));
assign N4thw6 = (~(Coxmz6[25] & Jcqhw6));
assign Vhh8v6 = (~(B5thw6 & I5thw6));
assign I5thw6 = (P5thw6 & W5thw6);
assign W5thw6 = (~(Wk47v6 & Obqhw6));
assign P5thw6 = (D6thw6 & K6thw6);
assign K6thw6 = (~(Cxxmz6[27] & Nkrhw6));
assign D6thw6 = (~(Krxmz6[26] & Hbqhw6));
assign B5thw6 = (R6thw6 & Y6thw6);
assign Y6thw6 = (~(Cxxmz6[26] & Edqhw6));
assign R6thw6 = (~(Coxmz6[26] & Jcqhw6));
assign Ohh8v6 = (~(F7thw6 & M7thw6));
assign M7thw6 = (T7thw6 & A8thw6);
assign A8thw6 = (~(Krxmz6[27] & Hbqhw6));
assign T7thw6 = (H8thw6 & Ejrhw6);
assign H8thw6 = (~(Cxxmz6[28] & Nkrhw6));
assign F7thw6 = (O8thw6 & V8thw6);
assign V8thw6 = (~(Cxxmz6[27] & Edqhw6));
assign O8thw6 = (~(Coxmz6[27] & Jcqhw6));
assign Hhh8v6 = (~(C9thw6 & J9thw6));
assign J9thw6 = (Q9thw6 & X9thw6);
assign X9thw6 = (~(Obqhw6 & Qm47v6));
assign Q9thw6 = (Eathw6 & Lathw6);
assign Lathw6 = (~(Cxxmz6[29] & Nkrhw6));
assign Eathw6 = (~(Krxmz6[28] & Hbqhw6));
assign C9thw6 = (Sathw6 & Zathw6);
assign Zathw6 = (~(Cxxmz6[28] & Edqhw6));
assign Sathw6 = (~(Coxmz6[28] & Jcqhw6));
assign Ahh8v6 = (~(Gbthw6 & Nbthw6));
assign Nbthw6 = (Ubthw6 & Bcthw6);
assign Bcthw6 = (~(Krxmz6[29] & Hbqhw6));
assign Ubthw6 = (Icthw6 & Ejrhw6);
assign Icthw6 = (~(Cxxmz6[30] & Nkrhw6));
assign Gbthw6 = (Pcthw6 & Wcthw6);
assign Wcthw6 = (~(Coxmz6[29] & Jcqhw6));
assign Pcthw6 = (Ddthw6 & Kdthw6);
assign Kdthw6 = (~(Obqhw6 & Gj47v6));
assign Ddthw6 = (~(Cxxmz6[29] & Edqhw6));
assign Tgh8v6 = (~(Rdthw6 & Ydthw6));
assign Ydthw6 = (Fethw6 & Methw6);
assign Methw6 = (~(Obqhw6 & Sl47v6));
assign Fethw6 = (Tethw6 & Afthw6);
assign Afthw6 = (~(Nkrhw6 & Cxxmz6[31]));
assign Tethw6 = (~(Krxmz6[30] & Hbqhw6));
assign Rdthw6 = (Hfthw6 & Ofthw6);
assign Ofthw6 = (~(Cxxmz6[30] & Edqhw6));
assign Hfthw6 = (~(Coxmz6[30] & Jcqhw6));
assign Mgh8v6 = (~(Vfthw6 & Cgthw6));
assign Cgthw6 = (Jgthw6 & Qgthw6);
assign Qgthw6 = (Xgthw6 & Ejrhw6);
assign Ejrhw6 = (~(Ehthw6 & Lhthw6));
assign Ehthw6 = (Shthw6 & Zhthw6);
assign Xgthw6 = (~(Ovxmz6[0] & Ljrhw6));
assign Ljrhw6 = (Githw6 & Lhthw6);
assign Jgthw6 = (Nithw6 & Uithw6);
assign Uithw6 = (~(Coxmz6[0] & Gkrhw6));
assign Gkrhw6 = (Bjthw6 & Xh1nv6);
assign Bjthw6 = (Ijthw6 & Pjthw6);
assign Nithw6 = (~(Nkrhw6 & Cxxmz6[1]));
assign Nkrhw6 = (~(Edqhw6 | Wjthw6));
assign Vfthw6 = (Dkthw6 & Kkthw6);
assign Kkthw6 = (~(Edqhw6 & Cxxmz6[0]));
assign Edqhw6 = (!Ijthw6);
assign Dkthw6 = (Rkthw6 & Ykthw6);
assign Ykthw6 = (~(Krxmz6[0] & Hbqhw6));
assign Hbqhw6 = (Flthw6 & Cl57v6);
assign Flthw6 = (Lhthw6 & Zhthw6);
assign Rkthw6 = (~(Fy47v6 & Obqhw6));
assign Obqhw6 = (~(Mlthw6 | Pm57v6));
assign Mlthw6 = (!Exrhw6);
assign Exrhw6 = (Tlthw6 & Yn57v6);
assign Tlthw6 = (Lhthw6 & Shthw6);
assign Lhthw6 = (Amthw6 & Xh1nv6);
assign Amthw6 = (Ijthw6 & Hmthw6);
assign Ijthw6 = (~(Omthw6 & Vmthw6));
assign Vmthw6 = (~(Cnthw6 & Jnthw6));
assign Jnthw6 = (~(Qnthw6 & Xnthw6));
assign Xnthw6 = (~(Eothw6 & Lothw6));
assign Qnthw6 = (~(Sothw6 | Zothw6));
assign Cnthw6 = (Gpthw6 & Npthw6);
assign Omthw6 = (~(Upthw6 & Bqthw6));
assign Fgh8v6 = (Pqthw6 ? Iqthw6 : Ovxmz6[1]);
assign Iqthw6 = (Cxxmz6[1] | Uc1nv6);
assign Yfh8v6 = (Pqthw6 ? Wqthw6 : Fuxmz6[1]);
assign Wqthw6 = (Cxxmz6[9] & Uia7z6);
assign Rfh8v6 = (Drthw6 ? Hf57v6 : Ab57v6);
assign Kfh8v6 = (Ii57v6 ? Rrthw6 : Krthw6);
assign Rrthw6 = (Yrthw6 & Fsthw6);
assign Fsthw6 = (~(Msthw6 & Tsthw6));
assign Tsthw6 = (Bqthw6 & Hf57v6);
assign Msthw6 = (Eothw6 & Ds57v6);
assign Yrthw6 = (Atthw6 | Wd1nv6);
assign Krthw6 = (~(Atthw6 | Wd1nv6));
assign Dfh8v6 = (~(Htthw6 & Otthw6));
assign Otthw6 = (~(Vtthw6 & Npthw6));
assign Vtthw6 = (Cuthw6 | Juthw6);
assign Juthw6 = (Sdqhw6 ? Xuthw6 : Quthw6);
assign Cuthw6 = (~(Evthw6 & Lvthw6));
assign Lvthw6 = (Svthw6 | Zvthw6);
assign Zvthw6 = (~(Ii57v6 | Tg57v6));
assign Svthw6 = (Sdqhw6 ? Nwthw6 : Gwthw6);
assign Gwthw6 = (Uwthw6 & Bxthw6);
assign Evthw6 = (~(Ixthw6 & Pxthw6));
assign Ixthw6 = (~(Wxthw6 | Uzxmz6[3]));
assign Htthw6 = (~(Tq57v6 & Atthw6));
assign Weh8v6 = (~(Dythw6 & Kythw6));
assign Kythw6 = (~(Rythw6 & Yythw6));
assign Peh8v6 = (~(Dythw6 & Fzthw6));
assign Fzthw6 = (~(Rythw6 & Mzthw6));
assign Mzthw6 = (Tzthw6 ^ Yythw6);
assign Yythw6 = (!B1ymz6[0]);
assign Ieh8v6 = (A0uhw6 & H0uhw6);
assign H0uhw6 = (B1ymz6[2] ^ O0uhw6);
assign Beh8v6 = (A0uhw6 & V0uhw6);
assign V0uhw6 = (B1ymz6[3] ^ C1uhw6);
assign A0uhw6 = (Rythw6 & Dythw6);
assign Dythw6 = (~(J1uhw6 & Rythw6));
assign Udh8v6 = (Rythw6 & Q1uhw6);
assign Q1uhw6 = (B1ymz6[4] ^ X1uhw6);
assign Ndh8v6 = (Rythw6 & E2uhw6);
assign E2uhw6 = (B1ymz6[5] ^ L2uhw6);
assign L2uhw6 = (X1uhw6 & B1ymz6[4]);
assign X1uhw6 = (C1uhw6 & B1ymz6[3]);
assign C1uhw6 = (O0uhw6 & B1ymz6[2]);
assign O0uhw6 = (B1ymz6[0] & B1ymz6[1]);
assign Rythw6 = (Ifh7v6 & S2uhw6);
assign Gdh8v6 = (Z2uhw6 ? Woxmz6[1] : Fqxmz6[1]);
assign Z2uhw6 = (!G3uhw6);
assign Zch8v6 = (G3uhw6 ? Fqxmz6[2] : Woxmz6[2]);
assign Sch8v6 = (G3uhw6 ? Fqxmz6[3] : Woxmz6[3]);
assign Lch8v6 = (G3uhw6 | Woxmz6[4]);
assign Ech8v6 = (G3uhw6 ? Fqxmz6[5] : Woxmz6[5]);
assign Xbh8v6 = (G3uhw6 ? Fqxmz6[0] : Woxmz6[0]);
assign G3uhw6 = (N3uhw6 & Fqxmz6[4]);
assign N3uhw6 = (Fqxmz6[0] ? B4uhw6 : U3uhw6);
assign B4uhw6 = (I4uhw6 & P4uhw6);
assign P4uhw6 = (W4uhw6 & Fqxmz6[2]);
assign W4uhw6 = (Fqxmz6[1] & Uia7z6);
assign I4uhw6 = (Fqxmz6[5] & Fqxmz6[3]);
assign U3uhw6 = (D5uhw6 & K5uhw6);
assign K5uhw6 = (~(R5uhw6 | Fqxmz6[2]));
assign R5uhw6 = (Fqxmz6[3] | Fqxmz6[5]);
assign D5uhw6 = (~(Nc1nv6 | Fqxmz6[1]));
assign Qbh8v6 = (~(Y5uhw6 & F6uhw6));
assign F6uhw6 = (~(G8ymz6[1] & M6uhw6));
assign Y5uhw6 = (~(G8ymz6[2] & Nx1nv6));
assign Jbh8v6 = (T6uhw6 | A7uhw6);
assign T6uhw6 = (Nx1nv6 ? G8ymz6[1] : G8ymz6[0]);
assign Cbh8v6 = (~(H7uhw6 & O7uhw6));
assign O7uhw6 = (~(G8ymz6[2] & M6uhw6));
assign H7uhw6 = (~(G8ymz6[3] & Nx1nv6));
assign Vah8v6 = (~(V7uhw6 & C8uhw6));
assign C8uhw6 = (~(G8ymz6[3] & M6uhw6));
assign M6uhw6 = (~(Nx1nv6 | A7uhw6));
assign V7uhw6 = (~(Nx1nv6 & TDI));
assign Nx1nv6 = (D567v6 & R9ymz6[3]);
assign Oah8v6 = (~(J8uhw6 & Q8uhw6));
assign Q8uhw6 = (Iy1nv6 | Jo1nv6);
assign J8uhw6 = (~(X8uhw6 & G8ymz6[0]));
assign Hah8v6 = (~(E9uhw6 & L9uhw6));
assign L9uhw6 = (~(X8uhw6 & G8ymz6[1]));
assign E9uhw6 = (S9uhw6 & Cja7z6);
assign S9uhw6 = (Iy1nv6 | An1nv6);
assign Aah8v6 = (~(Z9uhw6 & Gauhw6));
assign Gauhw6 = (~(X8uhw6 & G8ymz6[2]));
assign Z9uhw6 = (Nauhw6 & Cja7z6);
assign Nauhw6 = (Iy1nv6 | Mm1nv6);
assign T9h8v6 = (~(Uauhw6 & Bbuhw6));
assign Bbuhw6 = (~(X8uhw6 & G8ymz6[3]));
assign Uauhw6 = (Ibuhw6 & Cja7z6);
assign Ibuhw6 = (Iy1nv6 | Pbuhw6);
assign Pbuhw6 = (!W6ymz6[3]);
assign Iy1nv6 = (X8uhw6 | Nc1nv6);
assign X8uhw6 = (Wbuhw6 & Lw1nv6);
assign Wbuhw6 = (R9ymz6[3] & R9ymz6[2]);
assign M9h8v6 = (~(Dcuhw6 & Kcuhw6));
assign Kcuhw6 = (~(Smwnv6 & L5ymz6[1]));
assign Dcuhw6 = (Rcuhw6 & Ycuhw6);
assign Ycuhw6 = (Fduhw6 | Mduhw6);
assign Rcuhw6 = (~(Lmwnv6 & L5ymz6[0]));
assign F9h8v6 = (~(Tduhw6 & Aeuhw6));
assign Aeuhw6 = (Heuhw6 & Oeuhw6);
assign Oeuhw6 = (~(Coxmz6[30] & Qlwnv6));
assign Heuhw6 = (Veuhw6 & Cfuhw6);
assign Veuhw6 = (~(Uixmz6[30] & Jlwnv6));
assign Tduhw6 = (Jfuhw6 & Qfuhw6);
assign Qfuhw6 = (~(Smwnv6 & L5ymz6[34]));
assign Jfuhw6 = (Xfuhw6 & Eguhw6);
assign Eguhw6 = (~(Okwnv6 & Mg47v6));
assign Xfuhw6 = (~(L5ymz6[33] & Lmwnv6));
assign Y8h8v6 = (~(Lguhw6 & Sguhw6));
assign Sguhw6 = (Zguhw6 & Ghuhw6);
assign Ghuhw6 = (~(Okwnv6 & Gj47v6));
assign Zguhw6 = (Nhuhw6 & Uhuhw6);
assign Uhuhw6 = (~(Uixmz6[29] & Jlwnv6));
assign Nhuhw6 = (~(Coxmz6[29] & Qlwnv6));
assign Lguhw6 = (Biuhw6 & Iiuhw6);
assign Iiuhw6 = (~(L5ymz6[32] & Lmwnv6));
assign Biuhw6 = (~(L5ymz6[33] & Smwnv6));
assign R8h8v6 = (~(Piuhw6 & Wiuhw6));
assign Wiuhw6 = (Djuhw6 & Kjuhw6);
assign Kjuhw6 = (~(Okwnv6 & Kh47v6));
assign Djuhw6 = (Rjuhw6 & Yjuhw6);
assign Yjuhw6 = (~(Uixmz6[28] & Jlwnv6));
assign Rjuhw6 = (~(Coxmz6[28] & Qlwnv6));
assign Piuhw6 = (Fkuhw6 & Mkuhw6);
assign Mkuhw6 = (~(L5ymz6[31] & Lmwnv6));
assign Fkuhw6 = (~(L5ymz6[32] & Smwnv6));
assign K8h8v6 = (~(Tkuhw6 & Aluhw6));
assign Aluhw6 = (Hluhw6 & Oluhw6);
assign Oluhw6 = (~(Coxmz6[27] & Qlwnv6));
assign Hluhw6 = (Vluhw6 & Cfuhw6);
assign Vluhw6 = (~(Uixmz6[27] & Jlwnv6));
assign Tkuhw6 = (Cmuhw6 & Jmuhw6);
assign Jmuhw6 = (~(L5ymz6[30] & Lmwnv6));
assign Cmuhw6 = (~(L5ymz6[31] & Smwnv6));
assign D8h8v6 = (~(Qmuhw6 & Xmuhw6));
assign Xmuhw6 = (Enuhw6 & Lnuhw6);
assign Lnuhw6 = (~(Qf47v6 & Okwnv6));
assign Enuhw6 = (Snuhw6 & Znuhw6);
assign Znuhw6 = (~(Uixmz6[26] & Jlwnv6));
assign Snuhw6 = (~(Coxmz6[26] & Qlwnv6));
assign Qmuhw6 = (Gouhw6 & Nouhw6);
assign Nouhw6 = (~(L5ymz6[29] & Lmwnv6));
assign Gouhw6 = (~(L5ymz6[30] & Smwnv6));
assign W7h8v6 = (~(Uouhw6 & Bpuhw6));
assign Bpuhw6 = (Ipuhw6 & Ppuhw6);
assign Ppuhw6 = (~(Coxmz6[25] & Qlwnv6));
assign Ipuhw6 = (Wpuhw6 & Cfuhw6);
assign Wpuhw6 = (~(Uixmz6[25] & Jlwnv6));
assign Uouhw6 = (Dquhw6 & Kquhw6);
assign Kquhw6 = (~(L5ymz6[28] & Lmwnv6));
assign Dquhw6 = (~(L5ymz6[29] & Smwnv6));
assign P7h8v6 = (~(Rquhw6 & Yquhw6));
assign Yquhw6 = (Fruhw6 & Mruhw6);
assign Mruhw6 = (~(Coxmz6[24] & Qlwnv6));
assign Fruhw6 = (Truhw6 & Cfuhw6);
assign Truhw6 = (~(Uixmz6[24] & Jlwnv6));
assign Rquhw6 = (Asuhw6 & Hsuhw6);
assign Hsuhw6 = (~(L5ymz6[27] & Lmwnv6));
assign Asuhw6 = (~(L5ymz6[28] & Smwnv6));
assign I7h8v6 = (~(Osuhw6 & Vsuhw6));
assign Vsuhw6 = (Ctuhw6 & Jtuhw6);
assign Jtuhw6 = (~(Okwnv6 & Tfxmz6[11]));
assign Ctuhw6 = (Qtuhw6 & Cfuhw6);
assign Qtuhw6 = (~(Coxmz6[23] & Qlwnv6));
assign Osuhw6 = (Xtuhw6 & Euuhw6);
assign Euuhw6 = (~(Lmwnv6 & L5ymz6[26]));
assign Xtuhw6 = (~(L5ymz6[27] & Smwnv6));
assign B7h8v6 = (~(Luuhw6 & Suuhw6));
assign Suuhw6 = (Zuuhw6 & Gvuhw6);
assign Gvuhw6 = (~(Coxmz6[22] & Qlwnv6));
assign Zuuhw6 = (~(Tfxmz6[10] & Okwnv6));
assign Luuhw6 = (Nvuhw6 & Uvuhw6);
assign Uvuhw6 = (~(L5ymz6[25] & Lmwnv6));
assign Nvuhw6 = (~(Smwnv6 & L5ymz6[26]));
assign U6h8v6 = (~(Bwuhw6 & Iwuhw6));
assign Iwuhw6 = (Pwuhw6 & Wwuhw6);
assign Wwuhw6 = (~(Tfxmz6[9] & Okwnv6));
assign Pwuhw6 = (Dxuhw6 & Cfuhw6);
assign Dxuhw6 = (~(Coxmz6[21] & Qlwnv6));
assign Bwuhw6 = (Kxuhw6 & Rxuhw6);
assign Rxuhw6 = (~(L5ymz6[24] & Lmwnv6));
assign Kxuhw6 = (~(L5ymz6[25] & Smwnv6));
assign N6h8v6 = (~(Yxuhw6 & Fyuhw6));
assign Fyuhw6 = (Myuhw6 & Tyuhw6);
assign Tyuhw6 = (~(Coxmz6[20] & Qlwnv6));
assign Myuhw6 = (~(Tfxmz6[8] & Okwnv6));
assign Yxuhw6 = (Azuhw6 & Hzuhw6);
assign Hzuhw6 = (~(L5ymz6[23] & Lmwnv6));
assign Azuhw6 = (~(L5ymz6[24] & Smwnv6));
assign G6h8v6 = (~(Ozuhw6 & Vzuhw6));
assign Vzuhw6 = (C0vhw6 & J0vhw6);
assign J0vhw6 = (~(Coxmz6[19] & Qlwnv6));
assign C0vhw6 = (~(Tfxmz6[7] & Okwnv6));
assign Ozuhw6 = (Q0vhw6 & X0vhw6);
assign X0vhw6 = (~(L5ymz6[22] & Lmwnv6));
assign Q0vhw6 = (~(L5ymz6[23] & Smwnv6));
assign Z5h8v6 = (~(E1vhw6 & L1vhw6));
assign L1vhw6 = (S1vhw6 & Z1vhw6);
assign Z1vhw6 = (~(Coxmz6[18] & Qlwnv6));
assign S1vhw6 = (~(Tfxmz6[6] & Okwnv6));
assign E1vhw6 = (G2vhw6 & N2vhw6);
assign N2vhw6 = (~(L5ymz6[21] & Lmwnv6));
assign G2vhw6 = (~(L5ymz6[22] & Smwnv6));
assign S5h8v6 = (~(U2vhw6 & B3vhw6));
assign B3vhw6 = (I3vhw6 & P3vhw6);
assign P3vhw6 = (~(Coxmz6[17] & Qlwnv6));
assign I3vhw6 = (~(Tfxmz6[5] & Okwnv6));
assign U2vhw6 = (W3vhw6 & D4vhw6);
assign D4vhw6 = (~(L5ymz6[20] & Lmwnv6));
assign W3vhw6 = (~(L5ymz6[21] & Smwnv6));
assign L5h8v6 = (~(K4vhw6 & R4vhw6));
assign R4vhw6 = (Y4vhw6 & F5vhw6);
assign F5vhw6 = (~(Coxmz6[16] & Qlwnv6));
assign Y4vhw6 = (~(Tfxmz6[4] & Okwnv6));
assign K4vhw6 = (M5vhw6 & T5vhw6);
assign T5vhw6 = (~(L5ymz6[19] & Lmwnv6));
assign M5vhw6 = (~(L5ymz6[20] & Smwnv6));
assign E5h8v6 = (~(A6vhw6 & H6vhw6));
assign H6vhw6 = (O6vhw6 & V6vhw6);
assign V6vhw6 = (~(Coxmz6[15] & Qlwnv6));
assign O6vhw6 = (~(Tfxmz6[3] & Okwnv6));
assign A6vhw6 = (C7vhw6 & J7vhw6);
assign J7vhw6 = (~(L5ymz6[18] & Lmwnv6));
assign C7vhw6 = (~(L5ymz6[19] & Smwnv6));
assign X4h8v6 = (~(Q7vhw6 & X7vhw6));
assign X7vhw6 = (E8vhw6 & L8vhw6);
assign L8vhw6 = (~(Coxmz6[14] & Qlwnv6));
assign E8vhw6 = (~(Tfxmz6[2] & Okwnv6));
assign Q7vhw6 = (S8vhw6 & Z8vhw6);
assign Z8vhw6 = (~(L5ymz6[17] & Lmwnv6));
assign S8vhw6 = (~(L5ymz6[18] & Smwnv6));
assign Q4h8v6 = (~(G9vhw6 & N9vhw6));
assign N9vhw6 = (U9vhw6 & Bavhw6);
assign Bavhw6 = (~(Coxmz6[13] & Qlwnv6));
assign U9vhw6 = (~(Tfxmz6[1] & Okwnv6));
assign G9vhw6 = (Iavhw6 & Pavhw6);
assign Pavhw6 = (~(L5ymz6[16] & Lmwnv6));
assign Iavhw6 = (~(L5ymz6[17] & Smwnv6));
assign J4h8v6 = (~(Wavhw6 & Dbvhw6));
assign Dbvhw6 = (Kbvhw6 & Rbvhw6);
assign Rbvhw6 = (~(Coxmz6[12] & Qlwnv6));
assign Kbvhw6 = (~(Tfxmz6[0] & Okwnv6));
assign Wavhw6 = (Ybvhw6 & Fcvhw6);
assign Fcvhw6 = (~(L5ymz6[15] & Lmwnv6));
assign Ybvhw6 = (~(L5ymz6[16] & Smwnv6));
assign C4h8v6 = (~(Mcvhw6 & Tcvhw6));
assign Tcvhw6 = (Advhw6 & Hdvhw6);
assign Hdvhw6 = (~(Coxmz6[11] & Qlwnv6));
assign Advhw6 = (~(Ogxmz6[3] & Okwnv6));
assign Mcvhw6 = (Odvhw6 & Vdvhw6);
assign Vdvhw6 = (~(L5ymz6[14] & Lmwnv6));
assign Odvhw6 = (~(L5ymz6[15] & Smwnv6));
assign V3h8v6 = (~(Cevhw6 & Jevhw6));
assign Jevhw6 = (Qevhw6 & Xevhw6);
assign Xevhw6 = (~(Ogxmz6[2] & Okwnv6));
assign Qevhw6 = (Efvhw6 & Cfuhw6);
assign Efvhw6 = (~(Coxmz6[10] & Qlwnv6));
assign Cevhw6 = (Lfvhw6 & Sfvhw6);
assign Sfvhw6 = (~(L5ymz6[13] & Lmwnv6));
assign Lfvhw6 = (~(L5ymz6[14] & Smwnv6));
assign O3h8v6 = (~(Zfvhw6 & Ggvhw6));
assign Ggvhw6 = (Ngvhw6 & Ugvhw6);
assign Ugvhw6 = (~(Coxmz6[9] & Qlwnv6));
assign Ngvhw6 = (~(Ogxmz6[1] & Okwnv6));
assign Zfvhw6 = (Bhvhw6 & Ihvhw6);
assign Ihvhw6 = (~(L5ymz6[12] & Lmwnv6));
assign Bhvhw6 = (~(L5ymz6[13] & Smwnv6));
assign H3h8v6 = (~(Phvhw6 & Whvhw6));
assign Whvhw6 = (Divhw6 & Kivhw6);
assign Kivhw6 = (~(Coxmz6[8] & Qlwnv6));
assign Divhw6 = (~(Ogxmz6[0] & Okwnv6));
assign Phvhw6 = (Rivhw6 & Yivhw6);
assign Yivhw6 = (~(L5ymz6[11] & Lmwnv6));
assign Rivhw6 = (~(L5ymz6[12] & Smwnv6));
assign A3h8v6 = (~(Fjvhw6 & Mjvhw6));
assign Mjvhw6 = (Tjvhw6 & Akvhw6);
assign Akvhw6 = (~(Uixmz6[7] & Jlwnv6));
assign Tjvhw6 = (~(Coxmz6[7] & Qlwnv6));
assign Fjvhw6 = (Hkvhw6 & Okvhw6);
assign Okvhw6 = (~(L5ymz6[10] & Lmwnv6));
assign Hkvhw6 = (~(L5ymz6[11] & Smwnv6));
assign T2h8v6 = (~(Vkvhw6 & Clvhw6));
assign Clvhw6 = (Jlvhw6 & Qlvhw6);
assign Qlvhw6 = (~(Coxmz6[6] & Qlwnv6));
assign Jlvhw6 = (Xlvhw6 & Cfuhw6);
assign Xlvhw6 = (~(Uixmz6[6] & Jlwnv6));
assign Vkvhw6 = (Emvhw6 & Lmvhw6);
assign Lmvhw6 = (~(L5ymz6[9] & Lmwnv6));
assign Emvhw6 = (~(L5ymz6[10] & Smwnv6));
assign M2h8v6 = (~(Smvhw6 & Zmvhw6));
assign Zmvhw6 = (Gnvhw6 & Nnvhw6);
assign Nnvhw6 = (~(Coxmz6[5] & Qlwnv6));
assign Gnvhw6 = (Unvhw6 & Cfuhw6);
assign Unvhw6 = (~(Uixmz6[5] & Jlwnv6));
assign Smvhw6 = (Bovhw6 & Iovhw6);
assign Iovhw6 = (~(L5ymz6[9] & Smwnv6));
assign Bovhw6 = (Povhw6 & Wovhw6);
assign Wovhw6 = (~(S067v6 & Okwnv6));
assign Povhw6 = (~(L5ymz6[8] & Lmwnv6));
assign F2h8v6 = (~(Dpvhw6 & Kpvhw6));
assign Kpvhw6 = (Rpvhw6 & Ypvhw6);
assign Ypvhw6 = (~(Coxmz6[4] & Qlwnv6));
assign Rpvhw6 = (Fqvhw6 & Cfuhw6);
assign Fqvhw6 = (~(Uixmz6[4] & Jlwnv6));
assign Jlwnv6 = (Mqvhw6 & Tqvhw6);
assign Tqvhw6 = (~(Mduhw6 | Q2ymz6[0]));
assign Mqvhw6 = (Uu57v6 & Q2ymz6[1]);
assign Dpvhw6 = (Arvhw6 & Hrvhw6);
assign Hrvhw6 = (~(L5ymz6[8] & Smwnv6));
assign Arvhw6 = (Orvhw6 & Vrvhw6);
assign Vrvhw6 = (~(F267v6 & Okwnv6));
assign Orvhw6 = (~(L5ymz6[7] & Lmwnv6));
assign Y1h8v6 = (~(Csvhw6 & Jsvhw6));
assign Jsvhw6 = (Qsvhw6 & Xsvhw6);
assign Xsvhw6 = (~(Coxmz6[3] & Qlwnv6));
assign Qsvhw6 = (~(Hhxmz6[1] & Okwnv6));
assign Csvhw6 = (Etvhw6 & Ltvhw6);
assign Ltvhw6 = (~(L5ymz6[6] & Lmwnv6));
assign Etvhw6 = (~(L5ymz6[7] & Smwnv6));
assign R1h8v6 = (~(Stvhw6 & Ztvhw6));
assign Ztvhw6 = (Guvhw6 & Nuvhw6);
assign Nuvhw6 = (~(Hhxmz6[0] & Okwnv6));
assign Guvhw6 = (Uuvhw6 & Cfuhw6);
assign Uuvhw6 = (~(Coxmz6[2] & Qlwnv6));
assign Stvhw6 = (Bvvhw6 & Ivvhw6);
assign Ivvhw6 = (~(L5ymz6[5] & Lmwnv6));
assign Bvvhw6 = (~(L5ymz6[6] & Smwnv6));
assign K1h8v6 = (~(Pvvhw6 & Wvvhw6));
assign Wvvhw6 = (Dwvhw6 & Kwvhw6);
assign Kwvhw6 = (~(Okwnv6 & Sx57v6));
assign Dwvhw6 = (Rwvhw6 & Cfuhw6);
assign Rwvhw6 = (~(Coxmz6[1] & Qlwnv6));
assign Pvvhw6 = (Ywvhw6 & Fxvhw6);
assign Fxvhw6 = (~(L5ymz6[4] & Lmwnv6));
assign Ywvhw6 = (~(L5ymz6[5] & Smwnv6));
assign D1h8v6 = (~(Mxvhw6 & Txvhw6));
assign Txvhw6 = (Ayvhw6 & Hyvhw6);
assign Hyvhw6 = (~(Okwnv6 & Ez57v6));
assign Okwnv6 = (Oyvhw6 & Vyvhw6);
assign Vyvhw6 = (~(Mduhw6 | Q2ymz6[1]));
assign Oyvhw6 = (Q2ymz6[0] & Uu57v6);
assign Ayvhw6 = (Czvhw6 & Cfuhw6);
assign Cfuhw6 = (~(Jzvhw6 & Qzvhw6));
assign Qzvhw6 = (W6ymz6[2] & W6ymz6[3]);
assign Jzvhw6 = (Xzvhw6 & Tm1nv6);
assign Czvhw6 = (~(Coxmz6[0] & Qlwnv6));
assign Qlwnv6 = (~(Mduhw6 | Uu57v6));
assign Mxvhw6 = (E0whw6 & L0whw6);
assign L0whw6 = (~(L5ymz6[3] & Lmwnv6));
assign E0whw6 = (~(L5ymz6[4] & Smwnv6));
assign W0h8v6 = (~(S0whw6 & Z0whw6));
assign Z0whw6 = (~(L5ymz6[2] & Lmwnv6));
assign S0whw6 = (~(L5ymz6[3] & Smwnv6));
assign P0h8v6 = (~(G1whw6 & N1whw6));
assign N1whw6 = (~(L5ymz6[2] & Smwnv6));
assign G1whw6 = (U1whw6 & B2whw6);
assign B2whw6 = (Mduhw6 | I2whw6);
assign Mduhw6 = (~(P2whw6 & Xzvhw6));
assign U1whw6 = (~(Lmwnv6 & L5ymz6[1]));
assign Lmwnv6 = (W2whw6 & Cja7z6);
assign Cja7z6 = (!Nc1nv6);
assign Nc1nv6 = (R9ymz6[0] & A7uhw6);
assign A7uhw6 = (!Pr1nv6);
assign Pr1nv6 = (~(D3whw6 & R9ymz6[3]));
assign D3whw6 = (R9ymz6[2] & R9ymz6[1]);
assign W2whw6 = (~(Smwnv6 | Xzvhw6));
assign Smwnv6 = (D567v6 & K3whw6);
assign D567v6 = (R3whw6 & R9ymz6[1]);
assign R3whw6 = (Nq1nv6 & Zp1nv6);
assign Zp1nv6 = (!R9ymz6[2]);
assign I0h8v6 = (Pqthw6 ? Y3whw6 : Fuxmz6[0]);
assign Y3whw6 = (Cxxmz6[8] & Uia7z6);
assign B0h8v6 = (~(F4whw6 & M4whw6));
assign M4whw6 = (~(T4whw6 & Uia7z6));
assign F4whw6 = (~(J1uhw6 & Uzxmz6[1]));
assign Uzg8v6 = (~(A5whw6 & H5whw6));
assign H5whw6 = (~(O5whw6 & Uia7z6));
assign A5whw6 = (~(J1uhw6 & Uzxmz6[2]));
assign Nzg8v6 = (~(V5whw6 & C6whw6));
assign C6whw6 = (~(J6whw6 & Uia7z6));
assign J6whw6 = (~(Q6whw6 & X6whw6));
assign X6whw6 = (E7whw6 & L7whw6);
assign L7whw6 = (S7whw6 & Z7whw6);
assign S7whw6 = (G8whw6 & N8whw6);
assign E7whw6 = (U8whw6 & B9whw6);
assign U8whw6 = (!Quthw6);
assign Q6whw6 = (I9whw6 & P9whw6);
assign P9whw6 = (W9whw6 & Dawhw6);
assign Dawhw6 = (~(Kawhw6 & Rawhw6));
assign Kawhw6 = (Tq57v6 & Yawhw6);
assign Yawhw6 = (~(Sdqhw6 & Fbwhw6));
assign W9whw6 = (~(Mbwhw6 & Tbwhw6));
assign I9whw6 = (Wjthw6 & Acwhw6);
assign Acwhw6 = (~(Xuthw6 & Hcwhw6));
assign V5whw6 = (~(J1uhw6 & Uzxmz6[3]));
assign Gzg8v6 = (~(Ocwhw6 & Vcwhw6));
assign Vcwhw6 = (~(Cdwhw6 & Uia7z6));
assign Ocwhw6 = (~(J1uhw6 & Uzxmz6[4]));
assign Zyg8v6 = (~(Jdwhw6 & Qdwhw6));
assign Qdwhw6 = (Xdwhw6 | Uc1nv6);
assign Jdwhw6 = (~(J1uhw6 & Uzxmz6[0]));
assign Syg8v6 = (!Eewhw6);
assign Eewhw6 = (Zewhw6 ? Sewhw6 : Lewhw6);
assign Lyg8v6 = (!Gfwhw6);
assign Gfwhw6 = (Myxmz6[1] ? Ufwhw6 : Nfwhw6);
assign Nfwhw6 = (Sewhw6 | Zewhw6);
assign Zewhw6 = (!Myxmz6[0]);
assign Eyg8v6 = (Myxmz6[2] ? Igwhw6 : Bgwhw6);
assign Igwhw6 = (~(Ufwhw6 & Pgwhw6));
assign Pgwhw6 = (Sewhw6 | Myxmz6[1]);
assign Ufwhw6 = (Lewhw6 & Wgwhw6);
assign Wgwhw6 = (Sewhw6 | Myxmz6[0]);
assign Bgwhw6 = (Dhwhw6 & Khwhw6);
assign Xxg8v6 = (Myxmz6[3] ? Yhwhw6 : Rhwhw6);
assign Yhwhw6 = (~(Lewhw6 & Fiwhw6));
assign Fiwhw6 = (Sewhw6 | Miwhw6);
assign Rhwhw6 = (Khwhw6 & Miwhw6);
assign Qxg8v6 = (Myxmz6[4] ? Ajwhw6 : Tiwhw6);
assign Ajwhw6 = (~(Lewhw6 & Hjwhw6));
assign Hjwhw6 = (~(Khwhw6 & Ojwhw6));
assign Tiwhw6 = (Khwhw6 & Vjwhw6);
assign Khwhw6 = (!Sewhw6);
assign Sewhw6 = (~(Lewhw6 & Uia7z6));
assign Lewhw6 = (~(Ckwhw6 & Uia7z6));
assign Ckwhw6 = (~(Jkwhw6 & Uzxmz6[0]));
assign Jxg8v6 = (Qkwhw6 ? Cl57v6 : S2uhw6);
assign Cxg8v6 = (Qkwhw6 ? Yn57v6 : Cl57v6);
assign Vwg8v6 = (~(Xkwhw6 & Elwhw6));
assign Elwhw6 = (~(Llwhw6 & Slwhw6));
assign Llwhw6 = (~(Zlwhw6 & Gmwhw6));
assign Gmwhw6 = (~(Nmwhw6 & Zothw6));
assign Nmwhw6 = (~(Umwhw6 | Uj57v6));
assign Zlwhw6 = (Wxthw6 | Bnwhw6);
assign Bnwhw6 = (Inwhw6 & Ldqhw6);
assign Xkwhw6 = (~(Uj57v6 & Pnwhw6));
assign Pnwhw6 = (~(Slwhw6 & Wnwhw6));
assign Wnwhw6 = (~(Zothw6 & Umwhw6));
assign Slwhw6 = (~(Qkwhw6 & Dowhw6));
assign Dowhw6 = (~(Kowhw6 & Npthw6));
assign Kowhw6 = (~(Rowhw6 & Yowhw6));
assign Yowhw6 = (~(Uzxmz6[0] & Fpwhw6));
assign Fpwhw6 = (~(Mpwhw6 & Tpwhw6));
assign Rowhw6 = (Aqwhw6 & Hqwhw6);
assign Aqwhw6 = (~(Oqwhw6 & Vqwhw6));
assign Vqwhw6 = (Tbwhw6 | Crwhw6);
assign Qkwhw6 = (Bxthw6 | J1uhw6);
assign Owg8v6 = (~(Uia7z6 & Jrwhw6));
assign Jrwhw6 = (~(Tg57v6 & Qrwhw6));
assign Qrwhw6 = (~(Xrwhw6 & Eothw6));
assign Hwg8v6 = (Drthw6 ? D857v6 : Eswhw6);
assign Drthw6 = (~(Lswhw6 & Sswhw6));
assign Sswhw6 = (Xdwhw6 & Cdwhw6);
assign Cdwhw6 = (~(Zswhw6 & Gtwhw6));
assign Gtwhw6 = (Ntwhw6 & Utwhw6);
assign Utwhw6 = (Buwhw6 & Z7whw6);
assign Buwhw6 = (~(Iuwhw6 | Puwhw6));
assign Ntwhw6 = (Wuwhw6 & Dvwhw6);
assign Zswhw6 = (Kvwhw6 & Rvwhw6);
assign Rvwhw6 = (Yvwhw6 & Fwwhw6);
assign Fwwhw6 = (~(Mwwhw6 & Og1nv6));
assign Mwwhw6 = (Twwhw6 & Axwhw6);
assign Yvwhw6 = (Hxwhw6 & Oxwhw6);
assign Oxwhw6 = (~(Crwhw6 & Og1nv6));
assign Hxwhw6 = (~(Vxwhw6 & Xuthw6));
assign Vxwhw6 = (!Hcwhw6);
assign Hcwhw6 = (Fuxmz6[1] | Fuxmz6[0]);
assign Kvwhw6 = (Wjthw6 & Cywhw6);
assign Cywhw6 = (~(Jywhw6 & Qywhw6));
assign Jywhw6 = (Xywhw6 & Ezwhw6);
assign Xdwhw6 = (Lzwhw6 & Szwhw6);
assign Szwhw6 = (Zzwhw6 & G0xhw6);
assign G0xhw6 = (N0xhw6 & N8whw6);
assign N0xhw6 = (~(Puwhw6 | Ei1nv6));
assign Zzwhw6 = (U0xhw6 & Wuwhw6);
assign U0xhw6 = (~(B1xhw6 & I1xhw6));
assign B1xhw6 = (~(Dvwhw6 & P1xhw6));
assign Lzwhw6 = (W1xhw6 & D2xhw6);
assign D2xhw6 = (K2xhw6 & R2xhw6);
assign R2xhw6 = (~(Rawhw6 & Tq57v6));
assign K2xhw6 = (Y2xhw6 & F3xhw6);
assign F3xhw6 = (~(Sdqhw6 & M3xhw6));
assign M3xhw6 = (~(T3xhw6 & A4xhw6));
assign A4xhw6 = (~(Jkwhw6 & Twwhw6));
assign T3xhw6 = (H4xhw6 & Mpwhw6);
assign H4xhw6 = (~(O4xhw6 & Oqwhw6));
assign Y2xhw6 = (V4xhw6 | Wjthw6);
assign W1xhw6 = (C5xhw6 & J5xhw6);
assign C5xhw6 = (Twwhw6 ? Inwhw6 : Q5xhw6);
assign Inwhw6 = (Bxthw6 & X5xhw6);
assign X5xhw6 = (~(E6xhw6 & Oqwhw6));
assign E6xhw6 = (Uzxmz6[1] & L6xhw6);
assign Q5xhw6 = (~(Uzxmz6[3] & S6xhw6));
assign S6xhw6 = (Uzxmz6[1] ^ Axwhw6);
assign Lswhw6 = (Z6xhw6 & G7xhw6);
assign G7xhw6 = (!T4whw6);
assign T4whw6 = (~(N7xhw6 & U7xhw6));
assign U7xhw6 = (B8xhw6 & I8xhw6);
assign I8xhw6 = (P8xhw6 & W8xhw6);
assign P8xhw6 = (~(D9xhw6 | Xh1nv6));
assign B8xhw6 = (K9xhw6 & R9xhw6);
assign R9xhw6 = (~(S2uhw6 & Y9xhw6));
assign Y9xhw6 = (~(Faxhw6 & Maxhw6));
assign Maxhw6 = (~(Taxhw6 & Twwhw6));
assign Faxhw6 = (Abxhw6 & Hbxhw6);
assign Hbxhw6 = (~(Obxhw6 & Tbwhw6));
assign Obxhw6 = (Vbxhw6 & Ccxhw6);
assign Abxhw6 = (~(Rawhw6 & Jcxhw6));
assign Jcxhw6 = (~(Ii57v6 & Tq57v6));
assign K9xhw6 = (Qcxhw6 & Uwthw6);
assign Qcxhw6 = (~(V4xhw6 & Gpthw6));
assign Gpthw6 = (!Wjthw6);
assign Wjthw6 = (Xcxhw6 & Ldqhw6);
assign Ldqhw6 = (~(Jkwhw6 & Tbwhw6));
assign Jkwhw6 = (!Tpwhw6);
assign Tpwhw6 = (~(Edxhw6 & Uzxmz6[4]));
assign Edxhw6 = (Uzxmz6[3] & Vbxhw6);
assign V4xhw6 = (Myxmz6[4] & Vjwhw6);
assign Vjwhw6 = (!Ojwhw6);
assign Ojwhw6 = (~(Myxmz6[3] & Miwhw6));
assign Miwhw6 = (Dhwhw6 & Myxmz6[2]);
assign Dhwhw6 = (Myxmz6[1] & Myxmz6[0]);
assign N7xhw6 = (Ldxhw6 & Sdxhw6);
assign Sdxhw6 = (Zdxhw6 & Gexhw6);
assign Gexhw6 = (Bxthw6 | Twwhw6);
assign Zdxhw6 = (Nexhw6 & Uexhw6);
assign Uexhw6 = (~(Puwhw6 & Ezwhw6));
assign Nexhw6 = (Dvwhw6 | Fuxmz6[1]);
assign Ldxhw6 = (J5xhw6 & P1xhw6);
assign P1xhw6 = (~(Xuthw6 & Fuxmz6[1]));
assign J5xhw6 = (Bfxhw6 & G8whw6);
assign G8whw6 = (~(Mbwhw6 & Crwhw6));
assign Bfxhw6 = (~(Crwhw6 & Uzxmz6[2]));
assign Z6xhw6 = (!O5whw6);
assign O5whw6 = (~(Ifxhw6 & Pfxhw6));
assign Pfxhw6 = (Wfxhw6 & Dgxhw6);
assign Dgxhw6 = (Kgxhw6 & Xcxhw6);
assign Xcxhw6 = (!Zothw6);
assign Zothw6 = (Taxhw6 & Uzxmz6[0]);
assign Kgxhw6 = (~(Pxthw6 | Rgxhw6));
assign Pxthw6 = (Ygxhw6 & Crwhw6);
assign Ygxhw6 = (Uzxmz6[2] & Axwhw6);
assign Wfxhw6 = (Fhxhw6 & Mhxhw6);
assign Mhxhw6 = (~(Thxhw6 & Xuthw6));
assign Xuthw6 = (Mbwhw6 & Aixhw6);
assign Mbwhw6 = (Uzxmz6[3] & Axwhw6);
assign Thxhw6 = (~(I1xhw6 | Fuxmz6[1]));
assign I1xhw6 = (!Fuxmz6[0]);
assign Fhxhw6 = (Bxthw6 & Z7whw6);
assign Bxthw6 = (~(Hixhw6 & Vbxhw6));
assign Ifxhw6 = (Oixhw6 & Vixhw6);
assign Vixhw6 = (Cjxhw6 & Wuwhw6);
assign Wuwhw6 = (~(Jjxhw6 & Uj1nv6));
assign Jjxhw6 = (Uzxmz6[2] & Twwhw6);
assign Cjxhw6 = (~(Qjxhw6 | D9xhw6));
assign D9xhw6 = (Qywhw6 & Xjxhw6);
assign Xjxhw6 = (~(Xywhw6 & Ezwhw6));
assign Ezwhw6 = (!Upthw6);
assign Xywhw6 = (Ekxhw6 | Fy47v6);
assign Qywhw6 = (!N8whw6);
assign N8whw6 = (~(Lkxhw6 & Skxhw6));
assign Skxhw6 = (Uzxmz6[1] & Uzxmz6[2]);
assign Lkxhw6 = (Uj1nv6 & Uzxmz6[0]);
assign Qjxhw6 = (!Dvwhw6);
assign Dvwhw6 = (~(Zkxhw6 & Tbwhw6));
assign Zkxhw6 = (Uj1nv6 & Uzxmz6[1]);
assign Oixhw6 = (Glxhw6 & Nlxhw6);
assign Nlxhw6 = (~(Ulxhw6 & Bmxhw6));
assign Bmxhw6 = (S2uhw6 & Fbwhw6);
assign Fbwhw6 = (!Ii57v6);
assign Ulxhw6 = (Rawhw6 & Tq57v6);
assign Rawhw6 = (!Mpwhw6);
assign Mpwhw6 = (~(Imxhw6 & Uzxmz6[1]));
assign Imxhw6 = (Og1nv6 & Axwhw6);
assign Glxhw6 = (B9whw6 & W8xhw6);
assign W8xhw6 = (~(Pmxhw6 & Iuwhw6));
assign Pmxhw6 = (Uzxmz6[0] & Uzxmz6[2]);
assign B9whw6 = (~(Upthw6 & Puwhw6));
assign Eswhw6 = (~(Wmxhw6 | Sothw6));
assign Wmxhw6 = (Dnxhw6 & Knxhw6);
assign Knxhw6 = (~(Yn57v6 & Rnxhw6));
assign Rnxhw6 = (Lothw6 | Pm57v6);
assign Awg8v6 = (Jcqhw6 | Ynxhw6);
assign Ynxhw6 = (Yt47v6 & Foxhw6);
assign Foxhw6 = (~(Xrwhw6 & Moxhw6));
assign Xrwhw6 = (~(Lothw6 | Tq57v6));
assign Tvg8v6 = (Zdqhw6 ? Omxmz6[25] : Cxxmz6[25]);
assign Mvg8v6 = (Zdqhw6 ? Omxmz6[26] : Cxxmz6[26]);
assign Fvg8v6 = (Zdqhw6 ? Omxmz6[27] : Cxxmz6[27]);
assign Yug8v6 = (Zdqhw6 ? Omxmz6[28] : Cxxmz6[28]);
assign Rug8v6 = (Zdqhw6 ? Omxmz6[29] : Cxxmz6[29]);
assign Zdqhw6 = (!Toxhw6);
assign Kug8v6 = (Toxhw6 ? Cxxmz6[30] : Omxmz6[30]);
assign Dug8v6 = (Toxhw6 ? Cxxmz6[4] : Omxmz6[4]);
assign Wtg8v6 = (Toxhw6 ? Cxxmz6[5] : Omxmz6[5]);
assign Ptg8v6 = (Toxhw6 ? Cxxmz6[6] : Omxmz6[6]);
assign Itg8v6 = (Toxhw6 ? Cxxmz6[7] : Omxmz6[7]);
assign Btg8v6 = (Toxhw6 ? Cxxmz6[0] : Pm57v6);
assign Usg8v6 = (~(Apxhw6 & Hpxhw6));
assign Hpxhw6 = (~(Cxxmz6[13] & Scrhw6));
assign Apxhw6 = (Opxhw6 & Vpxhw6);
assign Vpxhw6 = (~(Ndrhw6 & Njxmz6[1]));
assign Opxhw6 = (~(Udrhw6 & Hnxmz6[1]));
assign Nsg8v6 = (~(Cqxhw6 & Jqxhw6));
assign Jqxhw6 = (~(Cxxmz6[14] & Scrhw6));
assign Cqxhw6 = (Qqxhw6 & Xqxhw6);
assign Xqxhw6 = (~(Ndrhw6 & Njxmz6[2]));
assign Qqxhw6 = (~(Udrhw6 & Hnxmz6[2]));
assign Gsg8v6 = (~(Erxhw6 & Lrxhw6));
assign Lrxhw6 = (~(Cxxmz6[15] & Scrhw6));
assign Erxhw6 = (Srxhw6 & Zrxhw6);
assign Zrxhw6 = (~(Ndrhw6 & Njxmz6[3]));
assign Srxhw6 = (~(Udrhw6 & Hnxmz6[3]));
assign Zrg8v6 = (~(Gsxhw6 & Nsxhw6));
assign Nsxhw6 = (~(Cxxmz6[16] & Scrhw6));
assign Gsxhw6 = (Usxhw6 & Btxhw6);
assign Btxhw6 = (~(Ndrhw6 & Njxmz6[4]));
assign Usxhw6 = (~(Udrhw6 & Hnxmz6[4]));
assign Srg8v6 = (~(Itxhw6 & Ptxhw6));
assign Ptxhw6 = (~(Cxxmz6[17] & Scrhw6));
assign Itxhw6 = (Wtxhw6 & Duxhw6);
assign Duxhw6 = (~(Ndrhw6 & Njxmz6[5]));
assign Wtxhw6 = (~(Udrhw6 & Hnxmz6[5]));
assign Lrg8v6 = (~(Kuxhw6 & Ruxhw6));
assign Ruxhw6 = (~(Cxxmz6[18] & Scrhw6));
assign Kuxhw6 = (Yuxhw6 & Fvxhw6);
assign Fvxhw6 = (~(Ndrhw6 & Njxmz6[6]));
assign Yuxhw6 = (~(Udrhw6 & Hnxmz6[6]));
assign Erg8v6 = (~(Mvxhw6 & Tvxhw6));
assign Tvxhw6 = (~(Cxxmz6[19] & Scrhw6));
assign Mvxhw6 = (Awxhw6 & Hwxhw6);
assign Hwxhw6 = (~(Ndrhw6 & Njxmz6[7]));
assign Awxhw6 = (~(Udrhw6 & Hnxmz6[7]));
assign Xqg8v6 = (~(Owxhw6 & Vwxhw6));
assign Vwxhw6 = (~(Cxxmz6[20] & Scrhw6));
assign Owxhw6 = (Cxxhw6 & Jxxhw6);
assign Jxxhw6 = (~(Ndrhw6 & Njxmz6[8]));
assign Cxxhw6 = (~(Udrhw6 & Hnxmz6[8]));
assign Qqg8v6 = (~(Qxxhw6 & Xxxhw6));
assign Xxxhw6 = (~(Cxxmz6[21] & Scrhw6));
assign Qxxhw6 = (Eyxhw6 & Lyxhw6);
assign Lyxhw6 = (~(Ndrhw6 & Njxmz6[9]));
assign Eyxhw6 = (~(Udrhw6 & Hnxmz6[9]));
assign Jqg8v6 = (~(Syxhw6 & Zyxhw6));
assign Zyxhw6 = (~(Cxxmz6[22] & Scrhw6));
assign Syxhw6 = (Gzxhw6 & Nzxhw6);
assign Nzxhw6 = (~(Ndrhw6 & Njxmz6[10]));
assign Gzxhw6 = (~(Udrhw6 & Hnxmz6[10]));
assign Cqg8v6 = (~(Uzxhw6 & B0yhw6));
assign B0yhw6 = (~(Cxxmz6[12] & Scrhw6));
assign Uzxhw6 = (I0yhw6 & P0yhw6);
assign P0yhw6 = (~(Ndrhw6 & Njxmz6[0]));
assign Ndrhw6 = (~(Udrhw6 | Scrhw6));
assign I0yhw6 = (~(Udrhw6 & Hnxmz6[0]));
assign Udrhw6 = (~(Yfrhw6 | Scrhw6));
assign Vpg8v6 = (W0yhw6 ? Blxmz6[0] : Cxxmz6[2]);
assign Opg8v6 = (W0yhw6 ? Blxmz6[1] : Cxxmz6[3]);
assign Hpg8v6 = (Z6qhw6 ? K1yhw6 : D1yhw6);
assign K1yhw6 = (Viqhw6 & R1yhw6);
assign Viqhw6 = (Y1yhw6 & F2yhw6);
assign F2yhw6 = (M2yhw6 & T2yhw6);
assign T2yhw6 = (~(A3yhw6 & H3yhw6));
assign H3yhw6 = (~(O3yhw6 & V3yhw6));
assign V3yhw6 = (C4yhw6 & J4yhw6);
assign J4yhw6 = (Q4yhw6 & X4yhw6);
assign X4yhw6 = (~(E5yhw6 ^ L5yhw6));
assign Q4yhw6 = (~(S5yhw6 ^ Z5yhw6));
assign C4yhw6 = (G6yhw6 & N6yhw6);
assign N6yhw6 = (~(U6yhw6 ^ B7yhw6));
assign G6yhw6 = (~(I7yhw6 ^ P7yhw6));
assign O3yhw6 = (W7yhw6 & D8yhw6);
assign D8yhw6 = (K8yhw6 & R8yhw6);
assign R8yhw6 = (~(Y8yhw6 ^ F9yhw6));
assign K8yhw6 = (M9yhw6 ^ T9yhw6);
assign W7yhw6 = (Aayhw6 & Hayhw6);
assign Hayhw6 = (~(Oayhw6 ^ Qswnv6));
assign Aayhw6 = (~(Vayhw6 ^ Cbyhw6));
assign A3yhw6 = (Dz1nv6 ? Ikxmz6[0] : Ogxmz6[0]);
assign M2yhw6 = (~(Jbyhw6 & Qbyhw6));
assign Qbyhw6 = (~(Xbyhw6 & Ecyhw6));
assign Ecyhw6 = (Lcyhw6 & Scyhw6);
assign Scyhw6 = (Zcyhw6 & Gdyhw6);
assign Gdyhw6 = (~(Ndyhw6 ^ Udyhw6));
assign Zcyhw6 = (~(Beyhw6 ^ Ieyhw6));
assign Lcyhw6 = (Peyhw6 & Weyhw6);
assign Weyhw6 = (~(Dfyhw6 ^ Kfyhw6));
assign Peyhw6 = (~(Rfyhw6 ^ Yfyhw6));
assign Xbyhw6 = (Fgyhw6 & Mgyhw6);
assign Mgyhw6 = (Tgyhw6 & Ahyhw6);
assign Ahyhw6 = (~(Hhyhw6 ^ Ohyhw6));
assign Tgyhw6 = (~(Vhyhw6 ^ Ciyhw6));
assign Fgyhw6 = (Jiyhw6 & Qiyhw6);
assign Qiyhw6 = (~(Xiyhw6 ^ Ejyhw6));
assign Jiyhw6 = (~(Ljyhw6 ^ Sjyhw6));
assign Jbyhw6 = (Dz1nv6 ? Ikxmz6[2] : Ogxmz6[2]);
assign Y1yhw6 = (Zjyhw6 & Gkyhw6);
assign Gkyhw6 = (~(Nkyhw6 & Ukyhw6));
assign Ukyhw6 = (~(Blyhw6 & Ilyhw6));
assign Ilyhw6 = (Plyhw6 & Wlyhw6);
assign Wlyhw6 = (Dmyhw6 & Kmyhw6);
assign Kmyhw6 = (~(Rmyhw6 ^ Ymyhw6));
assign Dmyhw6 = (~(Fnyhw6 ^ Mnyhw6));
assign Plyhw6 = (Tnyhw6 & Aoyhw6);
assign Aoyhw6 = (~(Hoyhw6 ^ Mcwnv6));
assign Mcwnv6 = (Dz1nv6 ? Ulxmz6[31] : Aixmz6[31]);
assign Tnyhw6 = (~(Ooyhw6 ^ Voyhw6));
assign Blyhw6 = (Cpyhw6 & Jpyhw6);
assign Jpyhw6 = (Qpyhw6 & Xpyhw6);
assign Xpyhw6 = (~(Eqyhw6 ^ Lqyhw6));
assign Qpyhw6 = (~(Sqyhw6 ^ Zqyhw6));
assign Cpyhw6 = (Gryhw6 & Nryhw6);
assign Nryhw6 = (~(Uryhw6 ^ Bsyhw6));
assign Gryhw6 = (~(Isyhw6 ^ Psyhw6));
assign Nkyhw6 = (Dz1nv6 ? Ikxmz6[3] : Ogxmz6[3]);
assign Zjyhw6 = (~(Wsyhw6 & Dtyhw6));
assign Dtyhw6 = (~(Ktyhw6 & Rtyhw6));
assign Rtyhw6 = (Ytyhw6 & Fuyhw6);
assign Fuyhw6 = (Muyhw6 & Tuyhw6);
assign Tuyhw6 = (~(Avyhw6 ^ Hvyhw6));
assign Muyhw6 = (~(Ovyhw6 ^ Vvyhw6));
assign Ytyhw6 = (Cwyhw6 & Jwyhw6);
assign Jwyhw6 = (~(Qwyhw6 ^ Xwyhw6));
assign Cwyhw6 = (~(Exyhw6 ^ Lxyhw6));
assign Ktyhw6 = (Sxyhw6 & Zxyhw6);
assign Zxyhw6 = (Gyyhw6 & Nyyhw6);
assign Nyyhw6 = (~(Uyyhw6 ^ Bzyhw6));
assign Gyyhw6 = (~(Izyhw6 ^ Pzyhw6));
assign Sxyhw6 = (Wzyhw6 & D0zhw6);
assign D0zhw6 = (~(K0zhw6 ^ R0zhw6));
assign Wzyhw6 = (~(Y0zhw6 ^ F1zhw6));
assign Wsyhw6 = (Dz1nv6 ? Ikxmz6[1] : Ogxmz6[1]);
assign D1yhw6 = (Cp47v6 & M1zhw6);
assign M1zhw6 = (R1yhw6 | T1zhw6);
assign Apg8v6 = (W0yhw6 ? Ikxmz6[0] : Cxxmz6[8]);
assign Tog8v6 = (W0yhw6 ? Ikxmz6[1] : Cxxmz6[9]);
assign Mog8v6 = (W0yhw6 ? Ikxmz6[2] : Cxxmz6[10]);
assign W0yhw6 = (!Scrhw6);
assign Fog8v6 = (Scrhw6 ? Cxxmz6[11] : Ikxmz6[3]);
assign Yng8v6 = (Scrhw6 ? Cxxmz6[26] : Wk47v6);
assign Rng8v6 = (Scrhw6 ? Cxxmz6[28] : Qm47v6);
assign Kng8v6 = (Scrhw6 ? Cxxmz6[30] : Sl47v6);
assign Dng8v6 = (Scrhw6 ? Cxxmz6[0] : Fy47v6);
assign Scrhw6 = (A2zhw6 & H2zhw6);
assign H2zhw6 = (~(Pm57v6 | Cl57v6));
assign A2zhw6 = (O2zhw6 & Yn57v6);
assign Wmg8v6 = (V2zhw6 ? S657v6 : Tgrhw6);
assign Pmg8v6 = (~(C3zhw6 & J3zhw6));
assign J3zhw6 = (~(Q3zhw6 & X3zhw6));
assign X3zhw6 = (~(E4zhw6 | J1uhw6));
assign Q3zhw6 = (Fy47v6 & Puwhw6);
assign Puwhw6 = (!Ke1nv6);
assign Ke1nv6 = (~(L4zhw6 & Uj1nv6));
assign C3zhw6 = (~(V357v6 & S4zhw6));
assign S4zhw6 = (~(Cxxmz6[4] & Z4zhw6));
assign Img8v6 = (N5zhw6 ? G5zhw6 : Ud57v6);
assign N5zhw6 = (Npthw6 & U5zhw6);
assign U5zhw6 = (~(B6zhw6 & I6zhw6));
assign I6zhw6 = (P6zhw6 | Z7whw6);
assign P6zhw6 = (Wxthw6 | V357v6);
assign Wxthw6 = (~(S2uhw6 ^ Uj57v6));
assign B6zhw6 = (W6zhw6 & Perhw6);
assign W6zhw6 = (~(D7zhw6 & K7zhw6));
assign K7zhw6 = (Eothw6 & R7zhw6);
assign D7zhw6 = (Cxxmz6[3] & Y7zhw6);
assign G5zhw6 = (!F8zhw6);
assign Bmg8v6 = (~(M8zhw6 & T8zhw6));
assign T8zhw6 = (~(A9zhw6 & H9zhw6));
assign H9zhw6 = (O9zhw6 & Kp57v6);
assign O9zhw6 = (~(D857v6 | Ud57v6));
assign A9zhw6 = (V9zhw6 & Cazhw6);
assign M8zhw6 = (Jazhw6 | Qazhw6);
assign Jazhw6 = (V9zhw6 ? Eothw6 : Xazhw6);
assign Xazhw6 = (~(Perhw6 & Werhw6));
assign Ulg8v6 = (Toxhw6 ? Cxxmz6[24] : Ebzhw6);
assign Toxhw6 = (Lbzhw6 & O2zhw6);
assign Lbzhw6 = (Cl57v6 & Zhthw6);
assign Ebzhw6 = (!S397z6);
assign Nlg8v6 = (Pqthw6 ? Sbzhw6 : Ovxmz6[0]);
assign Pqthw6 = (~(Zbzhw6 & Uia7z6));
assign Zbzhw6 = (~(Githw6 & O2zhw6));
assign O2zhw6 = (Gczhw6 & Nczhw6);
assign Nczhw6 = (Uczhw6 & Gj1nv6);
assign Uczhw6 = (~(Kp57v6 | Ud57v6));
assign Gczhw6 = (F8zhw6 & V9zhw6);
assign Githw6 = (Bdzhw6 & Pm57v6);
assign Bdzhw6 = (Yn57v6 & Shthw6);
assign Shthw6 = (!Cl57v6);
assign Sbzhw6 = (Cxxmz6[0] | Uc1nv6);
assign Glg8v6 = (~(Idzhw6 & Pdzhw6));
assign Pdzhw6 = (~(Uz47v6 & Wdzhw6));
assign Wdzhw6 = (~(Dfrhw6 & Dezhw6));
assign Idzhw6 = (Dezhw6 | Umwhw6);
assign Umwhw6 = (!Cxxmz6[0]);
assign Dezhw6 = (~(Kezhw6 & Rezhw6));
assign Rezhw6 = (Yezhw6 & Npthw6);
assign Yezhw6 = (~(Tq57v6 | Ud57v6));
assign Kezhw6 = (Ffzhw6 & F8zhw6);
assign F8zhw6 = (Z7whw6 & Perhw6);
assign Perhw6 = (~(Lc57v6 & Mfzhw6));
assign Mfzhw6 = (~(Tfzhw6 & Agzhw6));
assign Agzhw6 = (~(Tgrhw6 & Hgzhw6));
assign Hgzhw6 = (~(V2zhw6 & P8qhw6));
assign P8qhw6 = (!Io47v6);
assign V2zhw6 = (Tgrhw6 ? Vgzhw6 : Ogzhw6);
assign Vgzhw6 = (~(Chzhw6 & Jhzhw6));
assign Jhzhw6 = (~(Qhzhw6 & Xhzhw6));
assign Chzhw6 = (Cp47v6 ? Qhzhw6 : Xhzhw6);
assign Ogzhw6 = (~(Eizhw6 & Cxxmz6[1]));
assign Eizhw6 = (Z4zhw6 & Qh1nv6);
assign Z4zhw6 = (Lizhw6 & V9zhw6);
assign Lizhw6 = (Eothw6 & Wd1nv6);
assign Tfzhw6 = (Hhrhw6 & Sizhw6);
assign Sizhw6 = (~(Zizhw6 & Gjzhw6));
assign Gjzhw6 = (Hmthw6 & Ccxhw6);
assign Zizhw6 = (Ab57v6 & Ei1nv6);
assign Ei1nv6 = (Aixhw6 & Uzxmz6[4]);
assign Aixhw6 = (O4xhw6 & Twwhw6);
assign O4xhw6 = (Vbxhw6 & L6xhw6);
assign Hhrhw6 = (Ohrhw6 | Hmthw6);
assign Ohrhw6 = (~(Njzhw6 & Ujzhw6));
assign Ujzhw6 = (Bkzhw6 & Yfrhw6);
assign Yfrhw6 = (!Tgrhw6);
assign Tgrhw6 = (R957v6 & Ek47v6);
assign Bkzhw6 = (~(Ikzhw6 & Pkzhw6));
assign Pkzhw6 = (Hmthw6 | Cazhw6);
assign Ikzhw6 = (~(Cxxmz6[2] & Eothw6));
assign Njzhw6 = (V9zhw6 & Gj1nv6);
assign Gj1nv6 = (Qh1nv6 & Wd1nv6);
assign V9zhw6 = (Wkzhw6 & Y7zhw6);
assign Wkzhw6 = (Hf57v6 & Npthw6);
assign Z7whw6 = (~(Dlzhw6 & Klzhw6));
assign Klzhw6 = (Uzxmz6[3] & L6xhw6);
assign Dlzhw6 = (Crwhw6 & Uzxmz6[4]);
assign Ffzhw6 = (Y7zhw6 & Eothw6);
assign Y7zhw6 = (Rlzhw6 & Taxhw6);
assign Taxhw6 = (!Hqwhw6);
assign Hqwhw6 = (~(Li1nv6 & Uzxmz6[4]));
assign Li1nv6 = (Og1nv6 & Vbxhw6);
assign Og1nv6 = (~(Ccxhw6 | L6xhw6));
assign Rlzhw6 = (Lothw6 & Twwhw6);
assign Zkg8v6 = (Kfrhw6 ? On47v6 : Ylzhw6);
assign Ylzhw6 = (M257v6 & E157v6);
assign Skg8v6 = (Kfrhw6 ? Omxmz6[2] : Fmzhw6);
assign Kfrhw6 = (!Mmzhw6);
assign Fmzhw6 = (M257v6 ? Usxmz6[0] : Yn57v6);
assign Lkg8v6 = (Mmzhw6 ? Tmzhw6 : Omxmz6[3]);
assign Mmzhw6 = (Dfrhw6 & Wy1nv6);
assign Wy1nv6 = (Anzhw6 & Hnzhw6);
assign Anzhw6 = (~(Onzhw6 & Vnzhw6));
assign Vnzhw6 = (~(Cazhw6 & Cozhw6));
assign Cozhw6 = (~(Werhw6 & Jozhw6));
assign Jozhw6 = (~(Qozhw6 & Xozhw6));
assign Xozhw6 = (Epzhw6 & E4zhw6);
assign E4zhw6 = (Sothw6 & R7zhw6);
assign Sothw6 = (Lpzhw6 & Spzhw6);
assign Spzhw6 = (~(H557v6 | Ud57v6));
assign Lpzhw6 = (~(V357v6 | S657v6));
assign Epzhw6 = (Qhzhw6 & Xhzhw6);
assign Xhzhw6 = (!Blxmz6[1]);
assign Qhzhw6 = (!Blxmz6[0]);
assign Qozhw6 = (Zpzhw6 & Ds57v6);
assign Zpzhw6 = (Kp57v6 & Bqthw6);
assign Cazhw6 = (Qm47v6 & Gj47v6);
assign Tmzhw6 = (M257v6 ? Usxmz6[1] : Cl57v6);
assign Ekg8v6 = (~(Gqzhw6 & Nqzhw6));
assign Nqzhw6 = (~(Uqzhw6 & Ymyhw6));
assign Gqzhw6 = (~(Cozet6 & Brzhw6));
assign Xjg8v6 = (~(Irzhw6 & Przhw6));
assign Przhw6 = (~(Uqzhw6 & Bsyhw6));
assign Irzhw6 = (~(Qmzet6 & Brzhw6));
assign Qjg8v6 = (~(Wrzhw6 & Dszhw6));
assign Dszhw6 = (~(Kszhw6 & Uqzhw6));
assign Kszhw6 = (~(T9yhw6 | Rszhw6));
assign Wrzhw6 = (~(Gco7z6[4] & Brzhw6));
assign Jjg8v6 = (Brzhw6 ? Gco7z6[5] : Rszhw6);
assign Cjg8v6 = (~(Yszhw6 ^ Bizet6));
assign Vig8v6 = (Zmwnv6 ? U3o7z6[12] : Bzyhw6);
assign Oig8v6 = (Zmwnv6 ? U3o7z6[13] : Hvyhw6);
assign Hig8v6 = (Zmwnv6 ? U3o7z6[14] : Pzyhw6);
assign Aig8v6 = (Zmwnv6 ? U3o7z6[15] : Xwyhw6);
assign Thg8v6 = (Zmwnv6 ? U3o7z6[16] : Sjyhw6);
assign Mhg8v6 = (Zmwnv6 ? U3o7z6[17] : Ejyhw6);
assign Fhg8v6 = (Zmwnv6 ? U3o7z6[18] : Yfyhw6);
assign Ygg8v6 = (Zmwnv6 ? U3o7z6[19] : Ieyhw6);
assign Rgg8v6 = (Zmwnv6 ? U3o7z6[20] : Ciyhw6);
assign Kgg8v6 = (Zmwnv6 ? U3o7z6[21] : Udyhw6);
assign Dgg8v6 = (Zmwnv6 ? U3o7z6[22] : Ohyhw6);
assign Wfg8v6 = (Zmwnv6 ? U3o7z6[23] : Kfyhw6);
assign Pfg8v6 = (Zmwnv6 ? U3o7z6[24] : Psyhw6);
assign Ifg8v6 = (~(Ftzhw6 & Mtzhw6));
assign Mtzhw6 = (~(Ttzhw6 & Bsyhw6));
assign Ftzhw6 = (~(U3o7z6[25] & Zmwnv6));
assign Bfg8v6 = (Zmwnv6 ? U3o7z6[26] : Voyhw6);
assign Ueg8v6 = (Zmwnv6 ? U3o7z6[27] : Mnyhw6);
assign Neg8v6 = (Zmwnv6 ? U3o7z6[28] : Lqyhw6);
assign Geg8v6 = (~(Auzhw6 & Huzhw6));
assign Huzhw6 = (~(Ttzhw6 & Ymyhw6));
assign Auzhw6 = (~(U3o7z6[29] & Zmwnv6));
assign Zdg8v6 = (Zmwnv6 ? U3o7z6[30] : Zqyhw6);
assign Sdg8v6 = (~(Ouzhw6 & Vuzhw6));
assign Vuzhw6 = (~(Cvzhw6 & Uqzhw6));
assign Uqzhw6 = (!Brzhw6);
assign Cvzhw6 = (Qswnv6 & Jvzhw6);
assign Ouzhw6 = (~(Pl0ft6 & Brzhw6));
assign Ldg8v6 = (Brzhw6 ? O7o7z6[2] : Qvzhw6);
assign Brzhw6 = (~(Xvzhw6 & Ewzhw6));
assign Ewzhw6 = (~(Lwzhw6 | Bmqhw6));
assign Bmqhw6 = (!Rnqhw6);
assign Xvzhw6 = (~(Ulqhw6 | Swzhw6));
assign Edg8v6 = (~(Zwzhw6 & Gxzhw6));
assign Gxzhw6 = (~(Yszhw6 & Y9o7z6[0]));
assign Zwzhw6 = (Nxzhw6 & Uxzhw6);
assign Uxzhw6 = (~(Ttzhw6 & Qswnv6));
assign Qswnv6 = (JTAGNSW ? Aixmz6[0] : Ulxmz6[0]);
assign Nxzhw6 = (~(Pj0ft6 & Byzhw6));
assign Xcg8v6 = (~(Iyzhw6 & Pyzhw6));
assign Pyzhw6 = (~(Qvzhw6 & Ttzhw6));
assign Iyzhw6 = (Wyzhw6 & Dzzhw6);
assign Dzzhw6 = (~(Ph0ft6 & Byzhw6));
assign Wyzhw6 = (~(Yszhw6 & Y9o7z6[1]));
assign Qcg8v6 = (~(Kzzhw6 & Rzzhw6));
assign Rzzhw6 = (~(Ttzhw6 & P7yhw6));
assign Kzzhw6 = (Yzzhw6 & F00iw6);
assign F00iw6 = (~(Pf0ft6 & Byzhw6));
assign Yzzhw6 = (~(Yszhw6 & Y9o7z6[2]));
assign Jcg8v6 = (~(M00iw6 & T00iw6));
assign T00iw6 = (~(Ttzhw6 & Z5yhw6));
assign M00iw6 = (A10iw6 & H10iw6);
assign H10iw6 = (~(Pd0ft6 & Byzhw6));
assign A10iw6 = (~(Yszhw6 & Y9o7z6[3]));
assign Ccg8v6 = (~(O10iw6 & V10iw6));
assign V10iw6 = (~(Yszhw6 & U3o7z6[4]));
assign O10iw6 = (C20iw6 & J20iw6);
assign J20iw6 = (Zmwnv6 | T9yhw6);
assign T9yhw6 = (!Q20iw6);
assign C20iw6 = (~(Pb0ft6 & Byzhw6));
assign Vbg8v6 = (~(X20iw6 & E30iw6));
assign E30iw6 = (~(Rszhw6 & Ttzhw6));
assign X20iw6 = (L30iw6 & S30iw6);
assign S30iw6 = (~(P90ft6 & Byzhw6));
assign L30iw6 = (~(Yszhw6 & U3o7z6[5]));
assign Obg8v6 = (~(Z30iw6 & G40iw6));
assign G40iw6 = (~(Ttzhw6 & F9yhw6));
assign Z30iw6 = (N40iw6 & U40iw6);
assign U40iw6 = (~(P70ft6 & Byzhw6));
assign N40iw6 = (~(Yszhw6 & U3o7z6[6]));
assign Hbg8v6 = (~(B50iw6 & I50iw6));
assign I50iw6 = (~(Ttzhw6 & B7yhw6));
assign B50iw6 = (P50iw6 & W50iw6);
assign W50iw6 = (~(P50ft6 & Byzhw6));
assign P50iw6 = (~(Yszhw6 & U3o7z6[7]));
assign Abg8v6 = (~(D60iw6 & K60iw6));
assign K60iw6 = (~(Ttzhw6 & F1zhw6));
assign D60iw6 = (R60iw6 & Y60iw6);
assign Y60iw6 = (~(P30ft6 & Byzhw6));
assign R60iw6 = (~(Yszhw6 & U3o7z6[8]));
assign Tag8v6 = (~(F70iw6 & M70iw6));
assign M70iw6 = (~(Ttzhw6 & R0zhw6));
assign F70iw6 = (T70iw6 & A80iw6);
assign A80iw6 = (~(P10ft6 & Byzhw6));
assign T70iw6 = (~(Yszhw6 & U3o7z6[9]));
assign Mag8v6 = (~(H80iw6 & O80iw6));
assign O80iw6 = (~(Ttzhw6 & Lxyhw6));
assign H80iw6 = (V80iw6 & C90iw6);
assign C90iw6 = (~(Pzzet6 & Byzhw6));
assign V80iw6 = (~(Yszhw6 & U3o7z6[10]));
assign Fag8v6 = (~(J90iw6 & Q90iw6));
assign Q90iw6 = (~(Ttzhw6 & Vvyhw6));
assign J90iw6 = (X90iw6 & Ea0iw6);
assign Ea0iw6 = (~(Pxzet6 & Byzhw6));
assign Byzhw6 = (~(Yszhw6 | Ttzhw6));
assign Ttzhw6 = (!Zmwnv6);
assign X90iw6 = (~(Yszhw6 & U3o7z6[11]));
assign Yszhw6 = (La0iw6 & Zmwnv6);
assign Zmwnv6 = (~(Sa0iw6 & Za0iw6));
assign Za0iw6 = (Rnqhw6 & Ulqhw6);
assign Rnqhw6 = (Gb0iw6 & Kr97z6);
assign Gb0iw6 = (Kgqhw6 & Ekqhw6);
assign Ekqhw6 = (!Dbymz6[1]);
assign Sa0iw6 = (~(Swzhw6 | Lwzhw6));
assign La0iw6 = (~(Nb0iw6 & Ub0iw6));
assign Ub0iw6 = (Gco7z6[5] ? Ic0iw6 : Bc0iw6);
assign Bc0iw6 = (Pc0iw6 & Gco7z6[4]);
assign Nb0iw6 = (Oeo7z6[2] & Wc0iw6);
assign Y9g8v6 = (~(Dd0iw6 & Kd0iw6));
assign Kd0iw6 = (~(I2yet6 & Y2qhw6));
assign Dd0iw6 = (Rd0iw6 & Yd0iw6);
assign Yd0iw6 = (~(Fe0iw6 & L3bdt6));
assign Rd0iw6 = (~(R2qhw6 & Lhmov6));
assign R9g8v6 = (Me0iw6 ? Vayhw6 : Coxmz6[1]);
assign Vayhw6 = (~(Te0iw6 & Af0iw6));
assign Af0iw6 = (Hf0iw6 & Of0iw6);
assign Hf0iw6 = (~(O7o7z6[2] & Vf0iw6));
assign Te0iw6 = (Cg0iw6 & Jg0iw6);
assign Jg0iw6 = (~(Itb7z6[1] & Qg0iw6));
assign Cg0iw6 = (~(Y9o7z6[1] & Xg0iw6));
assign K9g8v6 = (Jcqhw6 ? Coxmz6[1] : Krxmz6[1]);
assign D9g8v6 = (Me0iw6 ? I7yhw6 : Coxmz6[2]);
assign I7yhw6 = (~(Eh0iw6 & Lh0iw6));
assign Lh0iw6 = (~(Itb7z6[2] & Qg0iw6));
assign Eh0iw6 = (~(Y9o7z6[2] & Xg0iw6));
assign W8g8v6 = (Jcqhw6 ? Coxmz6[2] : Krxmz6[2]);
assign P8g8v6 = (Me0iw6 ? S5yhw6 : Coxmz6[3]);
assign S5yhw6 = (~(Sh0iw6 & Zh0iw6));
assign Zh0iw6 = (~(Itb7z6[3] & Qg0iw6));
assign Sh0iw6 = (~(Y9o7z6[3] & Xg0iw6));
assign I8g8v6 = (Jcqhw6 ? Coxmz6[3] : Krxmz6[3]);
assign B8g8v6 = (Me0iw6 ? M9yhw6 : Coxmz6[4]);
assign M9yhw6 = (~(Gi0iw6 & Ni0iw6));
assign Ni0iw6 = (Ui0iw6 & Bj0iw6);
assign Ui0iw6 = (~(Gco7z6[4] & Vf0iw6));
assign Gi0iw6 = (Ij0iw6 & Pj0iw6);
assign Pj0iw6 = (~(Itb7z6[4] & Qg0iw6));
assign Ij0iw6 = (~(U3o7z6[4] & Xg0iw6));
assign U7g8v6 = (Jcqhw6 ? Coxmz6[4] : Krxmz6[4]);
assign N7g8v6 = (Me0iw6 ? E5yhw6 : Coxmz6[5]);
assign E5yhw6 = (~(Wj0iw6 & Dk0iw6));
assign Dk0iw6 = (~(U3o7z6[5] & Xg0iw6));
assign Wj0iw6 = (Kk0iw6 & Rk0iw6);
assign Rk0iw6 = (~(Gco7z6[5] & Vf0iw6));
assign Kk0iw6 = (~(Itb7z6[5] & Qg0iw6));
assign G7g8v6 = (Jcqhw6 ? Coxmz6[5] : Krxmz6[5]);
assign Z6g8v6 = (Me0iw6 ? Y8yhw6 : Coxmz6[6]);
assign Y8yhw6 = (~(Yk0iw6 & Fl0iw6));
assign Fl0iw6 = (~(U3o7z6[6] & Xg0iw6));
assign Yk0iw6 = (Ml0iw6 & Tl0iw6);
assign Tl0iw6 = (~(Vf0iw6 & Gco7z6[6]));
assign Ml0iw6 = (~(Itb7z6[6] & Qg0iw6));
assign S6g8v6 = (Jcqhw6 ? Coxmz6[6] : Krxmz6[6]);
assign L6g8v6 = (Me0iw6 ? U6yhw6 : Coxmz6[7]);
assign U6yhw6 = (~(Am0iw6 & Hm0iw6));
assign Hm0iw6 = (~(U3o7z6[7] & Xg0iw6));
assign Am0iw6 = (Om0iw6 & Vm0iw6);
assign Vm0iw6 = (Cn0iw6 | L6qhw6);
assign Om0iw6 = (~(Itb7z6[7] & Qg0iw6));
assign E6g8v6 = (Jcqhw6 ? Coxmz6[7] : Krxmz6[7]);
assign X5g8v6 = (Me0iw6 ? Y0zhw6 : Coxmz6[8]);
assign Y0zhw6 = (~(Jn0iw6 & Qn0iw6));
assign Qn0iw6 = (~(Itb7z6[8] & Qg0iw6));
assign Jn0iw6 = (~(U3o7z6[8] & Xg0iw6));
assign Q5g8v6 = (Jcqhw6 ? Coxmz6[8] : Krxmz6[8]);
assign J5g8v6 = (Me0iw6 ? K0zhw6 : Coxmz6[9]);
assign K0zhw6 = (~(Xn0iw6 & Eo0iw6));
assign Eo0iw6 = (~(Itb7z6[9] & Qg0iw6));
assign Xn0iw6 = (~(U3o7z6[9] & Xg0iw6));
assign C5g8v6 = (Jcqhw6 ? Coxmz6[9] : Krxmz6[9]);
assign V4g8v6 = (Me0iw6 ? Exyhw6 : Coxmz6[10]);
assign Exyhw6 = (~(Lo0iw6 & So0iw6));
assign So0iw6 = (~(Itb7z6[10] & Qg0iw6));
assign Lo0iw6 = (~(U3o7z6[10] & Xg0iw6));
assign O4g8v6 = (Jcqhw6 ? Coxmz6[10] : Krxmz6[10]);
assign H4g8v6 = (Me0iw6 ? Ovyhw6 : Coxmz6[11]);
assign Ovyhw6 = (~(Zo0iw6 & Gp0iw6));
assign Gp0iw6 = (~(Itb7z6[11] & Qg0iw6));
assign Zo0iw6 = (~(U3o7z6[11] & Xg0iw6));
assign A4g8v6 = (Jcqhw6 ? Coxmz6[11] : Krxmz6[11]);
assign T3g8v6 = (Me0iw6 ? Uyyhw6 : Coxmz6[12]);
assign Uyyhw6 = (~(Np0iw6 & Up0iw6));
assign Up0iw6 = (~(U3o7z6[12] & Xg0iw6));
assign Np0iw6 = (Bq0iw6 & Of0iw6);
assign Bq0iw6 = (~(Itb7z6[12] & Qg0iw6));
assign M3g8v6 = (Jcqhw6 ? Coxmz6[12] : Krxmz6[12]);
assign F3g8v6 = (Me0iw6 ? Avyhw6 : Coxmz6[13]);
assign Avyhw6 = (~(Iq0iw6 & Pq0iw6));
assign Pq0iw6 = (~(U3o7z6[13] & Xg0iw6));
assign Iq0iw6 = (Wq0iw6 & Of0iw6);
assign Wq0iw6 = (~(Itb7z6[13] & Qg0iw6));
assign Y2g8v6 = (Jcqhw6 ? Coxmz6[13] : Krxmz6[13]);
assign R2g8v6 = (Me0iw6 ? Izyhw6 : Coxmz6[14]);
assign Izyhw6 = (~(Dr0iw6 & Kr0iw6));
assign Kr0iw6 = (~(U3o7z6[14] & Xg0iw6));
assign Dr0iw6 = (Rr0iw6 & Of0iw6);
assign Rr0iw6 = (~(Itb7z6[14] & Qg0iw6));
assign K2g8v6 = (Jcqhw6 ? Coxmz6[14] : Krxmz6[14]);
assign D2g8v6 = (Me0iw6 ? Qwyhw6 : Coxmz6[15]);
assign Qwyhw6 = (~(Yr0iw6 & Fs0iw6));
assign Fs0iw6 = (~(U3o7z6[15] & Xg0iw6));
assign Yr0iw6 = (Ms0iw6 & Of0iw6);
assign Ms0iw6 = (~(Itb7z6[15] & Qg0iw6));
assign W1g8v6 = (Jcqhw6 ? Coxmz6[15] : Krxmz6[15]);
assign P1g8v6 = (Me0iw6 ? Ljyhw6 : Coxmz6[16]);
assign Ljyhw6 = (~(Ts0iw6 & At0iw6));
assign At0iw6 = (~(U3o7z6[16] & Xg0iw6));
assign Ts0iw6 = (Ht0iw6 & Ot0iw6);
assign Ht0iw6 = (~(Itb7z6[16] & Qg0iw6));
assign I1g8v6 = (Jcqhw6 ? Coxmz6[16] : Krxmz6[16]);
assign B1g8v6 = (Me0iw6 ? Xiyhw6 : Coxmz6[17]);
assign Xiyhw6 = (~(Vt0iw6 & Cu0iw6));
assign Cu0iw6 = (~(U3o7z6[17] & Xg0iw6));
assign Vt0iw6 = (Ju0iw6 & Ot0iw6);
assign Ju0iw6 = (~(Itb7z6[17] & Qg0iw6));
assign U0g8v6 = (Jcqhw6 ? Coxmz6[17] : Krxmz6[17]);
assign N0g8v6 = (Me0iw6 ? Rfyhw6 : Coxmz6[18]);
assign Rfyhw6 = (~(Qu0iw6 & Xu0iw6));
assign Xu0iw6 = (~(U3o7z6[18] & Xg0iw6));
assign Qu0iw6 = (Ev0iw6 & Ot0iw6);
assign Ev0iw6 = (~(Itb7z6[18] & Qg0iw6));
assign G0g8v6 = (Jcqhw6 ? Coxmz6[18] : Krxmz6[18]);
assign Zzf8v6 = (Me0iw6 ? Beyhw6 : Coxmz6[19]);
assign Beyhw6 = (~(Lv0iw6 & Sv0iw6));
assign Sv0iw6 = (~(U3o7z6[19] & Xg0iw6));
assign Lv0iw6 = (Zv0iw6 & Of0iw6);
assign Zv0iw6 = (~(Itb7z6[19] & Qg0iw6));
assign Szf8v6 = (Jcqhw6 ? Coxmz6[19] : Krxmz6[19]);
assign Lzf8v6 = (Me0iw6 ? Vhyhw6 : Coxmz6[20]);
assign Vhyhw6 = (~(Gw0iw6 & Nw0iw6));
assign Nw0iw6 = (~(U3o7z6[20] & Xg0iw6));
assign Gw0iw6 = (Uw0iw6 & Bj0iw6);
assign Uw0iw6 = (~(Itb7z6[20] & Qg0iw6));
assign Ezf8v6 = (Jcqhw6 ? Coxmz6[20] : Krxmz6[20]);
assign Xyf8v6 = (Me0iw6 ? Ndyhw6 : Coxmz6[21]);
assign Ndyhw6 = (~(Bx0iw6 & Ix0iw6));
assign Ix0iw6 = (~(U3o7z6[21] & Xg0iw6));
assign Bx0iw6 = (Px0iw6 & Bj0iw6);
assign Px0iw6 = (~(Itb7z6[21] & Qg0iw6));
assign Qyf8v6 = (Jcqhw6 ? Coxmz6[21] : Krxmz6[21]);
assign Jyf8v6 = (Me0iw6 ? Hhyhw6 : Coxmz6[22]);
assign Hhyhw6 = (~(Wx0iw6 & Dy0iw6));
assign Dy0iw6 = (~(U3o7z6[22] & Xg0iw6));
assign Wx0iw6 = (Ky0iw6 & Bj0iw6);
assign Ky0iw6 = (~(Itb7z6[22] & Qg0iw6));
assign Cyf8v6 = (Jcqhw6 ? Coxmz6[22] : Krxmz6[22]);
assign Vxf8v6 = (Me0iw6 ? Dfyhw6 : Coxmz6[23]);
assign Dfyhw6 = (~(Ry0iw6 & Yy0iw6));
assign Yy0iw6 = (~(Itb7z6[23] & Qg0iw6));
assign Ry0iw6 = (~(U3o7z6[23] & Xg0iw6));
assign Oxf8v6 = (Jcqhw6 ? Coxmz6[23] : Krxmz6[23]);
assign Hxf8v6 = (Me0iw6 ? Isyhw6 : Coxmz6[24]);
assign Isyhw6 = (~(Fz0iw6 & Mz0iw6));
assign Mz0iw6 = (~(U3o7z6[24] & Xg0iw6));
assign Fz0iw6 = (Tz0iw6 & Cn0iw6);
assign Cn0iw6 = (!Vf0iw6);
assign Tz0iw6 = (~(Itb7z6[24] & Qg0iw6));
assign Axf8v6 = (Jcqhw6 ? Coxmz6[24] : Krxmz6[24]);
assign Twf8v6 = (Me0iw6 ? Uryhw6 : Coxmz6[25]);
assign Uryhw6 = (~(A01iw6 & H01iw6));
assign H01iw6 = (~(U3o7z6[25] & Xg0iw6));
assign A01iw6 = (O01iw6 & V01iw6);
assign V01iw6 = (~(Qmzet6 & Vf0iw6));
assign O01iw6 = (~(Itb7z6[25] & Qg0iw6));
assign Mwf8v6 = (Jcqhw6 ? Coxmz6[25] : Krxmz6[25]);
assign Fwf8v6 = (Me0iw6 ? Ooyhw6 : Coxmz6[26]);
assign Ooyhw6 = (~(C11iw6 & J11iw6));
assign J11iw6 = (~(U3o7z6[26] & Xg0iw6));
assign C11iw6 = (Q11iw6 & Bj0iw6);
assign Bj0iw6 = (Ot0iw6 | X11iw6);
assign Q11iw6 = (~(Itb7z6[26] & Qg0iw6));
assign Yvf8v6 = (Jcqhw6 ? Coxmz6[26] : Krxmz6[26]);
assign Rvf8v6 = (Me0iw6 ? Fnyhw6 : Coxmz6[27]);
assign Fnyhw6 = (~(E21iw6 & L21iw6));
assign L21iw6 = (~(Itb7z6[27] & Qg0iw6));
assign E21iw6 = (~(U3o7z6[27] & Xg0iw6));
assign Kvf8v6 = (Jcqhw6 ? Coxmz6[27] : Krxmz6[27]);
assign Dvf8v6 = (Me0iw6 ? Eqyhw6 : Coxmz6[28]);
assign Eqyhw6 = (~(S21iw6 & Z21iw6));
assign Z21iw6 = (~(Itb7z6[28] & Qg0iw6));
assign S21iw6 = (~(U3o7z6[28] & Xg0iw6));
assign Wuf8v6 = (Jcqhw6 ? Coxmz6[28] : Krxmz6[28]);
assign Puf8v6 = (Me0iw6 ? Rmyhw6 : Coxmz6[29]);
assign Rmyhw6 = (~(G31iw6 & N31iw6));
assign N31iw6 = (U31iw6 & Ot0iw6);
assign U31iw6 = (~(Cozet6 & Vf0iw6));
assign G31iw6 = (B41iw6 & I41iw6);
assign I41iw6 = (~(Itb7z6[29] & Qg0iw6));
assign B41iw6 = (~(U3o7z6[29] & Xg0iw6));
assign Iuf8v6 = (Jcqhw6 ? Coxmz6[29] : Krxmz6[29]);
assign Buf8v6 = (Me0iw6 ? Sqyhw6 : Coxmz6[30]);
assign Sqyhw6 = (~(P41iw6 & W41iw6));
assign W41iw6 = (~(U3o7z6[30] & Xg0iw6));
assign P41iw6 = (D51iw6 & Of0iw6);
assign D51iw6 = (~(Itb7z6[30] & Qg0iw6));
assign Utf8v6 = (Jcqhw6 ? Coxmz6[30] : Krxmz6[30]);
assign Ntf8v6 = (Me0iw6 ? Hoyhw6 : Coxmz6[31]);
assign Hoyhw6 = (~(K51iw6 & R51iw6));
assign R51iw6 = (~(U3o7z6[31] & Xg0iw6));
assign K51iw6 = (Y51iw6 & Of0iw6);
assign Of0iw6 = (Ot0iw6 | F5o7z6[2]);
assign Y51iw6 = (~(Itb7z6[31] & Qg0iw6));
assign Gtf8v6 = (Jcqhw6 ? Coxmz6[31] : Krxmz6[31]);
assign Zsf8v6 = (Me0iw6 ? Oayhw6 : Coxmz6[0]);
assign Me0iw6 = (Z6qhw6 & Lwzhw6);
assign Lwzhw6 = (!F61iw6);
assign Z6qhw6 = (M61iw6 & T61iw6);
assign T61iw6 = (Dbymz6[0] & Glqhw6);
assign Glqhw6 = (R0bdt6 | A71iw6);
assign A71iw6 = (!Kgqhw6);
assign M61iw6 = (Kr97z6 & Dbymz6[1]);
assign Oayhw6 = (~(H71iw6 & O71iw6));
assign O71iw6 = (V71iw6 & Ot0iw6);
assign Ot0iw6 = (~(C81iw6 & J81iw6));
assign J81iw6 = (Q81iw6 & F5o7z6[4]);
assign Q81iw6 = (F5o7z6[3] & Kgqhw6);
assign C81iw6 = (X81iw6 & F5o7z6[7]);
assign X81iw6 = (F5o7z6[6] & F5o7z6[5]);
assign V71iw6 = (~(Vf0iw6 & Pl0ft6));
assign Vf0iw6 = (E91iw6 & L91iw6);
assign E91iw6 = (S91iw6 & X11iw6);
assign H71iw6 = (Z91iw6 & Ga1iw6);
assign Ga1iw6 = (~(Itb7z6[0] & Qg0iw6));
assign Qg0iw6 = (~(Na1iw6 & Ua1iw6));
assign Ua1iw6 = (~(Bb1iw6 & F5o7z6[3]));
assign Na1iw6 = (~(Ib1iw6 & Kgqhw6));
assign Z91iw6 = (~(Y9o7z6[0] & Xg0iw6));
assign Xg0iw6 = (Bb1iw6 & L91iw6);
assign L91iw6 = (~(F5o7z6[3] | F5o7z6[4]));
assign Bb1iw6 = (F5o7z6[2] & S91iw6);
assign S91iw6 = (Pb1iw6 & Kgqhw6);
assign Ssf8v6 = (Jcqhw6 ? Coxmz6[0] : Krxmz6[0]);
assign Jcqhw6 = (Moxhw6 & Upthw6);
assign Upthw6 = (Ekxhw6 & Ds57v6);
assign Moxhw6 = (Bqthw6 & Pjthw6);
assign Pjthw6 = (~(Hmthw6 & Wb1iw6));
assign Wb1iw6 = (~(Yn57v6 & Cl57v6));
assign Hmthw6 = (!Kp57v6);
assign Lsf8v6 = (Kc1iw6 ? Sx57v6 : Dc1iw6);
assign Kc1iw6 = (Rc1iw6 & Yc1iw6);
assign Yc1iw6 = (~(Fd1iw6 & I2whw6));
assign I2whw6 = (!Fduhw6);
assign Fd1iw6 = (Xzvhw6 & Ez57v6);
assign Rc1iw6 = (~(Md1iw6 & Td1iw6));
assign Td1iw6 = (~(L5ymz6[3] & Ae1iw6));
assign Ae1iw6 = (!L5ymz6[4]);
assign Md1iw6 = (!He1iw6);
assign Esf8v6 = (Oe1iw6 & Hnzhw6);
assign Oe1iw6 = (~(Ve1iw6 & Cf1iw6));
assign Cf1iw6 = (~(Jf1iw6 & Qf1iw6));
assign Qf1iw6 = (Xf1iw6 & Eg1iw6);
assign Jf1iw6 = (Lg1iw6 & Kh47v6);
assign Lg1iw6 = (Gj47v6 & R9qhw6);
assign Ve1iw6 = (~(Sg1iw6 | S367v6));
assign Xrf8v6 = (~(Zg1iw6 & Gh1iw6));
assign Gh1iw6 = (~(Nh1iw6 & Uh1iw6));
assign Uh1iw6 = (Bi1iw6 & Ii1iw6);
assign Ii1iw6 = (Hw57v6 | Pi1iw6);
assign Pi1iw6 = (S367v6 & Hnzhw6);
assign Bi1iw6 = (Jo1nv6 & An1nv6);
assign An1nv6 = (!W6ymz6[1]);
assign Nh1iw6 = (By1nv6 & Co1nv6);
assign Zg1iw6 = (~(Hw57v6 & Hnzhw6));
assign Qrf8v6 = (~(Wi1iw6 & Dj1iw6));
assign Dj1iw6 = (~(Tfxmz6[1] & Diwnv6));
assign Wi1iw6 = (Kj1iw6 & Rj1iw6);
assign Rj1iw6 = (~(Hnxmz6[1] & Yiwnv6));
assign Kj1iw6 = (~(L5ymz6[16] & Fjwnv6));
assign Jrf8v6 = (~(Yj1iw6 & Fk1iw6));
assign Fk1iw6 = (~(Tfxmz6[2] & Diwnv6));
assign Yj1iw6 = (Mk1iw6 & Tk1iw6);
assign Tk1iw6 = (~(Hnxmz6[2] & Yiwnv6));
assign Mk1iw6 = (~(L5ymz6[17] & Fjwnv6));
assign Crf8v6 = (~(Al1iw6 & Hl1iw6));
assign Hl1iw6 = (~(Tfxmz6[3] & Diwnv6));
assign Al1iw6 = (Ol1iw6 & Vl1iw6);
assign Vl1iw6 = (~(Hnxmz6[3] & Yiwnv6));
assign Ol1iw6 = (~(L5ymz6[18] & Fjwnv6));
assign Vqf8v6 = (~(Cm1iw6 & Jm1iw6));
assign Jm1iw6 = (~(Tfxmz6[4] & Diwnv6));
assign Cm1iw6 = (Qm1iw6 & Xm1iw6);
assign Xm1iw6 = (~(Hnxmz6[4] & Yiwnv6));
assign Qm1iw6 = (~(L5ymz6[19] & Fjwnv6));
assign Oqf8v6 = (~(En1iw6 & Ln1iw6));
assign Ln1iw6 = (~(Tfxmz6[5] & Diwnv6));
assign En1iw6 = (Sn1iw6 & Zn1iw6);
assign Zn1iw6 = (~(Hnxmz6[5] & Yiwnv6));
assign Sn1iw6 = (~(L5ymz6[20] & Fjwnv6));
assign Hqf8v6 = (~(Go1iw6 & No1iw6));
assign No1iw6 = (~(Tfxmz6[6] & Diwnv6));
assign Go1iw6 = (Uo1iw6 & Bp1iw6);
assign Bp1iw6 = (~(Hnxmz6[6] & Yiwnv6));
assign Uo1iw6 = (~(L5ymz6[21] & Fjwnv6));
assign Aqf8v6 = (~(Ip1iw6 & Pp1iw6));
assign Pp1iw6 = (~(Tfxmz6[7] & Diwnv6));
assign Ip1iw6 = (Wp1iw6 & Dq1iw6);
assign Dq1iw6 = (~(Hnxmz6[7] & Yiwnv6));
assign Wp1iw6 = (~(L5ymz6[22] & Fjwnv6));
assign Tpf8v6 = (~(Kq1iw6 & Rq1iw6));
assign Rq1iw6 = (~(Tfxmz6[8] & Diwnv6));
assign Kq1iw6 = (Yq1iw6 & Fr1iw6);
assign Fr1iw6 = (~(Hnxmz6[8] & Yiwnv6));
assign Yq1iw6 = (~(L5ymz6[23] & Fjwnv6));
assign Mpf8v6 = (~(Mr1iw6 & Tr1iw6));
assign Tr1iw6 = (~(Tfxmz6[9] & Diwnv6));
assign Mr1iw6 = (As1iw6 & Hs1iw6);
assign Hs1iw6 = (~(Hnxmz6[9] & Yiwnv6));
assign As1iw6 = (~(L5ymz6[24] & Fjwnv6));
assign Fpf8v6 = (~(Os1iw6 & Vs1iw6));
assign Vs1iw6 = (~(Tfxmz6[10] & Diwnv6));
assign Os1iw6 = (Ct1iw6 & Jt1iw6);
assign Jt1iw6 = (~(Hnxmz6[10] & Yiwnv6));
assign Ct1iw6 = (~(L5ymz6[25] & Fjwnv6));
assign Yof8v6 = (~(Qt1iw6 & Xt1iw6));
assign Xt1iw6 = (~(Tfxmz6[0] & Diwnv6));
assign Qt1iw6 = (Eu1iw6 & Lu1iw6);
assign Lu1iw6 = (~(Hnxmz6[0] & Yiwnv6));
assign Yiwnv6 = (~(Diwnv6 | Su1iw6));
assign Eu1iw6 = (~(L5ymz6[15] & Fjwnv6));
assign Fjwnv6 = (~(Dc1iw6 | Diwnv6));
assign Diwnv6 = (Zu1iw6 & He1iw6);
assign Zu1iw6 = (~(W8qhw6 & Dc1iw6));
assign Rof8v6 = (Gv1iw6 ? F267v6 : W8qhw6);
assign Gv1iw6 = (Nv1iw6 & Uv1iw6);
assign Uv1iw6 = (~(L5ymz6[7] & B8qhw6));
assign B8qhw6 = (~(He1iw6 | W8qhw6));
assign Nv1iw6 = (Bw1iw6 | Iw1iw6);
assign Iw1iw6 = (Cp47v6 ? Hhxmz6[0] : Hhxmz6[1]);
assign Bw1iw6 = (~(W8qhw6 & Pw1iw6));
assign Pw1iw6 = (Hhxmz6[0] | Hhxmz6[1]);
assign Kof8v6 = (Iownv6 | Ww1iw6);
assign Ww1iw6 = (Dx1iw6 & Q7wnv6);
assign Dof8v6 = (~(Kx1iw6 & Rx1iw6));
assign Rx1iw6 = (~(Yx1iw6 & Unwnv6));
assign Kx1iw6 = (~(Iownv6 & Dtm7z6[0]));
assign Wnf8v6 = (~(Fy1iw6 & My1iw6));
assign My1iw6 = (~(Ty1iw6 & Unwnv6));
assign Unwnv6 = (~(Az1iw6 | Iownv6));
assign Ty1iw6 = (Hz1iw6 & Oz1iw6);
assign Fy1iw6 = (~(Iownv6 & Dtm7z6[1]));
assign Pnf8v6 = (~(Vz1iw6 & C02iw6));
assign C02iw6 = (~(Hl9ov6 & Fbqnv6));
assign Vz1iw6 = (~(Dq9ov6 & Styet6));
assign Inf8v6 = (~(J02iw6 & Q02iw6));
assign Q02iw6 = (~(T3qhw6 & X02iw6));
assign J02iw6 = (~(H4qhw6 & Znn7z6[0]));
assign Bnf8v6 = (~(E12iw6 & L12iw6));
assign L12iw6 = (~(T3qhw6 & S12iw6));
assign E12iw6 = (~(H4qhw6 & Znn7z6[2]));
assign Umf8v6 = (~(Z12iw6 & G22iw6));
assign G22iw6 = (~(T3qhw6 & N22iw6));
assign T3qhw6 = (~(U22iw6 | H4qhw6));
assign Z12iw6 = (~(H4qhw6 & Znn7z6[3]));
assign H4qhw6 = (Jalov6 & B32iw6);
assign Nmf8v6 = (Q7wnv6 ? FIXMASTERTYPE : Lq0ft6);
assign Gmf8v6 = (~(I32iw6 & P32iw6));
assign P32iw6 = (~(W32iw6 & Lxbet6));
assign I32iw6 = (D42iw6 | K42iw6);
assign Zlf8v6 = (!R42iw6);
assign R42iw6 = (W32iw6 ? F52iw6 : Y42iw6);
assign Y42iw6 = (~(M52iw6 & T52iw6));
assign Slf8v6 = (H62iw6 ? A62iw6 : Toi7z6[11]);
assign Llf8v6 = (H62iw6 ? O62iw6 : Toi7z6[10]);
assign Elf8v6 = (H62iw6 ? V62iw6 : Toi7z6[9]);
assign Xkf8v6 = (H62iw6 ? C72iw6 : Toi7z6[8]);
assign Qkf8v6 = (H62iw6 ? J72iw6 : Toi7z6[7]);
assign Jkf8v6 = (H62iw6 ? Q72iw6 : Toi7z6[6]);
assign Ckf8v6 = (H62iw6 ? X72iw6 : Toi7z6[5]);
assign H62iw6 = (!W32iw6);
assign Vjf8v6 = (W32iw6 ? Toi7z6[4] : E82iw6);
assign Ojf8v6 = (W32iw6 ? Toi7z6[3] : L82iw6);
assign Hjf8v6 = (W32iw6 ? Toi7z6[2] : S82iw6);
assign Ajf8v6 = (Z82iw6 & Lxbet6);
assign Z82iw6 = (~(G92iw6 | N92iw6));
assign Tif8v6 = (~(U92iw6 & Ba2iw6));
assign Ba2iw6 = (~(Ia2iw6 & Pa2iw6));
assign U92iw6 = (~(W32iw6 & Bqi7z6[3]));
assign Mif8v6 = (~(Wa2iw6 & Db2iw6));
assign Db2iw6 = (~(Ia2iw6 & Kb2iw6));
assign Wa2iw6 = (~(W32iw6 & Bqi7z6[2]));
assign Fif8v6 = (~(Rb2iw6 & Yb2iw6));
assign Yb2iw6 = (~(Ia2iw6 & Fc2iw6));
assign Rb2iw6 = (~(W32iw6 & Bqi7z6[1]));
assign Yhf8v6 = (~(Mc2iw6 & Tc2iw6));
assign Tc2iw6 = (~(Ia2iw6 & Ujlov6));
assign Ia2iw6 = (~(K42iw6 | Ad2iw6));
assign Mc2iw6 = (~(W32iw6 & Bqi7z6[0]));
assign W32iw6 = (K42iw6 & Hd2iw6);
assign Hd2iw6 = (~(Od2iw6 & Vd2iw6));
assign Od2iw6 = (~(Ce2iw6 & Je2iw6));
assign Ce2iw6 = (!Q22nv6);
assign K42iw6 = (Qe2iw6 | Xe2iw6);
assign Qe2iw6 = (~(Ef2iw6 & Vd2iw6));
assign Rhf8v6 = (~(Lf2iw6 & Sf2iw6));
assign Sf2iw6 = (~(Lgj7z6[11] & Zf2iw6));
assign Lf2iw6 = (~(Gg2iw6 & Ng2iw6));
assign Khf8v6 = (~(Ug2iw6 & Bh2iw6));
assign Bh2iw6 = (~(Lgj7z6[23] & Ih2iw6));
assign Ug2iw6 = (~(Ph2iw6 & Gg2iw6));
assign Dhf8v6 = (~(Wh2iw6 & Di2iw6));
assign Di2iw6 = (~(Lgj7z6[35] & Ki2iw6));
assign Wh2iw6 = (~(Ri2iw6 & Gg2iw6));
assign Wgf8v6 = (~(Yi2iw6 & Fj2iw6));
assign Fj2iw6 = (~(Lgj7z6[47] & Mj2iw6));
assign Yi2iw6 = (~(Tj2iw6 & Gg2iw6));
assign Pgf8v6 = (~(Ak2iw6 & Hk2iw6));
assign Hk2iw6 = (~(Lgj7z6[59] & Ok2iw6));
assign Ak2iw6 = (~(Vk2iw6 & Gg2iw6));
assign Igf8v6 = (~(Cl2iw6 & Jl2iw6));
assign Jl2iw6 = (~(Lgj7z6[71] & Ql2iw6));
assign Cl2iw6 = (~(Xl2iw6 & Gg2iw6));
assign Bgf8v6 = (~(Em2iw6 & Lm2iw6));
assign Lm2iw6 = (~(Lgj7z6[83] & Sm2iw6));
assign Em2iw6 = (~(Zm2iw6 & Gg2iw6));
assign Uff8v6 = (~(Gn2iw6 & Nn2iw6));
assign Nn2iw6 = (~(Lgj7z6[95] & Un2iw6));
assign Gn2iw6 = (~(Bo2iw6 & Gg2iw6));
assign Nff8v6 = (~(Io2iw6 & Po2iw6));
assign Po2iw6 = (~(Lgj7z6[107] & Wo2iw6));
assign Io2iw6 = (~(Dp2iw6 & Gg2iw6));
assign Gff8v6 = (~(Kp2iw6 & Rp2iw6));
assign Rp2iw6 = (~(Lgj7z6[119] & Yp2iw6));
assign Kp2iw6 = (~(Fq2iw6 & Gg2iw6));
assign Zef8v6 = (~(Mq2iw6 & Tq2iw6));
assign Tq2iw6 = (~(Lgj7z6[131] & Ar2iw6));
assign Mq2iw6 = (~(Hr2iw6 & Gg2iw6));
assign Sef8v6 = (~(Or2iw6 & Vr2iw6));
assign Vr2iw6 = (~(Lgj7z6[143] & Cs2iw6));
assign Or2iw6 = (~(Js2iw6 & Gg2iw6));
assign Lef8v6 = (~(Qs2iw6 & Xs2iw6));
assign Xs2iw6 = (~(Lgj7z6[155] & Et2iw6));
assign Qs2iw6 = (~(Lt2iw6 & Gg2iw6));
assign Eef8v6 = (~(St2iw6 & Zt2iw6));
assign Zt2iw6 = (~(Lgj7z6[167] & Gu2iw6));
assign St2iw6 = (~(Nu2iw6 & Gg2iw6));
assign Xdf8v6 = (~(Uu2iw6 & Bv2iw6));
assign Bv2iw6 = (~(Lgj7z6[179] & Iv2iw6));
assign Uu2iw6 = (~(Pv2iw6 & Gg2iw6));
assign Qdf8v6 = (~(Wv2iw6 & Dw2iw6));
assign Dw2iw6 = (~(Lgj7z6[191] & Kw2iw6));
assign Wv2iw6 = (~(Rw2iw6 & Gg2iw6));
assign Jdf8v6 = (~(Yw2iw6 & Fx2iw6));
assign Fx2iw6 = (~(Ohj7z6[63] & Mx2iw6));
assign Mx2iw6 = (~(Tx2iw6 & X0hov6));
assign Yw2iw6 = (~(Ay2iw6 & Gg2iw6));
assign Cdf8v6 = (~(Hy2iw6 & Oy2iw6));
assign Oy2iw6 = (~(Ohj7z6[31] & Vy2iw6));
assign Vy2iw6 = (~(Cz2iw6 & X0hov6));
assign Hy2iw6 = (~(Jz2iw6 & Gg2iw6));
assign Ocf8v6 = (~(Vcf8v6 & Qz2iw6));
assign Qz2iw6 = (~(P8adt6 & Xz2iw6));
assign Xz2iw6 = (~(O9adt6 & E03iw6));
assign E03iw6 = (Ef2iw6 | Xe2iw6);
assign Vcf8v6 = (~(L03iw6 & S03iw6));
assign S03iw6 = (O9adt6 & Vd2iw6);
assign L03iw6 = (~(Ef2iw6 | Xe2iw6));
assign Xe2iw6 = (~(Z03iw6 & G13iw6));
assign Z03iw6 = (~(N13iw6 | U13iw6));
assign Ef2iw6 = (~(B23iw6 & I23iw6));
assign I23iw6 = (~(P23iw6 & W23iw6));
assign W23iw6 = (D33iw6 & K33iw6);
assign K33iw6 = (R33iw6 & A62iw6);
assign R33iw6 = (O62iw6 & V62iw6);
assign D33iw6 = (O6cet6 & C72iw6);
assign P23iw6 = (Y33iw6 & F43iw6);
assign F43iw6 = (~(M43iw6 | L82iw6));
assign M43iw6 = (T43iw6 | Q72iw6);
assign Y33iw6 = (~(J72iw6 | S82iw6));
assign Acf8v6 = (~(Hcf8v6 & A53iw6));
assign A53iw6 = (~(Euget6 & H53iw6));
assign H53iw6 = (!Orget6);
assign Hcf8v6 = (~(O53iw6 & V53iw6));
assign V53iw6 = (Wdlov6 & Orget6);
assign Wdlov6 = (~(Iu4ov6 | C63iw6));
assign Tbf8v6 = (~(J63iw6 & Q63iw6));
assign Q63iw6 = (~(Njlov6 & Pa2iw6));
assign J63iw6 = (~(Bklov6 & Pvj7z6[3]));
assign Mbf8v6 = (~(X63iw6 & E73iw6));
assign E73iw6 = (~(Ad2iw6 & L73iw6));
assign X63iw6 = (~(Bklov6 & Rmget6));
assign Fbf8v6 = (Z73iw6 ? S73iw6 : Hkget6);
assign S73iw6 = (G83iw6 & N83iw6);
assign Yaf8v6 = (Z73iw6 ? X72iw6 : Dtj7z6[5]);
assign Raf8v6 = (Z73iw6 ? E82iw6 : Dtj7z6[4]);
assign Kaf8v6 = (Z73iw6 ? L82iw6 : Dtj7z6[3]);
assign Daf8v6 = (Z73iw6 ? S82iw6 : Dtj7z6[2]);
assign W9f8v6 = (~(U83iw6 & B93iw6));
assign B93iw6 = (~(Njlov6 & Kb2iw6));
assign U83iw6 = (~(Bklov6 & Pvj7z6[2]));
assign P9f8v6 = (~(I93iw6 & P93iw6));
assign P93iw6 = (~(Njlov6 & Fc2iw6));
assign Njlov6 = (L73iw6 & D42iw6);
assign L73iw6 = (O53iw6 & W93iw6);
assign W93iw6 = (~(Da3iw6 | Bklov6));
assign I93iw6 = (~(Bklov6 & Pvj7z6[1]));
assign Bklov6 = (!Z73iw6);
assign Z73iw6 = (~(Ka3iw6 & Ra3iw6));
assign Ra3iw6 = (~(O53iw6 & Ya3iw6));
assign Ya3iw6 = (~(Da3iw6 | MPUDISABLE));
assign O53iw6 = (G13iw6 & N13iw6);
assign Ka3iw6 = (~(Fb3iw6 & Mb3iw6));
assign Mb3iw6 = (~(Tb3iw6 & Ac3iw6));
assign Ac3iw6 = (~(Hc3iw6 | Rmget6));
assign Tb3iw6 = (Oc3iw6 & Vc3iw6);
assign Oc3iw6 = (~(Cd3iw6 & Jd3iw6));
assign Jd3iw6 = (Pvj7z6[1] | Pvj7z6[2]);
assign Fb3iw6 = (~(Pdlov6 | MPUDISABLE));
assign I9f8v6 = (Vd2iw6 ? Qd3iw6 : C1o7z6[1]);
assign Qd3iw6 = (M52iw6 & D42iw6);
assign B9f8v6 = (!Xd3iw6);
assign Xd3iw6 = (Pdlov6 ? Q497z6 : Ee3iw6);
assign U8f8v6 = (Vd2iw6 ? Le3iw6 : C1o7z6[0]);
assign Le3iw6 = (Se3iw6 & D42iw6);
assign N8f8v6 = (~(Ze3iw6 & Gf3iw6));
assign Gf3iw6 = (~(Lgj7z6[190] & Kw2iw6));
assign Ze3iw6 = (~(Nf3iw6 & Rw2iw6));
assign G8f8v6 = (~(Uf3iw6 & Bg3iw6));
assign Bg3iw6 = (~(Lgj7z6[178] & Iv2iw6));
assign Uf3iw6 = (~(Nf3iw6 & Pv2iw6));
assign Z7f8v6 = (~(Ig3iw6 & Pg3iw6));
assign Pg3iw6 = (~(Lgj7z6[166] & Gu2iw6));
assign Ig3iw6 = (~(Nf3iw6 & Nu2iw6));
assign S7f8v6 = (~(Wg3iw6 & Dh3iw6));
assign Dh3iw6 = (~(Lgj7z6[154] & Et2iw6));
assign Wg3iw6 = (~(Nf3iw6 & Lt2iw6));
assign L7f8v6 = (~(Kh3iw6 & Rh3iw6));
assign Rh3iw6 = (~(Lgj7z6[142] & Cs2iw6));
assign Kh3iw6 = (~(Nf3iw6 & Js2iw6));
assign E7f8v6 = (~(Yh3iw6 & Fi3iw6));
assign Fi3iw6 = (~(Lgj7z6[130] & Ar2iw6));
assign Yh3iw6 = (~(Nf3iw6 & Hr2iw6));
assign X6f8v6 = (~(Mi3iw6 & Ti3iw6));
assign Ti3iw6 = (~(Lgj7z6[118] & Yp2iw6));
assign Mi3iw6 = (~(Nf3iw6 & Fq2iw6));
assign Q6f8v6 = (~(Aj3iw6 & Hj3iw6));
assign Hj3iw6 = (~(Lgj7z6[106] & Wo2iw6));
assign Aj3iw6 = (~(Nf3iw6 & Dp2iw6));
assign J6f8v6 = (~(Oj3iw6 & Vj3iw6));
assign Vj3iw6 = (~(Lgj7z6[94] & Un2iw6));
assign Oj3iw6 = (~(Nf3iw6 & Bo2iw6));
assign C6f8v6 = (~(Ck3iw6 & Jk3iw6));
assign Jk3iw6 = (~(Lgj7z6[82] & Sm2iw6));
assign Ck3iw6 = (~(Nf3iw6 & Zm2iw6));
assign V5f8v6 = (~(Qk3iw6 & Xk3iw6));
assign Xk3iw6 = (~(Lgj7z6[70] & Ql2iw6));
assign Qk3iw6 = (~(Nf3iw6 & Xl2iw6));
assign O5f8v6 = (~(El3iw6 & Ll3iw6));
assign Ll3iw6 = (~(Lgj7z6[58] & Ok2iw6));
assign El3iw6 = (~(Nf3iw6 & Vk2iw6));
assign H5f8v6 = (~(Sl3iw6 & Zl3iw6));
assign Zl3iw6 = (~(Lgj7z6[46] & Mj2iw6));
assign Sl3iw6 = (~(Nf3iw6 & Tj2iw6));
assign A5f8v6 = (~(Gm3iw6 & Nm3iw6));
assign Nm3iw6 = (~(Lgj7z6[34] & Ki2iw6));
assign Gm3iw6 = (~(Nf3iw6 & Ri2iw6));
assign T4f8v6 = (~(Um3iw6 & Bn3iw6));
assign Bn3iw6 = (~(Lgj7z6[22] & Ih2iw6));
assign Um3iw6 = (~(Nf3iw6 & Ph2iw6));
assign M4f8v6 = (~(In3iw6 & Pn3iw6));
assign Pn3iw6 = (~(Lgj7z6[10] & Zf2iw6));
assign In3iw6 = (~(Nf3iw6 & Ng2iw6));
assign F4f8v6 = (~(Wn3iw6 & Do3iw6));
assign Do3iw6 = (~(Ohj7z6[30] & Ko3iw6));
assign Ko3iw6 = (~(Cz2iw6 & Ro3iw6));
assign Wn3iw6 = (~(Nf3iw6 & Jz2iw6));
assign Y3f8v6 = (~(Yo3iw6 & Fp3iw6));
assign Fp3iw6 = (~(Ohj7z6[62] & Mp3iw6));
assign Mp3iw6 = (~(Tx2iw6 & Ro3iw6));
assign Yo3iw6 = (~(Nf3iw6 & Ay2iw6));
assign R3f8v6 = (~(Tp3iw6 & Aq3iw6));
assign Aq3iw6 = (~(Lgj7z6[189] & Kw2iw6));
assign Kw2iw6 = (~(Rw2iw6 & Bqi7z6[3]));
assign Tp3iw6 = (~(Rw2iw6 & Hq3iw6));
assign K3f8v6 = (~(Oq3iw6 & Vq3iw6));
assign Vq3iw6 = (~(Lgj7z6[177] & Iv2iw6));
assign Iv2iw6 = (~(Pv2iw6 & Bqi7z6[3]));
assign Oq3iw6 = (~(Pv2iw6 & Hq3iw6));
assign D3f8v6 = (~(Cr3iw6 & Jr3iw6));
assign Jr3iw6 = (~(Lgj7z6[165] & Gu2iw6));
assign Gu2iw6 = (~(Nu2iw6 & Bqi7z6[3]));
assign Cr3iw6 = (~(Nu2iw6 & Hq3iw6));
assign W2f8v6 = (~(Qr3iw6 & Xr3iw6));
assign Xr3iw6 = (~(Lgj7z6[153] & Et2iw6));
assign Et2iw6 = (~(Lt2iw6 & Bqi7z6[3]));
assign Qr3iw6 = (~(Lt2iw6 & Hq3iw6));
assign P2f8v6 = (~(Es3iw6 & Ls3iw6));
assign Ls3iw6 = (~(Lgj7z6[141] & Cs2iw6));
assign Cs2iw6 = (~(Js2iw6 & Bqi7z6[3]));
assign Es3iw6 = (~(Js2iw6 & Hq3iw6));
assign I2f8v6 = (~(Ss3iw6 & Zs3iw6));
assign Zs3iw6 = (~(Lgj7z6[129] & Ar2iw6));
assign Ar2iw6 = (~(Hr2iw6 & Bqi7z6[3]));
assign Ss3iw6 = (~(Hr2iw6 & Hq3iw6));
assign B2f8v6 = (~(Gt3iw6 & Nt3iw6));
assign Nt3iw6 = (~(Lgj7z6[117] & Yp2iw6));
assign Yp2iw6 = (~(Fq2iw6 & Bqi7z6[3]));
assign Gt3iw6 = (~(Fq2iw6 & Hq3iw6));
assign U1f8v6 = (~(Ut3iw6 & Bu3iw6));
assign Bu3iw6 = (~(Lgj7z6[105] & Wo2iw6));
assign Wo2iw6 = (~(Dp2iw6 & Bqi7z6[3]));
assign Ut3iw6 = (~(Dp2iw6 & Hq3iw6));
assign N1f8v6 = (~(Iu3iw6 & Pu3iw6));
assign Pu3iw6 = (~(Lgj7z6[93] & Un2iw6));
assign Un2iw6 = (Wu3iw6 | Dv3iw6);
assign Iu3iw6 = (~(Bo2iw6 & Hq3iw6));
assign G1f8v6 = (~(Kv3iw6 & Rv3iw6));
assign Rv3iw6 = (~(Lgj7z6[81] & Sm2iw6));
assign Sm2iw6 = (~(Zm2iw6 & Bqi7z6[3]));
assign Kv3iw6 = (~(Zm2iw6 & Hq3iw6));
assign Z0f8v6 = (~(Yv3iw6 & Fw3iw6));
assign Fw3iw6 = (~(Lgj7z6[69] & Ql2iw6));
assign Ql2iw6 = (~(Xl2iw6 & Bqi7z6[3]));
assign Yv3iw6 = (~(Xl2iw6 & Hq3iw6));
assign S0f8v6 = (~(Mw3iw6 & Tw3iw6));
assign Tw3iw6 = (~(Lgj7z6[57] & Ok2iw6));
assign Ok2iw6 = (~(Vk2iw6 & Bqi7z6[3]));
assign Mw3iw6 = (~(Vk2iw6 & Hq3iw6));
assign L0f8v6 = (~(Ax3iw6 & Hx3iw6));
assign Hx3iw6 = (~(Lgj7z6[45] & Mj2iw6));
assign Mj2iw6 = (~(Tj2iw6 & Bqi7z6[3]));
assign Ax3iw6 = (~(Tj2iw6 & Hq3iw6));
assign E0f8v6 = (~(Ox3iw6 & Vx3iw6));
assign Vx3iw6 = (~(Lgj7z6[33] & Ki2iw6));
assign Ki2iw6 = (~(Ri2iw6 & Bqi7z6[3]));
assign Ox3iw6 = (~(Ri2iw6 & Hq3iw6));
assign Xze8v6 = (~(Cy3iw6 & Jy3iw6));
assign Jy3iw6 = (~(Lgj7z6[21] & Ih2iw6));
assign Ih2iw6 = (~(Ph2iw6 & Bqi7z6[3]));
assign Cy3iw6 = (~(Ph2iw6 & Hq3iw6));
assign Qze8v6 = (~(Qy3iw6 & Xy3iw6));
assign Xy3iw6 = (~(Lgj7z6[9] & Zf2iw6));
assign Zf2iw6 = (~(Ng2iw6 & Bqi7z6[3]));
assign Qy3iw6 = (~(Ng2iw6 & Hq3iw6));
assign Jze8v6 = (~(Ez3iw6 & Lz3iw6));
assign Lz3iw6 = (~(Ohj7z6[29] & Sz3iw6));
assign Sz3iw6 = (~(Cz2iw6 & Zz3iw6));
assign Ez3iw6 = (~(Jz2iw6 & Hq3iw6));
assign Cze8v6 = (~(G04iw6 & N04iw6));
assign N04iw6 = (~(Ohj7z6[61] & U04iw6));
assign U04iw6 = (~(Tx2iw6 & Zz3iw6));
assign G04iw6 = (~(Ay2iw6 & Hq3iw6));
assign Vye8v6 = (~(B14iw6 & I14iw6));
assign I14iw6 = (~(Ohj7z6[28] & P14iw6));
assign P14iw6 = (~(Cz2iw6 & W14iw6));
assign B14iw6 = (~(D24iw6 & W14iw6));
assign Oye8v6 = (~(K24iw6 & R24iw6));
assign R24iw6 = (~(Ohj7z6[60] & Y24iw6));
assign Y24iw6 = (~(Tx2iw6 & W14iw6));
assign K24iw6 = (~(F34iw6 & W14iw6));
assign Hye8v6 = (~(M34iw6 & T34iw6));
assign T34iw6 = (~(Ohj7z6[27] & A44iw6));
assign A44iw6 = (~(Cz2iw6 & H44iw6));
assign M34iw6 = (~(D24iw6 & H44iw6));
assign Aye8v6 = (~(O44iw6 & V44iw6));
assign V44iw6 = (~(Ohj7z6[59] & C54iw6));
assign C54iw6 = (~(Tx2iw6 & H44iw6));
assign O44iw6 = (~(F34iw6 & H44iw6));
assign Txe8v6 = (~(J54iw6 & Q54iw6));
assign Q54iw6 = (~(Ohj7z6[26] & X54iw6));
assign X54iw6 = (~(Cz2iw6 & E64iw6));
assign J54iw6 = (~(D24iw6 & E64iw6));
assign Mxe8v6 = (~(L64iw6 & S64iw6));
assign S64iw6 = (~(Ohj7z6[58] & Z64iw6));
assign Z64iw6 = (~(Tx2iw6 & E64iw6));
assign L64iw6 = (~(F34iw6 & E64iw6));
assign Fxe8v6 = (~(G74iw6 & N74iw6));
assign N74iw6 = (~(Ohj7z6[25] & U74iw6));
assign U74iw6 = (~(Cz2iw6 & Iklov6));
assign G74iw6 = (~(D24iw6 & Iklov6));
assign Ywe8v6 = (~(B84iw6 & I84iw6));
assign I84iw6 = (~(Ohj7z6[57] & P84iw6));
assign P84iw6 = (~(Tx2iw6 & Iklov6));
assign B84iw6 = (~(F34iw6 & Iklov6));
assign Rwe8v6 = (!W84iw6);
assign W84iw6 = (K94iw6 ? Pfh7v6 : D94iw6);
assign Kwe8v6 = (!R94iw6);
assign R94iw6 = (K94iw6 ? Cjh7v6 : Y94iw6);
assign Dwe8v6 = (K94iw6 ? HTMDHPROT[1] : Hjqnv6);
assign Wve8v6 = (K94iw6 ? Fa4iw6 : Anehw6);
assign Pve8v6 = (!Ma4iw6);
assign Ma4iw6 = (K94iw6 ? Kgh7v6 : Ta4iw6);
assign Ive8v6 = (!Ab4iw6);
assign Ab4iw6 = (Ob4iw6 ? Hb4iw6 : Dgh7v6);
assign Hb4iw6 = (~(Aeonv6 & Vb4iw6));
assign Bve8v6 = (K94iw6 ? HTMDHTRANS[0] : Cc4iw6);
assign Cc4iw6 = (Jc4iw6 & Aeonv6);
assign Uue8v6 = (K94iw6 ? HTMDHADDR[31] : Cmm7z6[31]);
assign Nue8v6 = (K94iw6 ? HTMDHADDR[30] : Cmm7z6[30]);
assign Gue8v6 = (K94iw6 ? HTMDHADDR[29] : Cmm7z6[29]);
assign Zte8v6 = (K94iw6 ? HTMDHADDR[28] : Cmm7z6[28]);
assign Ste8v6 = (K94iw6 ? HTMDHADDR[27] : Cmm7z6[27]);
assign Lte8v6 = (K94iw6 ? HTMDHADDR[26] : Cmm7z6[26]);
assign Ete8v6 = (K94iw6 ? HTMDHADDR[25] : Cmm7z6[25]);
assign Xse8v6 = (K94iw6 ? HTMDHADDR[24] : Cmm7z6[24]);
assign Qse8v6 = (K94iw6 ? HTMDHADDR[23] : Cmm7z6[23]);
assign Jse8v6 = (K94iw6 ? HTMDHADDR[22] : Cmm7z6[22]);
assign Cse8v6 = (K94iw6 ? HTMDHADDR[21] : Cmm7z6[21]);
assign Vre8v6 = (K94iw6 ? HTMDHADDR[20] : Cmm7z6[20]);
assign Ore8v6 = (K94iw6 ? HTMDHADDR[19] : Cmm7z6[19]);
assign Hre8v6 = (K94iw6 ? HTMDHADDR[18] : Cmm7z6[18]);
assign Are8v6 = (K94iw6 ? HTMDHADDR[17] : Cmm7z6[17]);
assign Tqe8v6 = (K94iw6 ? HTMDHADDR[16] : Cmm7z6[16]);
assign Mqe8v6 = (K94iw6 ? HTMDHADDR[15] : Cmm7z6[15]);
assign Fqe8v6 = (K94iw6 ? HTMDHADDR[14] : Cmm7z6[14]);
assign Ype8v6 = (K94iw6 ? HTMDHADDR[13] : Cmm7z6[13]);
assign Rpe8v6 = (K94iw6 ? HTMDHADDR[12] : Cmm7z6[12]);
assign Kpe8v6 = (K94iw6 ? HTMDHADDR[11] : Cmm7z6[11]);
assign Dpe8v6 = (K94iw6 ? HTMDHADDR[10] : Cmm7z6[10]);
assign Woe8v6 = (K94iw6 ? HTMDHADDR[9] : Cmm7z6[9]);
assign Poe8v6 = (K94iw6 ? HTMDHADDR[8] : Cmm7z6[8]);
assign Ioe8v6 = (K94iw6 ? HTMDHADDR[7] : Cmm7z6[7]);
assign Boe8v6 = (K94iw6 ? HTMDHADDR[6] : Cmm7z6[6]);
assign Une8v6 = (K94iw6 ? HTMDHADDR[5] : Cmm7z6[5]);
assign Nne8v6 = (K94iw6 ? HTMDHADDR[4] : Cmm7z6[4]);
assign Gne8v6 = (K94iw6 ? HTMDHADDR[3] : Cmm7z6[3]);
assign Zme8v6 = (K94iw6 ? HTMDHADDR[2] : Yefnv6);
assign Sme8v6 = (!Qc4iw6);
assign Qc4iw6 = (K94iw6 ? Rgh7v6 : Xc4iw6);
assign Lme8v6 = (!Ed4iw6);
assign Ed4iw6 = (Ob4iw6 ? Sd4iw6 : Ld4iw6);
assign Sd4iw6 = (~(Zd4iw6 & Ge4iw6));
assign Ge4iw6 = (~(Kgh7v6 & Wfh7v6));
assign Zd4iw6 = (~(Pfh7v6 | Dgh7v6));
assign Eme8v6 = (!Ne4iw6);
assign Ne4iw6 = (Ob4iw6 ? Bf4iw6 : Ue4iw6);
assign Bf4iw6 = (~(If4iw6 & Pf4iw6));
assign Pf4iw6 = (~(Dgh7v6 | Rgh7v6));
assign If4iw6 = (Kgh7v6 & Fa4iw6);
assign Fa4iw6 = (!Wfh7v6);
assign Qle8v6 = (Dg4iw6 ? Wf4iw6 : Dri7z6[24]);
assign Jle8v6 = (Dg4iw6 ? Iklov6 : Dri7z6[25]);
assign Cle8v6 = (Dg4iw6 ? E64iw6 : Dri7z6[26]);
assign Vke8v6 = (Dg4iw6 ? H44iw6 : Dri7z6[27]);
assign Oke8v6 = (Dg4iw6 ? W14iw6 : Dri7z6[28]);
assign Hke8v6 = (Dg4iw6 ? Zz3iw6 : Dri7z6[29]);
assign Ake8v6 = (Dg4iw6 ? Ro3iw6 : Dri7z6[30]);
assign Tje8v6 = (Dg4iw6 ? X0hov6 : Dri7z6[31]);
assign Dg4iw6 = (~(Kg4iw6 | Dv3iw6));
assign Mje8v6 = (~(Rg4iw6 & Yg4iw6));
assign Yg4iw6 = (~(Ohj7z6[24] & Fh4iw6));
assign Fh4iw6 = (~(Cz2iw6 & Wf4iw6));
assign Cz2iw6 = (~(Mh4iw6 | Dv3iw6));
assign Rg4iw6 = (~(D24iw6 & Wf4iw6));
assign D24iw6 = (Jz2iw6 & Bqi7z6[3]);
assign Fje8v6 = (~(Th4iw6 & Ai4iw6));
assign Ai4iw6 = (~(Ohj7z6[56] & Hi4iw6));
assign Hi4iw6 = (~(Tx2iw6 & Wf4iw6));
assign Tx2iw6 = (~(Oi4iw6 | Dv3iw6));
assign Th4iw6 = (~(F34iw6 & Wf4iw6));
assign F34iw6 = (Ay2iw6 & Bqi7z6[3]);
assign Yie8v6 = (~(Vi4iw6 & Cj4iw6));
assign Cj4iw6 = (~(Lgj7z6[188] & Jj4iw6));
assign Vi4iw6 = (~(Qj4iw6 & Rw2iw6));
assign Rie8v6 = (~(Xj4iw6 & Ek4iw6));
assign Ek4iw6 = (~(Lgj7z6[176] & Lk4iw6));
assign Xj4iw6 = (~(Qj4iw6 & Pv2iw6));
assign Kie8v6 = (~(Sk4iw6 & Zk4iw6));
assign Zk4iw6 = (~(Lgj7z6[164] & Gl4iw6));
assign Sk4iw6 = (~(Qj4iw6 & Nu2iw6));
assign Die8v6 = (~(Nl4iw6 & Ul4iw6));
assign Ul4iw6 = (~(Lgj7z6[152] & Bm4iw6));
assign Nl4iw6 = (~(Qj4iw6 & Lt2iw6));
assign Whe8v6 = (~(Im4iw6 & Pm4iw6));
assign Pm4iw6 = (~(Lgj7z6[140] & Wm4iw6));
assign Im4iw6 = (~(Qj4iw6 & Js2iw6));
assign Phe8v6 = (~(Dn4iw6 & Kn4iw6));
assign Kn4iw6 = (~(Lgj7z6[128] & Rn4iw6));
assign Dn4iw6 = (~(Qj4iw6 & Hr2iw6));
assign Ihe8v6 = (~(Yn4iw6 & Fo4iw6));
assign Fo4iw6 = (~(Lgj7z6[116] & Mo4iw6));
assign Yn4iw6 = (~(Qj4iw6 & Fq2iw6));
assign Bhe8v6 = (~(To4iw6 & Ap4iw6));
assign Ap4iw6 = (~(Lgj7z6[104] & Hp4iw6));
assign To4iw6 = (~(Qj4iw6 & Dp2iw6));
assign Uge8v6 = (~(Op4iw6 & Vp4iw6));
assign Vp4iw6 = (~(Lgj7z6[92] & Cq4iw6));
assign Op4iw6 = (~(Qj4iw6 & Bo2iw6));
assign Nge8v6 = (~(Jq4iw6 & Qq4iw6));
assign Qq4iw6 = (~(Lgj7z6[80] & Xq4iw6));
assign Jq4iw6 = (~(Qj4iw6 & Zm2iw6));
assign Gge8v6 = (~(Er4iw6 & Lr4iw6));
assign Lr4iw6 = (~(Lgj7z6[68] & Sr4iw6));
assign Er4iw6 = (~(Qj4iw6 & Xl2iw6));
assign Zfe8v6 = (~(Zr4iw6 & Gs4iw6));
assign Gs4iw6 = (~(Lgj7z6[56] & Ns4iw6));
assign Zr4iw6 = (~(Qj4iw6 & Vk2iw6));
assign Sfe8v6 = (~(Us4iw6 & Bt4iw6));
assign Bt4iw6 = (~(Lgj7z6[44] & It4iw6));
assign Us4iw6 = (~(Qj4iw6 & Tj2iw6));
assign Lfe8v6 = (~(Pt4iw6 & Wt4iw6));
assign Wt4iw6 = (~(Lgj7z6[32] & Du4iw6));
assign Pt4iw6 = (~(Qj4iw6 & Ri2iw6));
assign Efe8v6 = (~(Ku4iw6 & Ru4iw6));
assign Ru4iw6 = (~(Lgj7z6[20] & Yu4iw6));
assign Ku4iw6 = (~(Qj4iw6 & Ph2iw6));
assign Xee8v6 = (~(Fv4iw6 & Mv4iw6));
assign Mv4iw6 = (~(Lgj7z6[8] & Tv4iw6));
assign Fv4iw6 = (~(Qj4iw6 & Ng2iw6));
assign Qee8v6 = (~(Aw4iw6 & Hw4iw6));
assign Hw4iw6 = (~(Ohj7z6[23] & Ow4iw6));
assign Ow4iw6 = (~(Vw4iw6 & Cx4iw6));
assign Aw4iw6 = (~(Qj4iw6 & Jz2iw6));
assign Jee8v6 = (~(Jx4iw6 & Qx4iw6));
assign Qx4iw6 = (~(Ohj7z6[55] & Xx4iw6));
assign Xx4iw6 = (~(Ey4iw6 & Cx4iw6));
assign Jx4iw6 = (~(Qj4iw6 & Ay2iw6));
assign Cee8v6 = (~(Ly4iw6 & Sy4iw6));
assign Sy4iw6 = (~(Lgj7z6[187] & Jj4iw6));
assign Ly4iw6 = (~(Rw2iw6 & Zy4iw6));
assign Vde8v6 = (~(Gz4iw6 & Nz4iw6));
assign Nz4iw6 = (~(Lgj7z6[175] & Lk4iw6));
assign Gz4iw6 = (~(Pv2iw6 & Zy4iw6));
assign Ode8v6 = (~(Uz4iw6 & B05iw6));
assign B05iw6 = (~(Lgj7z6[163] & Gl4iw6));
assign Uz4iw6 = (~(Nu2iw6 & Zy4iw6));
assign Hde8v6 = (~(I05iw6 & P05iw6));
assign P05iw6 = (~(Lgj7z6[151] & Bm4iw6));
assign I05iw6 = (~(Lt2iw6 & Zy4iw6));
assign Ade8v6 = (~(W05iw6 & D15iw6));
assign D15iw6 = (~(Lgj7z6[139] & Wm4iw6));
assign W05iw6 = (~(Js2iw6 & Zy4iw6));
assign Tce8v6 = (~(K15iw6 & R15iw6));
assign R15iw6 = (~(Lgj7z6[127] & Rn4iw6));
assign K15iw6 = (~(Hr2iw6 & Zy4iw6));
assign Mce8v6 = (~(Y15iw6 & F25iw6));
assign F25iw6 = (~(Lgj7z6[115] & Mo4iw6));
assign Y15iw6 = (~(Fq2iw6 & Zy4iw6));
assign Fce8v6 = (~(M25iw6 & T25iw6));
assign T25iw6 = (~(Lgj7z6[103] & Hp4iw6));
assign M25iw6 = (~(Dp2iw6 & Zy4iw6));
assign Ybe8v6 = (~(A35iw6 & H35iw6));
assign H35iw6 = (~(Lgj7z6[91] & Cq4iw6));
assign A35iw6 = (~(Bo2iw6 & Zy4iw6));
assign Rbe8v6 = (~(O35iw6 & V35iw6));
assign V35iw6 = (~(Lgj7z6[79] & Xq4iw6));
assign O35iw6 = (~(Zm2iw6 & Zy4iw6));
assign Kbe8v6 = (~(C45iw6 & J45iw6));
assign J45iw6 = (~(Lgj7z6[67] & Sr4iw6));
assign C45iw6 = (~(Xl2iw6 & Zy4iw6));
assign Dbe8v6 = (~(Q45iw6 & X45iw6));
assign X45iw6 = (~(Lgj7z6[55] & Ns4iw6));
assign Q45iw6 = (~(Vk2iw6 & Zy4iw6));
assign Wae8v6 = (~(E55iw6 & L55iw6));
assign L55iw6 = (~(Lgj7z6[43] & It4iw6));
assign E55iw6 = (~(Tj2iw6 & Zy4iw6));
assign Pae8v6 = (~(S55iw6 & Z55iw6));
assign Z55iw6 = (~(Lgj7z6[31] & Du4iw6));
assign S55iw6 = (~(Ri2iw6 & Zy4iw6));
assign Iae8v6 = (~(G65iw6 & N65iw6));
assign N65iw6 = (~(Lgj7z6[19] & Yu4iw6));
assign G65iw6 = (~(Ph2iw6 & Zy4iw6));
assign Bae8v6 = (~(U65iw6 & B75iw6));
assign B75iw6 = (~(Lgj7z6[7] & Tv4iw6));
assign U65iw6 = (~(Ng2iw6 & Zy4iw6));
assign U9e8v6 = (~(I75iw6 & P75iw6));
assign P75iw6 = (~(Ohj7z6[22] & W75iw6));
assign W75iw6 = (~(Vw4iw6 & D85iw6));
assign I75iw6 = (~(Jz2iw6 & Zy4iw6));
assign N9e8v6 = (~(K85iw6 & R85iw6));
assign R85iw6 = (~(Ohj7z6[54] & Y85iw6));
assign Y85iw6 = (~(Ey4iw6 & D85iw6));
assign K85iw6 = (~(Ay2iw6 & Zy4iw6));
assign G9e8v6 = (~(F95iw6 & M95iw6));
assign M95iw6 = (~(Lgj7z6[186] & Jj4iw6));
assign Jj4iw6 = (~(Rw2iw6 & Bqi7z6[2]));
assign F95iw6 = (~(T95iw6 & Rw2iw6));
assign Z8e8v6 = (~(Aa5iw6 & Ha5iw6));
assign Ha5iw6 = (~(Lgj7z6[174] & Lk4iw6));
assign Lk4iw6 = (~(Pv2iw6 & Bqi7z6[2]));
assign Aa5iw6 = (~(T95iw6 & Pv2iw6));
assign S8e8v6 = (~(Oa5iw6 & Va5iw6));
assign Va5iw6 = (~(Lgj7z6[162] & Gl4iw6));
assign Gl4iw6 = (~(Nu2iw6 & Bqi7z6[2]));
assign Oa5iw6 = (~(T95iw6 & Nu2iw6));
assign L8e8v6 = (~(Cb5iw6 & Jb5iw6));
assign Jb5iw6 = (~(Lgj7z6[150] & Bm4iw6));
assign Bm4iw6 = (~(Lt2iw6 & Bqi7z6[2]));
assign Cb5iw6 = (~(T95iw6 & Lt2iw6));
assign E8e8v6 = (~(Qb5iw6 & Xb5iw6));
assign Xb5iw6 = (~(Lgj7z6[138] & Wm4iw6));
assign Wm4iw6 = (~(Js2iw6 & Bqi7z6[2]));
assign Qb5iw6 = (~(T95iw6 & Js2iw6));
assign X7e8v6 = (~(Ec5iw6 & Lc5iw6));
assign Lc5iw6 = (~(Lgj7z6[126] & Rn4iw6));
assign Rn4iw6 = (~(Hr2iw6 & Bqi7z6[2]));
assign Ec5iw6 = (~(T95iw6 & Hr2iw6));
assign Q7e8v6 = (~(Sc5iw6 & Zc5iw6));
assign Zc5iw6 = (~(Lgj7z6[114] & Mo4iw6));
assign Mo4iw6 = (~(Fq2iw6 & Bqi7z6[2]));
assign Sc5iw6 = (~(T95iw6 & Fq2iw6));
assign J7e8v6 = (~(Gd5iw6 & Nd5iw6));
assign Nd5iw6 = (~(Lgj7z6[102] & Hp4iw6));
assign Hp4iw6 = (~(Dp2iw6 & Bqi7z6[2]));
assign Gd5iw6 = (~(T95iw6 & Dp2iw6));
assign C7e8v6 = (~(Ud5iw6 & Be5iw6));
assign Be5iw6 = (~(Lgj7z6[90] & Cq4iw6));
assign Cq4iw6 = (Wu3iw6 | Ie5iw6);
assign Ud5iw6 = (~(T95iw6 & Bo2iw6));
assign V6e8v6 = (~(Pe5iw6 & We5iw6));
assign We5iw6 = (~(Lgj7z6[78] & Xq4iw6));
assign Xq4iw6 = (~(Zm2iw6 & Bqi7z6[2]));
assign Pe5iw6 = (~(T95iw6 & Zm2iw6));
assign O6e8v6 = (~(Df5iw6 & Kf5iw6));
assign Kf5iw6 = (~(Lgj7z6[66] & Sr4iw6));
assign Sr4iw6 = (~(Xl2iw6 & Bqi7z6[2]));
assign Df5iw6 = (~(T95iw6 & Xl2iw6));
assign H6e8v6 = (~(Rf5iw6 & Yf5iw6));
assign Yf5iw6 = (~(Lgj7z6[54] & Ns4iw6));
assign Ns4iw6 = (~(Vk2iw6 & Bqi7z6[2]));
assign Rf5iw6 = (~(T95iw6 & Vk2iw6));
assign A6e8v6 = (~(Fg5iw6 & Mg5iw6));
assign Mg5iw6 = (~(Lgj7z6[42] & It4iw6));
assign It4iw6 = (~(Tj2iw6 & Bqi7z6[2]));
assign Fg5iw6 = (~(T95iw6 & Tj2iw6));
assign T5e8v6 = (~(Tg5iw6 & Ah5iw6));
assign Ah5iw6 = (~(Lgj7z6[30] & Du4iw6));
assign Du4iw6 = (~(Ri2iw6 & Bqi7z6[2]));
assign Tg5iw6 = (~(T95iw6 & Ri2iw6));
assign M5e8v6 = (~(Hh5iw6 & Oh5iw6));
assign Oh5iw6 = (~(Lgj7z6[18] & Yu4iw6));
assign Yu4iw6 = (~(Ph2iw6 & Bqi7z6[2]));
assign Hh5iw6 = (~(T95iw6 & Ph2iw6));
assign F5e8v6 = (~(Vh5iw6 & Ci5iw6));
assign Ci5iw6 = (~(Lgj7z6[6] & Tv4iw6));
assign Tv4iw6 = (~(Ng2iw6 & Bqi7z6[2]));
assign Vh5iw6 = (~(T95iw6 & Ng2iw6));
assign Y4e8v6 = (~(Ji5iw6 & Qi5iw6));
assign Qi5iw6 = (~(Ohj7z6[21] & Xi5iw6));
assign Xi5iw6 = (~(Vw4iw6 & Ej5iw6));
assign Ji5iw6 = (~(T95iw6 & Jz2iw6));
assign R4e8v6 = (~(Lj5iw6 & Sj5iw6));
assign Sj5iw6 = (~(Ohj7z6[53] & Zj5iw6));
assign Zj5iw6 = (~(Ey4iw6 & Ej5iw6));
assign Lj5iw6 = (~(T95iw6 & Ay2iw6));
assign K4e8v6 = (~(Gk5iw6 & Nk5iw6));
assign Nk5iw6 = (~(Ohj7z6[20] & Uk5iw6));
assign Uk5iw6 = (~(Vw4iw6 & Bl5iw6));
assign Gk5iw6 = (~(Il5iw6 & Bl5iw6));
assign D4e8v6 = (~(Pl5iw6 & Wl5iw6));
assign Wl5iw6 = (~(Ohj7z6[52] & Dm5iw6));
assign Dm5iw6 = (~(Ey4iw6 & Bl5iw6));
assign Pl5iw6 = (~(Km5iw6 & Bl5iw6));
assign W3e8v6 = (~(Rm5iw6 & Ym5iw6));
assign Ym5iw6 = (~(Ohj7z6[19] & Fn5iw6));
assign Fn5iw6 = (~(Vw4iw6 & Mn5iw6));
assign Rm5iw6 = (~(Il5iw6 & Mn5iw6));
assign P3e8v6 = (~(Tn5iw6 & Ao5iw6));
assign Ao5iw6 = (~(Ohj7z6[51] & Ho5iw6));
assign Ho5iw6 = (~(Ey4iw6 & Mn5iw6));
assign Tn5iw6 = (~(Km5iw6 & Mn5iw6));
assign I3e8v6 = (~(Oo5iw6 & Vo5iw6));
assign Vo5iw6 = (~(Ohj7z6[18] & Cp5iw6));
assign Cp5iw6 = (~(Vw4iw6 & Jp5iw6));
assign Oo5iw6 = (~(Il5iw6 & Jp5iw6));
assign B3e8v6 = (~(Qp5iw6 & Xp5iw6));
assign Xp5iw6 = (~(Ohj7z6[50] & Eq5iw6));
assign Eq5iw6 = (~(Ey4iw6 & Jp5iw6));
assign Qp5iw6 = (~(Km5iw6 & Jp5iw6));
assign U2e8v6 = (~(Lq5iw6 & Sq5iw6));
assign Sq5iw6 = (~(Ohj7z6[17] & Zq5iw6));
assign Zq5iw6 = (~(Vw4iw6 & Gr5iw6));
assign Lq5iw6 = (~(Il5iw6 & Gr5iw6));
assign N2e8v6 = (~(Nr5iw6 & Ur5iw6));
assign Ur5iw6 = (~(Ohj7z6[49] & Bs5iw6));
assign Bs5iw6 = (~(Ey4iw6 & Gr5iw6));
assign Nr5iw6 = (~(Km5iw6 & Gr5iw6));
assign G2e8v6 = (Ps5iw6 ? Is5iw6 : Dri7z6[16]);
assign Z1e8v6 = (Ps5iw6 ? Gr5iw6 : Dri7z6[17]);
assign S1e8v6 = (Ps5iw6 ? Jp5iw6 : Dri7z6[18]);
assign L1e8v6 = (Ps5iw6 ? Mn5iw6 : Dri7z6[19]);
assign E1e8v6 = (Ps5iw6 ? Bl5iw6 : Dri7z6[20]);
assign X0e8v6 = (Ps5iw6 ? Ej5iw6 : Dri7z6[21]);
assign Q0e8v6 = (Ps5iw6 ? D85iw6 : Dri7z6[22]);
assign J0e8v6 = (Ps5iw6 ? Cx4iw6 : Dri7z6[23]);
assign Ps5iw6 = (~(Kg4iw6 | Ie5iw6));
assign C0e8v6 = (~(Ws5iw6 & Dt5iw6));
assign Dt5iw6 = (~(Ohj7z6[16] & Kt5iw6));
assign Kt5iw6 = (~(Vw4iw6 & Is5iw6));
assign Vw4iw6 = (~(Mh4iw6 | Ie5iw6));
assign Ws5iw6 = (~(Il5iw6 & Is5iw6));
assign Il5iw6 = (Jz2iw6 & Bqi7z6[2]);
assign Vzd8v6 = (~(Rt5iw6 & Yt5iw6));
assign Yt5iw6 = (~(Ohj7z6[48] & Fu5iw6));
assign Fu5iw6 = (~(Ey4iw6 & Is5iw6));
assign Ey4iw6 = (~(Oi4iw6 | Ie5iw6));
assign Rt5iw6 = (~(Km5iw6 & Is5iw6));
assign Km5iw6 = (Ay2iw6 & Bqi7z6[2]);
assign Ozd8v6 = (~(Mu5iw6 & Tu5iw6));
assign Tu5iw6 = (~(Lgj7z6[185] & Av5iw6));
assign Mu5iw6 = (~(Hv5iw6 & Rw2iw6));
assign Hzd8v6 = (~(Ov5iw6 & Vv5iw6));
assign Vv5iw6 = (~(Lgj7z6[173] & Cw5iw6));
assign Ov5iw6 = (~(Hv5iw6 & Pv2iw6));
assign Azd8v6 = (~(Jw5iw6 & Qw5iw6));
assign Qw5iw6 = (~(Lgj7z6[161] & Xw5iw6));
assign Jw5iw6 = (~(Hv5iw6 & Nu2iw6));
assign Tyd8v6 = (~(Ex5iw6 & Lx5iw6));
assign Lx5iw6 = (~(Lgj7z6[149] & Sx5iw6));
assign Ex5iw6 = (~(Hv5iw6 & Lt2iw6));
assign Myd8v6 = (~(Zx5iw6 & Gy5iw6));
assign Gy5iw6 = (~(Lgj7z6[137] & Ny5iw6));
assign Zx5iw6 = (~(Hv5iw6 & Js2iw6));
assign Fyd8v6 = (~(Uy5iw6 & Bz5iw6));
assign Bz5iw6 = (~(Lgj7z6[125] & Iz5iw6));
assign Uy5iw6 = (~(Hv5iw6 & Hr2iw6));
assign Yxd8v6 = (~(Pz5iw6 & Wz5iw6));
assign Wz5iw6 = (~(Lgj7z6[113] & D06iw6));
assign Pz5iw6 = (~(Hv5iw6 & Fq2iw6));
assign Rxd8v6 = (~(K06iw6 & R06iw6));
assign R06iw6 = (~(Lgj7z6[101] & Y06iw6));
assign K06iw6 = (~(Hv5iw6 & Dp2iw6));
assign Kxd8v6 = (~(F16iw6 & M16iw6));
assign M16iw6 = (T16iw6 | A26iw6);
assign F16iw6 = (~(Hv5iw6 & Bo2iw6));
assign Dxd8v6 = (~(H26iw6 & O26iw6));
assign O26iw6 = (~(Lgj7z6[77] & V26iw6));
assign H26iw6 = (~(Hv5iw6 & Zm2iw6));
assign Wwd8v6 = (~(C36iw6 & J36iw6));
assign J36iw6 = (~(Lgj7z6[65] & Q36iw6));
assign C36iw6 = (~(Hv5iw6 & Xl2iw6));
assign Pwd8v6 = (~(X36iw6 & E46iw6));
assign E46iw6 = (~(Lgj7z6[53] & L46iw6));
assign X36iw6 = (~(Hv5iw6 & Vk2iw6));
assign Iwd8v6 = (~(S46iw6 & Z46iw6));
assign Z46iw6 = (~(Lgj7z6[41] & G56iw6));
assign S46iw6 = (~(Hv5iw6 & Tj2iw6));
assign Bwd8v6 = (~(N56iw6 & U56iw6));
assign U56iw6 = (~(Lgj7z6[29] & B66iw6));
assign N56iw6 = (~(Hv5iw6 & Ri2iw6));
assign Uvd8v6 = (~(I66iw6 & P66iw6));
assign P66iw6 = (~(Lgj7z6[17] & W66iw6));
assign I66iw6 = (~(Hv5iw6 & Ph2iw6));
assign Nvd8v6 = (~(D76iw6 & K76iw6));
assign K76iw6 = (~(Lgj7z6[5] & R76iw6));
assign D76iw6 = (~(Hv5iw6 & Ng2iw6));
assign Gvd8v6 = (~(Y76iw6 & F86iw6));
assign F86iw6 = (~(Ohj7z6[15] & M86iw6));
assign M86iw6 = (~(T86iw6 & Z0iov6));
assign Y76iw6 = (~(Hv5iw6 & Jz2iw6));
assign Zud8v6 = (~(A96iw6 & H96iw6));
assign H96iw6 = (~(Ohj7z6[47] & O96iw6));
assign O96iw6 = (~(V96iw6 & Z0iov6));
assign A96iw6 = (~(Hv5iw6 & Ay2iw6));
assign Sud8v6 = (~(Ca6iw6 & Ja6iw6));
assign Ja6iw6 = (~(Lgj7z6[184] & Av5iw6));
assign Ca6iw6 = (~(Qa6iw6 & Rw2iw6));
assign Lud8v6 = (~(Xa6iw6 & Eb6iw6));
assign Eb6iw6 = (~(Lgj7z6[172] & Cw5iw6));
assign Xa6iw6 = (~(Qa6iw6 & Pv2iw6));
assign Eud8v6 = (~(Lb6iw6 & Sb6iw6));
assign Sb6iw6 = (~(Lgj7z6[160] & Xw5iw6));
assign Lb6iw6 = (~(Qa6iw6 & Nu2iw6));
assign Xtd8v6 = (~(Zb6iw6 & Gc6iw6));
assign Gc6iw6 = (~(Lgj7z6[148] & Sx5iw6));
assign Zb6iw6 = (~(Qa6iw6 & Lt2iw6));
assign Qtd8v6 = (~(Nc6iw6 & Uc6iw6));
assign Uc6iw6 = (~(Lgj7z6[136] & Ny5iw6));
assign Nc6iw6 = (~(Qa6iw6 & Js2iw6));
assign Jtd8v6 = (~(Bd6iw6 & Id6iw6));
assign Id6iw6 = (~(Lgj7z6[124] & Iz5iw6));
assign Bd6iw6 = (~(Qa6iw6 & Hr2iw6));
assign Ctd8v6 = (~(Pd6iw6 & Wd6iw6));
assign Wd6iw6 = (~(Lgj7z6[112] & D06iw6));
assign Pd6iw6 = (~(Qa6iw6 & Fq2iw6));
assign Vsd8v6 = (~(De6iw6 & Ke6iw6));
assign Ke6iw6 = (~(Lgj7z6[100] & Y06iw6));
assign De6iw6 = (~(Qa6iw6 & Dp2iw6));
assign Osd8v6 = (~(Re6iw6 & Ye6iw6));
assign Ye6iw6 = (Ff6iw6 | A26iw6);
assign Re6iw6 = (~(Qa6iw6 & Bo2iw6));
assign Hsd8v6 = (~(Mf6iw6 & Tf6iw6));
assign Tf6iw6 = (~(Lgj7z6[76] & V26iw6));
assign Mf6iw6 = (~(Qa6iw6 & Zm2iw6));
assign Asd8v6 = (~(Ag6iw6 & Hg6iw6));
assign Hg6iw6 = (~(Lgj7z6[64] & Q36iw6));
assign Ag6iw6 = (~(Qa6iw6 & Xl2iw6));
assign Trd8v6 = (~(Og6iw6 & Vg6iw6));
assign Vg6iw6 = (~(Lgj7z6[52] & L46iw6));
assign Og6iw6 = (~(Qa6iw6 & Vk2iw6));
assign Mrd8v6 = (~(Ch6iw6 & Jh6iw6));
assign Jh6iw6 = (~(Lgj7z6[40] & G56iw6));
assign Ch6iw6 = (~(Qa6iw6 & Tj2iw6));
assign Frd8v6 = (~(Qh6iw6 & Xh6iw6));
assign Xh6iw6 = (~(Lgj7z6[28] & B66iw6));
assign Qh6iw6 = (~(Qa6iw6 & Ri2iw6));
assign Yqd8v6 = (~(Ei6iw6 & Li6iw6));
assign Li6iw6 = (~(Lgj7z6[16] & W66iw6));
assign Ei6iw6 = (~(Qa6iw6 & Ph2iw6));
assign Rqd8v6 = (~(Si6iw6 & Zi6iw6));
assign Zi6iw6 = (~(Lgj7z6[4] & R76iw6));
assign Si6iw6 = (~(Qa6iw6 & Ng2iw6));
assign Kqd8v6 = (~(Gj6iw6 & Nj6iw6));
assign Nj6iw6 = (~(Ohj7z6[14] & Uj6iw6));
assign Uj6iw6 = (~(T86iw6 & Bk6iw6));
assign Gj6iw6 = (~(Qa6iw6 & Jz2iw6));
assign Dqd8v6 = (~(Ik6iw6 & Pk6iw6));
assign Pk6iw6 = (~(Ohj7z6[46] & Wk6iw6));
assign Wk6iw6 = (~(V96iw6 & Bk6iw6));
assign Ik6iw6 = (~(Qa6iw6 & Ay2iw6));
assign Wpd8v6 = (~(Dl6iw6 & Kl6iw6));
assign Kl6iw6 = (~(Lgj7z6[183] & Av5iw6));
assign Av5iw6 = (~(Rw2iw6 & Bqi7z6[1]));
assign Dl6iw6 = (~(Rl6iw6 & Rw2iw6));
assign Ppd8v6 = (~(Yl6iw6 & Fm6iw6));
assign Fm6iw6 = (~(Lgj7z6[171] & Cw5iw6));
assign Cw5iw6 = (~(Pv2iw6 & Bqi7z6[1]));
assign Yl6iw6 = (~(Rl6iw6 & Pv2iw6));
assign Ipd8v6 = (~(Mm6iw6 & Tm6iw6));
assign Tm6iw6 = (~(Lgj7z6[159] & Xw5iw6));
assign Xw5iw6 = (~(Nu2iw6 & Bqi7z6[1]));
assign Mm6iw6 = (~(Rl6iw6 & Nu2iw6));
assign Bpd8v6 = (~(An6iw6 & Hn6iw6));
assign Hn6iw6 = (~(Lgj7z6[147] & Sx5iw6));
assign Sx5iw6 = (~(Lt2iw6 & Bqi7z6[1]));
assign An6iw6 = (~(Rl6iw6 & Lt2iw6));
assign Uod8v6 = (~(On6iw6 & Vn6iw6));
assign Vn6iw6 = (~(Lgj7z6[135] & Ny5iw6));
assign Ny5iw6 = (~(Js2iw6 & Bqi7z6[1]));
assign On6iw6 = (~(Rl6iw6 & Js2iw6));
assign Nod8v6 = (~(Co6iw6 & Jo6iw6));
assign Jo6iw6 = (~(Lgj7z6[123] & Iz5iw6));
assign Iz5iw6 = (~(Hr2iw6 & Bqi7z6[1]));
assign Co6iw6 = (~(Rl6iw6 & Hr2iw6));
assign God8v6 = (~(Qo6iw6 & Xo6iw6));
assign Xo6iw6 = (~(Lgj7z6[111] & D06iw6));
assign D06iw6 = (~(Fq2iw6 & Bqi7z6[1]));
assign Qo6iw6 = (~(Rl6iw6 & Fq2iw6));
assign Znd8v6 = (~(Ep6iw6 & Lp6iw6));
assign Lp6iw6 = (~(Lgj7z6[99] & Y06iw6));
assign Y06iw6 = (~(Dp2iw6 & Bqi7z6[1]));
assign Ep6iw6 = (~(Rl6iw6 & Dp2iw6));
assign Snd8v6 = (~(Sp6iw6 & Zp6iw6));
assign Zp6iw6 = (Gq6iw6 | A26iw6);
assign A26iw6 = (~(Wu3iw6 | Nq6iw6));
assign Wu3iw6 = (!Bo2iw6);
assign Sp6iw6 = (~(Rl6iw6 & Bo2iw6));
assign Lnd8v6 = (~(Uq6iw6 & Br6iw6));
assign Br6iw6 = (~(Lgj7z6[75] & V26iw6));
assign V26iw6 = (~(Zm2iw6 & Bqi7z6[1]));
assign Uq6iw6 = (~(Rl6iw6 & Zm2iw6));
assign End8v6 = (~(Ir6iw6 & Pr6iw6));
assign Pr6iw6 = (~(Lgj7z6[63] & Q36iw6));
assign Q36iw6 = (~(Xl2iw6 & Bqi7z6[1]));
assign Ir6iw6 = (~(Rl6iw6 & Xl2iw6));
assign Xmd8v6 = (~(Wr6iw6 & Ds6iw6));
assign Ds6iw6 = (~(Lgj7z6[51] & L46iw6));
assign L46iw6 = (~(Vk2iw6 & Bqi7z6[1]));
assign Wr6iw6 = (~(Rl6iw6 & Vk2iw6));
assign Qmd8v6 = (~(Ks6iw6 & Rs6iw6));
assign Rs6iw6 = (~(Lgj7z6[39] & G56iw6));
assign G56iw6 = (~(Tj2iw6 & Bqi7z6[1]));
assign Ks6iw6 = (~(Rl6iw6 & Tj2iw6));
assign Jmd8v6 = (~(Ys6iw6 & Ft6iw6));
assign Ft6iw6 = (~(Lgj7z6[27] & B66iw6));
assign B66iw6 = (~(Ri2iw6 & Bqi7z6[1]));
assign Ys6iw6 = (~(Rl6iw6 & Ri2iw6));
assign Cmd8v6 = (~(Mt6iw6 & Tt6iw6));
assign Tt6iw6 = (~(Lgj7z6[15] & W66iw6));
assign W66iw6 = (~(Ph2iw6 & Bqi7z6[1]));
assign Mt6iw6 = (~(Rl6iw6 & Ph2iw6));
assign Vld8v6 = (~(Au6iw6 & Hu6iw6));
assign Hu6iw6 = (~(Lgj7z6[3] & R76iw6));
assign R76iw6 = (~(Ng2iw6 & Bqi7z6[1]));
assign Au6iw6 = (~(Rl6iw6 & Ng2iw6));
assign Old8v6 = (~(Ou6iw6 & Vu6iw6));
assign Vu6iw6 = (~(Ohj7z6[13] & Cv6iw6));
assign Cv6iw6 = (~(T86iw6 & Guhov6));
assign Ou6iw6 = (~(Rl6iw6 & Jz2iw6));
assign Hld8v6 = (~(Jv6iw6 & Qv6iw6));
assign Qv6iw6 = (~(Ohj7z6[45] & Xv6iw6));
assign Xv6iw6 = (~(V96iw6 & Guhov6));
assign Jv6iw6 = (~(Rl6iw6 & Ay2iw6));
assign Ald8v6 = (~(Ew6iw6 & Lw6iw6));
assign Lw6iw6 = (~(Ohj7z6[12] & Sw6iw6));
assign Sw6iw6 = (~(T86iw6 & Emhov6));
assign Ew6iw6 = (~(Zw6iw6 & Emhov6));
assign Tkd8v6 = (~(Gx6iw6 & Nx6iw6));
assign Nx6iw6 = (~(Ohj7z6[44] & Ux6iw6));
assign Ux6iw6 = (~(V96iw6 & Emhov6));
assign Gx6iw6 = (~(By6iw6 & Emhov6));
assign Mkd8v6 = (~(Iy6iw6 & Py6iw6));
assign Py6iw6 = (~(Ohj7z6[11] & Wy6iw6));
assign Wy6iw6 = (~(T86iw6 & Dz6iw6));
assign Iy6iw6 = (~(Zw6iw6 & Dz6iw6));
assign Fkd8v6 = (~(Kz6iw6 & Rz6iw6));
assign Rz6iw6 = (~(Ohj7z6[43] & Yz6iw6));
assign Yz6iw6 = (~(V96iw6 & Dz6iw6));
assign Kz6iw6 = (~(By6iw6 & Dz6iw6));
assign Yjd8v6 = (Kkd7v6 ? F07iw6 : N6dov6);
assign F07iw6 = (~(C4dov6 | C477v6));
assign Rjd8v6 = (~(M07iw6 & T07iw6));
assign T07iw6 = (~(Ohj7z6[10] & A17iw6));
assign A17iw6 = (~(T86iw6 & H17iw6));
assign M07iw6 = (~(Zw6iw6 & H17iw6));
assign Kjd8v6 = (~(O17iw6 & V17iw6));
assign V17iw6 = (~(Ohj7z6[42] & C27iw6));
assign C27iw6 = (~(V96iw6 & H17iw6));
assign O17iw6 = (~(By6iw6 & H17iw6));
assign Djd8v6 = (X27iw6 ? Q27iw6 : J27iw6);
assign Q27iw6 = (Dtadt6 | Cr97z6);
assign Wid8v6 = (~(E37iw6 & L37iw6));
assign L37iw6 = (~(Ohj7z6[9] & S37iw6));
assign S37iw6 = (~(T86iw6 & J27iw6));
assign E37iw6 = (~(Zw6iw6 & J27iw6));
assign Pid8v6 = (~(Z37iw6 & G47iw6));
assign G47iw6 = (~(Ohj7z6[41] & N47iw6));
assign N47iw6 = (~(V96iw6 & J27iw6));
assign Z37iw6 = (~(By6iw6 & J27iw6));
assign Iid8v6 = (B57iw6 ? U47iw6 : Dri7z6[8]);
assign Bid8v6 = (B57iw6 ? J27iw6 : Dri7z6[9]);
assign Uhd8v6 = (B57iw6 ? H17iw6 : Dri7z6[10]);
assign Nhd8v6 = (B57iw6 ? Dz6iw6 : Dri7z6[11]);
assign Ghd8v6 = (B57iw6 ? Emhov6 : Dri7z6[12]);
assign Zgd8v6 = (B57iw6 ? Guhov6 : Dri7z6[13]);
assign Sgd8v6 = (B57iw6 ? Bk6iw6 : Dri7z6[14]);
assign Lgd8v6 = (B57iw6 ? Z0iov6 : Dri7z6[15]);
assign B57iw6 = (I57iw6 & Bqi7z6[1]);
assign I57iw6 = (!Kg4iw6);
assign Egd8v6 = (~(P57iw6 & W57iw6));
assign W57iw6 = (~(Ohj7z6[8] & D67iw6));
assign D67iw6 = (~(T86iw6 & U47iw6));
assign T86iw6 = (K67iw6 & Bqi7z6[1]);
assign K67iw6 = (!Mh4iw6);
assign P57iw6 = (~(Zw6iw6 & U47iw6));
assign Zw6iw6 = (Jz2iw6 & Bqi7z6[1]);
assign Xfd8v6 = (~(R67iw6 & Y67iw6));
assign Y67iw6 = (~(Ohj7z6[40] & F77iw6));
assign F77iw6 = (~(V96iw6 & U47iw6));
assign V96iw6 = (M77iw6 & Bqi7z6[1]);
assign M77iw6 = (!Oi4iw6);
assign R67iw6 = (~(By6iw6 & U47iw6));
assign By6iw6 = (Ay2iw6 & Bqi7z6[1]);
assign Qfd8v6 = (~(T77iw6 & A87iw6));
assign A87iw6 = (~(Lgj7z6[182] & H87iw6));
assign T77iw6 = (~(O87iw6 & Rw2iw6));
assign Jfd8v6 = (~(V87iw6 & C97iw6));
assign C97iw6 = (~(Lgj7z6[170] & J97iw6));
assign V87iw6 = (~(O87iw6 & Pv2iw6));
assign Cfd8v6 = (~(Q97iw6 & X97iw6));
assign X97iw6 = (~(Lgj7z6[158] & Ea7iw6));
assign Q97iw6 = (~(O87iw6 & Nu2iw6));
assign Ved8v6 = (~(La7iw6 & Sa7iw6));
assign Sa7iw6 = (~(Lgj7z6[146] & Za7iw6));
assign La7iw6 = (~(O87iw6 & Lt2iw6));
assign Oed8v6 = (~(Gb7iw6 & Nb7iw6));
assign Nb7iw6 = (Ub7iw6 | Bc7iw6);
assign Gb7iw6 = (~(O87iw6 & Js2iw6));
assign Hed8v6 = (~(Ic7iw6 & Pc7iw6));
assign Pc7iw6 = (Wc7iw6 | Dd7iw6);
assign Ic7iw6 = (~(O87iw6 & Hr2iw6));
assign Aed8v6 = (~(Kd7iw6 & Rd7iw6));
assign Rd7iw6 = (Yd7iw6 | Fe7iw6);
assign Kd7iw6 = (~(O87iw6 & Fq2iw6));
assign Tdd8v6 = (~(Me7iw6 & Te7iw6));
assign Te7iw6 = (Af7iw6 | Hf7iw6);
assign Af7iw6 = (!Lgj7z6[98]);
assign Me7iw6 = (~(O87iw6 & Dp2iw6));
assign Mdd8v6 = (~(Of7iw6 & Vf7iw6));
assign Vf7iw6 = (~(Lgj7z6[86] & Cg7iw6));
assign Of7iw6 = (~(O87iw6 & Bo2iw6));
assign Fdd8v6 = (~(Jg7iw6 & Qg7iw6));
assign Qg7iw6 = (~(Lgj7z6[74] & Xg7iw6));
assign Jg7iw6 = (~(O87iw6 & Zm2iw6));
assign Ycd8v6 = (~(Eh7iw6 & Lh7iw6));
assign Lh7iw6 = (Sh7iw6 | Zh7iw6);
assign Eh7iw6 = (~(O87iw6 & Xl2iw6));
assign Rcd8v6 = (~(Gi7iw6 & Ni7iw6));
assign Ni7iw6 = (~(Lgj7z6[50] & Ui7iw6));
assign Gi7iw6 = (~(O87iw6 & Vk2iw6));
assign Kcd8v6 = (~(Bj7iw6 & Ij7iw6));
assign Ij7iw6 = (~(Lgj7z6[38] & Pj7iw6));
assign Bj7iw6 = (~(O87iw6 & Tj2iw6));
assign Dcd8v6 = (~(Wj7iw6 & Dk7iw6));
assign Dk7iw6 = (Kk7iw6 | Rk7iw6);
assign Wj7iw6 = (~(O87iw6 & Ri2iw6));
assign Wbd8v6 = (~(Yk7iw6 & Fl7iw6));
assign Fl7iw6 = (Ml7iw6 | Tl7iw6);
assign Yk7iw6 = (~(O87iw6 & Ph2iw6));
assign Pbd8v6 = (~(Am7iw6 & Hm7iw6));
assign Hm7iw6 = (~(Lgj7z6[2] & Om7iw6));
assign Am7iw6 = (~(O87iw6 & Ng2iw6));
assign Ibd8v6 = (~(Vm7iw6 & Cn7iw6));
assign Cn7iw6 = (~(Ohj7z6[7] & Jn7iw6));
assign Jn7iw6 = (~(Qn7iw6 & R62nv6));
assign Vm7iw6 = (~(O87iw6 & Jz2iw6));
assign Bbd8v6 = (~(Xn7iw6 & Eo7iw6));
assign Eo7iw6 = (~(Ohj7z6[39] & Lo7iw6));
assign Lo7iw6 = (~(So7iw6 & R62nv6));
assign Xn7iw6 = (~(O87iw6 & Ay2iw6));
assign Uad8v6 = (~(Zo7iw6 & Gp7iw6));
assign Gp7iw6 = (~(Lgj7z6[181] & H87iw6));
assign Zo7iw6 = (~(Np7iw6 & Rw2iw6));
assign Nad8v6 = (~(Up7iw6 & Bq7iw6));
assign Bq7iw6 = (~(Lgj7z6[169] & J97iw6));
assign Up7iw6 = (~(Np7iw6 & Pv2iw6));
assign Gad8v6 = (~(Iq7iw6 & Pq7iw6));
assign Pq7iw6 = (~(Lgj7z6[157] & Ea7iw6));
assign Iq7iw6 = (~(Np7iw6 & Nu2iw6));
assign Z9d8v6 = (~(Wq7iw6 & Dr7iw6));
assign Dr7iw6 = (~(Lgj7z6[145] & Za7iw6));
assign Wq7iw6 = (~(Np7iw6 & Lt2iw6));
assign S9d8v6 = (~(Kr7iw6 & Rr7iw6));
assign Rr7iw6 = (Yr7iw6 | Bc7iw6);
assign Kr7iw6 = (~(Np7iw6 & Js2iw6));
assign L9d8v6 = (~(Fs7iw6 & Ms7iw6));
assign Ms7iw6 = (Ts7iw6 | Dd7iw6);
assign Fs7iw6 = (~(Np7iw6 & Hr2iw6));
assign E9d8v6 = (~(At7iw6 & Ht7iw6));
assign Ht7iw6 = (Ot7iw6 | Fe7iw6);
assign At7iw6 = (~(Np7iw6 & Fq2iw6));
assign X8d8v6 = (~(Vt7iw6 & Cu7iw6));
assign Cu7iw6 = (Ju7iw6 | Hf7iw6);
assign Vt7iw6 = (~(Np7iw6 & Dp2iw6));
assign Q8d8v6 = (~(Qu7iw6 & Xu7iw6));
assign Xu7iw6 = (~(Lgj7z6[85] & Cg7iw6));
assign Qu7iw6 = (~(Np7iw6 & Bo2iw6));
assign J8d8v6 = (~(Ev7iw6 & Lv7iw6));
assign Lv7iw6 = (~(Lgj7z6[73] & Xg7iw6));
assign Ev7iw6 = (~(Np7iw6 & Zm2iw6));
assign C8d8v6 = (~(Sv7iw6 & Zv7iw6));
assign Zv7iw6 = (Gw7iw6 | Zh7iw6);
assign Sv7iw6 = (~(Np7iw6 & Xl2iw6));
assign V7d8v6 = (~(Nw7iw6 & Uw7iw6));
assign Uw7iw6 = (~(Lgj7z6[49] & Ui7iw6));
assign Nw7iw6 = (~(Np7iw6 & Vk2iw6));
assign O7d8v6 = (~(Bx7iw6 & Ix7iw6));
assign Ix7iw6 = (~(Lgj7z6[37] & Pj7iw6));
assign Bx7iw6 = (~(Np7iw6 & Tj2iw6));
assign H7d8v6 = (~(Px7iw6 & Wx7iw6));
assign Wx7iw6 = (Dy7iw6 | Rk7iw6);
assign Px7iw6 = (~(Np7iw6 & Ri2iw6));
assign A7d8v6 = (~(Ky7iw6 & Ry7iw6));
assign Ry7iw6 = (Yy7iw6 | Tl7iw6);
assign Ky7iw6 = (~(Np7iw6 & Ph2iw6));
assign T6d8v6 = (~(Fz7iw6 & Mz7iw6));
assign Mz7iw6 = (~(Lgj7z6[1] & Om7iw6));
assign Fz7iw6 = (~(Np7iw6 & Ng2iw6));
assign M6d8v6 = (~(Tz7iw6 & A08iw6));
assign A08iw6 = (~(Ohj7z6[6] & H08iw6));
assign H08iw6 = (~(Qn7iw6 & K62nv6));
assign Tz7iw6 = (~(Np7iw6 & Jz2iw6));
assign F6d8v6 = (~(O08iw6 & V08iw6));
assign V08iw6 = (~(Ohj7z6[38] & C18iw6));
assign C18iw6 = (~(So7iw6 & K62nv6));
assign O08iw6 = (~(Np7iw6 & Ay2iw6));
assign Y5d8v6 = (~(J18iw6 & Q18iw6));
assign Q18iw6 = (~(Lgj7z6[180] & H87iw6));
assign H87iw6 = (~(Rw2iw6 & Bqi7z6[0]));
assign J18iw6 = (~(X18iw6 & Rw2iw6));
assign Rw2iw6 = (E28iw6 & L28iw6);
assign R5d8v6 = (~(S28iw6 & Z28iw6));
assign Z28iw6 = (~(Lgj7z6[168] & J97iw6));
assign J97iw6 = (~(Pv2iw6 & Bqi7z6[0]));
assign S28iw6 = (~(X18iw6 & Pv2iw6));
assign Pv2iw6 = (~(G38iw6 | N38iw6));
assign K5d8v6 = (~(U38iw6 & B48iw6));
assign B48iw6 = (~(Lgj7z6[156] & Ea7iw6));
assign Ea7iw6 = (~(Nu2iw6 & Bqi7z6[0]));
assign U38iw6 = (~(X18iw6 & Nu2iw6));
assign Nu2iw6 = (~(I48iw6 | P48iw6));
assign D5d8v6 = (~(W48iw6 & D58iw6));
assign D58iw6 = (~(Lgj7z6[144] & Za7iw6));
assign Za7iw6 = (~(Lt2iw6 & Bqi7z6[0]));
assign W48iw6 = (~(X18iw6 & Lt2iw6));
assign Lt2iw6 = (K58iw6 & R58iw6);
assign K58iw6 = (!G38iw6);
assign W4d8v6 = (~(Y58iw6 & F68iw6));
assign F68iw6 = (M68iw6 | Bc7iw6);
assign Bc7iw6 = (Js2iw6 & Bqi7z6[0]);
assign Y58iw6 = (~(X18iw6 & Js2iw6));
assign Js2iw6 = (E28iw6 & T68iw6);
assign E28iw6 = (!I48iw6);
assign P4d8v6 = (~(A78iw6 & H78iw6));
assign H78iw6 = (O78iw6 | Dd7iw6);
assign Dd7iw6 = (Hr2iw6 & Bqi7z6[0]);
assign A78iw6 = (~(X18iw6 & Hr2iw6));
assign Hr2iw6 = (~(G38iw6 | V78iw6));
assign I4d8v6 = (~(C88iw6 & J88iw6));
assign J88iw6 = (Q88iw6 | Fe7iw6);
assign Fe7iw6 = (Fq2iw6 & Bqi7z6[0]);
assign C88iw6 = (~(X18iw6 & Fq2iw6));
assign Fq2iw6 = (~(I48iw6 | X88iw6));
assign I48iw6 = (~(E98iw6 & L98iw6));
assign L98iw6 = (S98iw6 & Toi7z6[10]);
assign E98iw6 = (Z98iw6 & Toi7z6[2]);
assign B4d8v6 = (~(Ga8iw6 & Na8iw6));
assign Na8iw6 = (Ua8iw6 | Hf7iw6);
assign Hf7iw6 = (Dp2iw6 & Bqi7z6[0]);
assign Ga8iw6 = (~(X18iw6 & Dp2iw6));
assign Dp2iw6 = (~(G38iw6 | X88iw6));
assign G38iw6 = (~(Bb8iw6 & Ib8iw6));
assign Ib8iw6 = (Toi7z6[10] & Pb8iw6);
assign Bb8iw6 = (Z98iw6 & S98iw6);
assign U3d8v6 = (~(Wb8iw6 & Dc8iw6));
assign Dc8iw6 = (~(Lgj7z6[84] & Cg7iw6));
assign Cg7iw6 = (~(Bo2iw6 & Bqi7z6[0]));
assign Wb8iw6 = (~(X18iw6 & Bo2iw6));
assign Bo2iw6 = (~(N38iw6 | Kc8iw6));
assign N3d8v6 = (~(Rc8iw6 & Yc8iw6));
assign Yc8iw6 = (~(Lgj7z6[72] & Xg7iw6));
assign Xg7iw6 = (~(Zm2iw6 & Bqi7z6[0]));
assign Rc8iw6 = (~(X18iw6 & Zm2iw6));
assign Zm2iw6 = (~(N38iw6 | Fd8iw6));
assign N38iw6 = (!L28iw6);
assign G3d8v6 = (~(Md8iw6 & Td8iw6));
assign Td8iw6 = (Ae8iw6 | Zh7iw6);
assign Zh7iw6 = (Xl2iw6 & Bqi7z6[0]);
assign Md8iw6 = (~(X18iw6 & Xl2iw6));
assign Xl2iw6 = (~(Kc8iw6 | P48iw6));
assign Z2d8v6 = (~(He8iw6 & Oe8iw6));
assign Oe8iw6 = (~(Lgj7z6[48] & Ui7iw6));
assign Ui7iw6 = (~(Vk2iw6 & Bqi7z6[0]));
assign He8iw6 = (~(X18iw6 & Vk2iw6));
assign Vk2iw6 = (Ve8iw6 & R58iw6);
assign S2d8v6 = (~(Cf8iw6 & Jf8iw6));
assign Jf8iw6 = (~(Lgj7z6[36] & Pj7iw6));
assign Pj7iw6 = (~(Tj2iw6 & Bqi7z6[0]));
assign Cf8iw6 = (~(X18iw6 & Tj2iw6));
assign Tj2iw6 = (~(Kc8iw6 | V78iw6));
assign L2d8v6 = (~(Qf8iw6 & Xf8iw6));
assign Xf8iw6 = (Eg8iw6 | Rk7iw6);
assign Rk7iw6 = (Ri2iw6 & Bqi7z6[0]);
assign Qf8iw6 = (~(X18iw6 & Ri2iw6));
assign Ri2iw6 = (~(Fd8iw6 | V78iw6));
assign V78iw6 = (!T68iw6);
assign E2d8v6 = (~(Lg8iw6 & Sg8iw6));
assign Sg8iw6 = (Zg8iw6 | Tl7iw6);
assign Tl7iw6 = (Ph2iw6 & Bqi7z6[0]);
assign Lg8iw6 = (~(X18iw6 & Ph2iw6));
assign Ph2iw6 = (~(Kc8iw6 | X88iw6));
assign Kc8iw6 = (Gh8iw6 | Pb8iw6);
assign X1d8v6 = (~(Nh8iw6 & Uh8iw6));
assign Uh8iw6 = (~(Lgj7z6[0] & Om7iw6));
assign Om7iw6 = (~(Ng2iw6 & Bqi7z6[0]));
assign Nh8iw6 = (~(X18iw6 & Ng2iw6));
assign Ng2iw6 = (~(Fd8iw6 | X88iw6));
assign Fd8iw6 = (!Ve8iw6);
assign Ve8iw6 = (Bi8iw6 & Pb8iw6);
assign Bi8iw6 = (!Gh8iw6);
assign Gh8iw6 = (~(Ii8iw6 & Z98iw6));
assign Ii8iw6 = (Pi8iw6 & Toi7z6[10]);
assign Q1d8v6 = (~(Wi8iw6 & Dj8iw6));
assign Dj8iw6 = (~(Ohj7z6[5] & Kj8iw6));
assign Kj8iw6 = (~(Qn7iw6 & D62nv6));
assign Wi8iw6 = (~(X18iw6 & Jz2iw6));
assign J1d8v6 = (~(Rj8iw6 & Yj8iw6));
assign Yj8iw6 = (~(Ohj7z6[37] & Fk8iw6));
assign Fk8iw6 = (~(So7iw6 & D62nv6));
assign Rj8iw6 = (~(X18iw6 & Ay2iw6));
assign C1d8v6 = (Al8iw6 ? Tk8iw6 : Mk8iw6);
assign Al8iw6 = (Hl8iw6 & Esadt6);
assign Hl8iw6 = (Rabov6 & Mrnov6);
assign Mk8iw6 = (Cngdt6 & Ol8iw6);
assign V0d8v6 = (Vl8iw6 & Rabov6);
assign Vl8iw6 = (Tk8iw6 & Cm8iw6);
assign Cm8iw6 = (~(Jm8iw6 & Qm8iw6));
assign Qm8iw6 = (~(Esadt6 & Mrnov6));
assign O0d8v6 = (~(Xm8iw6 & En8iw6));
assign En8iw6 = (~(Bxi7z6[4] & Ln8iw6));
assign Ln8iw6 = (~(O8fov6 & W52nv6));
assign Xm8iw6 = (~(C9fov6 & Sn8iw6));
assign C9fov6 = (~(Zn8iw6 & Go8iw6));
assign Go8iw6 = (~(Q7hov6 & Vm2nv6));
assign Zn8iw6 = (~(Fe2nv6 & Ldo7v6));
assign H0d8v6 = (~(No8iw6 & Uo8iw6));
assign Uo8iw6 = (~(Ohj7z6[4] & Bp8iw6));
assign Bp8iw6 = (~(Qn7iw6 & W52nv6));
assign No8iw6 = (~(Ip8iw6 & W52nv6));
assign A0d8v6 = (~(Pp8iw6 & Wp8iw6));
assign Wp8iw6 = (~(Ohj7z6[36] & Dq8iw6));
assign Dq8iw6 = (~(So7iw6 & W52nv6));
assign Pp8iw6 = (~(Kq8iw6 & W52nv6));
assign Tzc8v6 = (~(Rq8iw6 & Yq8iw6));
assign Yq8iw6 = (~(Fr8iw6 & B8cdt6));
assign Fr8iw6 = (Mr8iw6 & Tr8iw6);
assign Mr8iw6 = (~(As8iw6 & Hs8iw6));
assign Hs8iw6 = (~(Mqhhw6 | Wwvnv6));
assign As8iw6 = (Os8iw6 & Vs8iw6);
assign Vs8iw6 = (~(Dradt6 & Ct8iw6));
assign Ct8iw6 = (Yqvnv6 | Kxvnv6);
assign Os8iw6 = (~(Yqvnv6 & Mzfhw6));
assign Rq8iw6 = (~(W5fhw6 & Ez2et6));
assign W5fhw6 = (~(Jt8iw6 | Qt8iw6));
assign Qt8iw6 = (~(Gaonv6 | Zwehw6));
assign Jt8iw6 = (I2jnv6 ? Gr2et6 : Xt8iw6);
assign Xt8iw6 = (Tfh7z6[0] | Tfh7z6[1]);
assign Mzc8v6 = (~(Eu8iw6 & Lu8iw6));
assign Lu8iw6 = (~(Ohj7z6[3] & Su8iw6));
assign Su8iw6 = (~(Qn7iw6 & P52nv6));
assign Eu8iw6 = (~(Ip8iw6 & P52nv6));
assign Fzc8v6 = (~(Zu8iw6 & Gv8iw6));
assign Gv8iw6 = (~(Ohj7z6[35] & Nv8iw6));
assign Nv8iw6 = (~(So7iw6 & P52nv6));
assign Zu8iw6 = (~(Kq8iw6 & P52nv6));
assign Yyc8v6 = (Uv8iw6 ? Apget6 : I52nv6);
assign Ryc8v6 = (~(Bw8iw6 & Iw8iw6));
assign Iw8iw6 = (~(Ohj7z6[2] & Pw8iw6));
assign Pw8iw6 = (~(Qn7iw6 & I52nv6));
assign Bw8iw6 = (~(Ip8iw6 & I52nv6));
assign Kyc8v6 = (~(Ww8iw6 & Dx8iw6));
assign Dx8iw6 = (~(Ohj7z6[34] & Kx8iw6));
assign Kx8iw6 = (~(So7iw6 & I52nv6));
assign Ww8iw6 = (~(Kq8iw6 & I52nv6));
assign Dyc8v6 = (Uv8iw6 ? Weget6 : B52nv6);
assign Uv8iw6 = (!Rx8iw6);
assign Wxc8v6 = (~(Yx8iw6 & Fy8iw6));
assign Fy8iw6 = (~(Ohj7z6[1] & My8iw6));
assign My8iw6 = (~(Qn7iw6 & B52nv6));
assign Yx8iw6 = (~(Ip8iw6 & B52nv6));
assign Pxc8v6 = (~(Ty8iw6 & Az8iw6));
assign Az8iw6 = (~(Ohj7z6[33] & Hz8iw6));
assign Hz8iw6 = (~(So7iw6 & B52nv6));
assign Ty8iw6 = (~(Kq8iw6 & B52nv6));
assign Ixc8v6 = (!Oz8iw6);
assign Oz8iw6 = (J09iw6 ? C09iw6 : Vz8iw6);
assign Bxc8v6 = (~(Q09iw6 & X09iw6));
assign X09iw6 = (E19iw6 | L19iw6);
assign Q09iw6 = (~(J09iw6 & Hyj7z6[6]));
assign Uwc8v6 = (~(S19iw6 & Z19iw6));
assign Z19iw6 = (B52nv6 | E19iw6);
assign E19iw6 = (~(G29iw6 & Orhov6));
assign G29iw6 = (N29iw6 & I52nv6);
assign S19iw6 = (~(J09iw6 & Hyj7z6[4]));
assign Nwc8v6 = (~(U29iw6 & B39iw6));
assign B39iw6 = (~(I39iw6 & P39iw6));
assign U29iw6 = (~(J09iw6 & Hyj7z6[2]));
assign Gwc8v6 = (~(W39iw6 & D49iw6));
assign D49iw6 = (~(K49iw6 & P39iw6));
assign W39iw6 = (~(J09iw6 & Hyj7z6[0]));
assign Zvc8v6 = (Rx8iw6 ? U42nv6 : Phget6);
assign Rx8iw6 = (R49iw6 & Y49iw6);
assign Y49iw6 = (F59iw6 & Dtj7z6[4]);
assign F59iw6 = (M59iw6 & T59iw6);
assign R49iw6 = (Hc3iw6 & Dtj7z6[2]);
assign Svc8v6 = (~(A69iw6 & H69iw6));
assign H69iw6 = (~(O69iw6 & V69iw6));
assign V69iw6 = (C79iw6 & J79iw6);
assign O69iw6 = (Q79iw6 & Jjbdt6);
assign A69iw6 = (~(X79iw6 & E89iw6));
assign E89iw6 = (~(L89iw6 & C79iw6));
assign C79iw6 = (S89iw6 & Jolov6);
assign S89iw6 = (~(Gr2et6 & Puphw6));
assign L89iw6 = (Q79iw6 & J79iw6);
assign J79iw6 = (~(Zgnov6 & J2cdt6));
assign Zgnov6 = (Z89iw6 & G99iw6);
assign G99iw6 = (~(Z7edt6 | Tnzdt6));
assign Z89iw6 = (Ibe7z6[4] & N99iw6);
assign Q79iw6 = (U99iw6 & Ba9iw6);
assign Ba9iw6 = (~(Ia9iw6 & Eyknv6));
assign Ia9iw6 = (O5a7z6 & Venov6);
assign U99iw6 = (Pa9iw6 & Lhfov6);
assign Pa9iw6 = (~(Tnzdt6 & Wa9iw6));
assign Wa9iw6 = (~(Db9iw6 & Kb9iw6));
assign Db9iw6 = (~(Rb9iw6 & Kioov6));
assign X79iw6 = (~(Yb9iw6 & Fc9iw6));
assign Fc9iw6 = (~(Ibe7z6[4] & E3c7z6[1]));
assign Yb9iw6 = (Mc9iw6 & Tc9iw6);
assign Tc9iw6 = (Jolov6 | Ad9iw6);
assign Jolov6 = (Dxvnv6 | Hd9iw6);
assign Mc9iw6 = (~(Rkfov6 & Od9iw6));
assign Rkfov6 = (!Lhfov6);
assign Lhfov6 = (~(Vd9iw6 & Ce9iw6));
assign Vd9iw6 = (Qij7z6[2] & Gvvnv6);
assign Lvc8v6 = (~(Je9iw6 & Qe9iw6));
assign Qe9iw6 = (Xe9iw6 & Ef9iw6);
assign Ef9iw6 = (~(Ohe7z6[5] & Okaov6));
assign Okaov6 = (N4mov6 | Upfov6);
assign Xe9iw6 = (Lf9iw6 & Sf9iw6);
assign Sf9iw6 = (~(Jlaov6 & Zec7z6[5]));
assign Lf9iw6 = (~(Qlaov6 & Xumov6));
assign Je9iw6 = (Zf9iw6 & Gg9iw6);
assign Gg9iw6 = (Smaov6 | Ivaov6);
assign Ivaov6 = (!Ng9iw6);
assign Zf9iw6 = (~(Gnaov6 & Zec7z6[21]));
assign Evc8v6 = (~(B5mov6 & Ug9iw6));
assign Ug9iw6 = (~(Upfov6 & Ohe7z6[4]));
assign B5mov6 = (Bh9iw6 & Ih9iw6);
assign Ih9iw6 = (~(Ph9iw6 & X2mov6));
assign Bh9iw6 = (Wh9iw6 & Di9iw6);
assign Di9iw6 = (~(Ki9iw6 & Z3mov6));
assign Ki9iw6 = (G4mov6 ? Zec7z6[3] : Zec7z6[19]);
assign Wh9iw6 = (~(N4mov6 & Ohe7z6[3]));
assign Xuc8v6 = (~(Ri9iw6 & Yi9iw6));
assign Yi9iw6 = (Fj9iw6 & Mj9iw6);
assign Mj9iw6 = (Smaov6 | Bvaov6);
assign Bvaov6 = (!Tj9iw6);
assign Smaov6 = (~(X2mov6 & Ak9iw6));
assign Ak9iw6 = (~(Staov6 & Hk9iw6));
assign Staov6 = (Ok9iw6 & Vk9iw6);
assign Vk9iw6 = (Cl9iw6 & Jl9iw6);
assign Ok9iw6 = (Ql9iw6 & Xl9iw6);
assign Fj9iw6 = (Em9iw6 & Lm9iw6);
assign Lm9iw6 = (~(Jlaov6 & Zec7z6[4]));
assign Jlaov6 = (~(P5mov6 | Gnaov6));
assign Em9iw6 = (~(Qlaov6 & Pxmov6));
assign Qlaov6 = (~(Hk9iw6 | Hulov6));
assign Ri9iw6 = (Sm9iw6 & Zm9iw6);
assign Zm9iw6 = (~(Gnaov6 & Zec7z6[20]));
assign Gnaov6 = (!G4mov6);
assign Sm9iw6 = (Gn9iw6 & Nn9iw6);
assign Nn9iw6 = (~(Upfov6 & N0gdt6));
assign Gn9iw6 = (~(N4mov6 & Ohe7z6[4]));
assign Quc8v6 = (~(U4mov6 & Un9iw6));
assign Un9iw6 = (~(Upfov6 & Ohe7z6[1]));
assign U4mov6 = (Bo9iw6 & Io9iw6);
assign Io9iw6 = (~(Od9iw6 & X2mov6));
assign X2mov6 = (~(Po9iw6 & Wo9iw6));
assign Wo9iw6 = (~(Dp9iw6 & Hulov6));
assign Dp9iw6 = (!Hk9iw6);
assign Hk9iw6 = (~(Kp9iw6 & Rp9iw6));
assign Rp9iw6 = (Yp9iw6 & Kb9iw6);
assign Yp9iw6 = (Fiihw6 & Elphw6);
assign Kp9iw6 = (Fq9iw6 & Mq9iw6);
assign Fq9iw6 = (Tq9iw6 & Ar9iw6);
assign Ar9iw6 = (!M0mov6);
assign Bo9iw6 = (~(Hr9iw6 & Z3mov6));
assign Z3mov6 = (!P5mov6);
assign Hr9iw6 = (G4mov6 ? Zec7z6[0] : Zec7z6[16]);
assign Juc8v6 = (Qu1ov6 ? Or9iw6 : Qmb7z6[1]);
assign Cuc8v6 = (Qu1ov6 ? Vr9iw6 : Qmb7z6[2]);
assign Vtc8v6 = (Qu1ov6 ? Cs9iw6 : Qmb7z6[3]);
assign Otc8v6 = (Qu1ov6 ? Js9iw6 : Qmb7z6[4]);
assign Htc8v6 = (Qu1ov6 ? Qs9iw6 : Qmb7z6[5]);
assign Atc8v6 = (Qu1ov6 ? Xs9iw6 : Qmb7z6[6]);
assign Tsc8v6 = (Qu1ov6 ? Zwlov6 : Qmb7z6[7]);
assign Msc8v6 = (Qu1ov6 ? Et9iw6 : Qmb7z6[8]);
assign Fsc8v6 = (Qu1ov6 ? Swlov6 : Qmb7z6[0]);
assign Rrc8v6 = (~(Lt9iw6 & St9iw6));
assign St9iw6 = (~(Zt9iw6 & A0j7z6[0]));
assign Lt9iw6 = (Gu9iw6 & Nu9iw6);
assign Nu9iw6 = (~(Uu9iw6 & H1j7z6[0]));
assign Gu9iw6 = (~(Oldet6 & Bv9iw6));
assign Krc8v6 = (~(Iv9iw6 & Pv9iw6));
assign Pv9iw6 = (~(Zt9iw6 & A0j7z6[1]));
assign Iv9iw6 = (Wv9iw6 & Dw9iw6);
assign Dw9iw6 = (~(Uu9iw6 & H1j7z6[1]));
assign Wv9iw6 = (~(Akdet6 & Bv9iw6));
assign Drc8v6 = (~(Kw9iw6 & Rw9iw6));
assign Rw9iw6 = (~(Zt9iw6 & A0j7z6[2]));
assign Kw9iw6 = (Yw9iw6 & Fx9iw6);
assign Fx9iw6 = (~(Uu9iw6 & H1j7z6[2]));
assign Yw9iw6 = (~(Midet6 & Bv9iw6));
assign Wqc8v6 = (~(Mx9iw6 & Tx9iw6));
assign Tx9iw6 = (~(Zt9iw6 & A0j7z6[3]));
assign Mx9iw6 = (Ay9iw6 & Hy9iw6);
assign Hy9iw6 = (~(Uu9iw6 & H1j7z6[3]));
assign Ay9iw6 = (~(Ygdet6 & Bv9iw6));
assign Pqc8v6 = (~(Oy9iw6 & Vy9iw6));
assign Vy9iw6 = (~(Zt9iw6 & A0j7z6[4]));
assign Oy9iw6 = (Cz9iw6 & Jz9iw6);
assign Jz9iw6 = (~(Uu9iw6 & H1j7z6[4]));
assign Cz9iw6 = (~(Kfdet6 & Bv9iw6));
assign Iqc8v6 = (~(Qz9iw6 & Xz9iw6));
assign Xz9iw6 = (~(Zt9iw6 & A0j7z6[5]));
assign Qz9iw6 = (E0aiw6 & L0aiw6);
assign L0aiw6 = (~(Uu9iw6 & H1j7z6[5]));
assign E0aiw6 = (~(Wddet6 & Bv9iw6));
assign Bqc8v6 = (~(S0aiw6 & Z0aiw6));
assign Z0aiw6 = (~(Zt9iw6 & A0j7z6[6]));
assign S0aiw6 = (G1aiw6 & N1aiw6);
assign N1aiw6 = (~(Uu9iw6 & H1j7z6[6]));
assign G1aiw6 = (~(Icdet6 & Bv9iw6));
assign Upc8v6 = (~(U1aiw6 & B2aiw6));
assign B2aiw6 = (~(Zt9iw6 & A0j7z6[7]));
assign U1aiw6 = (I2aiw6 & P2aiw6);
assign P2aiw6 = (~(Uu9iw6 & H1j7z6[7]));
assign I2aiw6 = (~(Uadet6 & Bv9iw6));
assign Npc8v6 = (~(W2aiw6 & D3aiw6));
assign D3aiw6 = (~(Zt9iw6 & A0j7z6[8]));
assign W2aiw6 = (K3aiw6 & R3aiw6);
assign R3aiw6 = (~(Uu9iw6 & H1j7z6[8]));
assign K3aiw6 = (~(G9det6 & Bv9iw6));
assign Gpc8v6 = (~(Y3aiw6 & F4aiw6));
assign F4aiw6 = (~(Zt9iw6 & A0j7z6[9]));
assign Y3aiw6 = (M4aiw6 & T4aiw6);
assign T4aiw6 = (~(Uu9iw6 & H1j7z6[9]));
assign M4aiw6 = (~(S7det6 & Bv9iw6));
assign Zoc8v6 = (~(A5aiw6 & H5aiw6));
assign H5aiw6 = (~(Zt9iw6 & A0j7z6[10]));
assign A5aiw6 = (O5aiw6 & V5aiw6);
assign V5aiw6 = (~(Uu9iw6 & H1j7z6[10]));
assign O5aiw6 = (~(E6det6 & Bv9iw6));
assign Soc8v6 = (~(C6aiw6 & J6aiw6));
assign J6aiw6 = (~(Zt9iw6 & A0j7z6[11]));
assign C6aiw6 = (Q6aiw6 & X6aiw6);
assign X6aiw6 = (~(Uu9iw6 & H1j7z6[11]));
assign Q6aiw6 = (~(Q4det6 & Bv9iw6));
assign Loc8v6 = (~(E7aiw6 & L7aiw6));
assign L7aiw6 = (~(Zt9iw6 & A0j7z6[12]));
assign E7aiw6 = (S7aiw6 & Z7aiw6);
assign Z7aiw6 = (~(Uu9iw6 & H1j7z6[12]));
assign S7aiw6 = (~(C3det6 & Bv9iw6));
assign Eoc8v6 = (~(G8aiw6 & N8aiw6));
assign N8aiw6 = (~(Zt9iw6 & A0j7z6[13]));
assign G8aiw6 = (U8aiw6 & B9aiw6);
assign B9aiw6 = (~(Uu9iw6 & H1j7z6[13]));
assign U8aiw6 = (~(O1det6 & Bv9iw6));
assign Xnc8v6 = (~(I9aiw6 & P9aiw6));
assign P9aiw6 = (~(Zt9iw6 & A0j7z6[14]));
assign I9aiw6 = (W9aiw6 & Daaiw6);
assign Daaiw6 = (~(Uu9iw6 & H1j7z6[14]));
assign W9aiw6 = (~(A0det6 & Bv9iw6));
assign Qnc8v6 = (~(Kaaiw6 & Raaiw6));
assign Raaiw6 = (~(Zt9iw6 & A0j7z6[15]));
assign Kaaiw6 = (Yaaiw6 & Fbaiw6);
assign Fbaiw6 = (~(Uu9iw6 & H1j7z6[15]));
assign Yaaiw6 = (~(Mycet6 & Bv9iw6));
assign Jnc8v6 = (~(Mbaiw6 & Tbaiw6));
assign Tbaiw6 = (~(Zt9iw6 & A0j7z6[16]));
assign Mbaiw6 = (Acaiw6 & Hcaiw6);
assign Hcaiw6 = (~(Uu9iw6 & H1j7z6[16]));
assign Acaiw6 = (~(Ywcet6 & Bv9iw6));
assign Cnc8v6 = (~(Ocaiw6 & Vcaiw6));
assign Vcaiw6 = (~(Zt9iw6 & A0j7z6[17]));
assign Ocaiw6 = (Cdaiw6 & Jdaiw6);
assign Jdaiw6 = (~(Uu9iw6 & H1j7z6[17]));
assign Cdaiw6 = (~(Kvcet6 & Bv9iw6));
assign Vmc8v6 = (~(Qdaiw6 & Xdaiw6));
assign Xdaiw6 = (~(Zt9iw6 & A0j7z6[18]));
assign Qdaiw6 = (Eeaiw6 & Leaiw6);
assign Leaiw6 = (~(Uu9iw6 & H1j7z6[18]));
assign Eeaiw6 = (~(Wtcet6 & Bv9iw6));
assign Omc8v6 = (~(Seaiw6 & Zeaiw6));
assign Zeaiw6 = (~(Zt9iw6 & A0j7z6[19]));
assign Seaiw6 = (Gfaiw6 & Nfaiw6);
assign Nfaiw6 = (~(Uu9iw6 & H1j7z6[19]));
assign Gfaiw6 = (~(Iscet6 & Bv9iw6));
assign Hmc8v6 = (~(Ufaiw6 & Bgaiw6));
assign Bgaiw6 = (~(Zt9iw6 & A0j7z6[20]));
assign Ufaiw6 = (Igaiw6 & Pgaiw6);
assign Pgaiw6 = (~(Uu9iw6 & H1j7z6[20]));
assign Igaiw6 = (~(Uqcet6 & Bv9iw6));
assign Amc8v6 = (~(Wgaiw6 & Dhaiw6));
assign Dhaiw6 = (~(Zt9iw6 & A0j7z6[21]));
assign Wgaiw6 = (Khaiw6 & Rhaiw6);
assign Rhaiw6 = (~(Uu9iw6 & H1j7z6[21]));
assign Khaiw6 = (~(Gpcet6 & Bv9iw6));
assign Tlc8v6 = (~(Yhaiw6 & Fiaiw6));
assign Fiaiw6 = (~(Zt9iw6 & A0j7z6[22]));
assign Yhaiw6 = (Miaiw6 & Tiaiw6);
assign Tiaiw6 = (~(Uu9iw6 & H1j7z6[22]));
assign Miaiw6 = (~(Sncet6 & Bv9iw6));
assign Mlc8v6 = (~(Ajaiw6 & Hjaiw6));
assign Hjaiw6 = (~(Zt9iw6 & A0j7z6[23]));
assign Ajaiw6 = (Ojaiw6 & Vjaiw6);
assign Vjaiw6 = (~(Uu9iw6 & H1j7z6[23]));
assign Uu9iw6 = (~(Ckaiw6 | Jkaiw6));
assign Ckaiw6 = (Zt9iw6 | Qkaiw6);
assign Ojaiw6 = (~(Emcet6 & Bv9iw6));
assign Bv9iw6 = (Xkaiw6 & Jkaiw6);
assign Jkaiw6 = (~(Elaiw6 & Llaiw6));
assign Llaiw6 = (!A0j7z6[0]);
assign Xkaiw6 = (~(Zt9iw6 | Qkaiw6));
assign Zt9iw6 = (~(Slaiw6 | Qkaiw6));
assign Qkaiw6 = (!Zlaiw6);
assign Flc8v6 = (~(Gmaiw6 & Nmaiw6));
assign Nmaiw6 = (~(Umaiw6 & Macet6));
assign Umaiw6 = (Bnaiw6 & Zlaiw6);
assign Bnaiw6 = (~(Inaiw6 & Pnaiw6));
assign Pnaiw6 = (F52iw6 & Wnaiw6);
assign Inaiw6 = (Doaiw6 & Koaiw6);
assign Gmaiw6 = (~(Roaiw6 & Slaiw6));
assign Roaiw6 = (Elaiw6 & A0j7z6[0]);
assign Ykc8v6 = (Yoaiw6 & Fpaiw6);
assign Fpaiw6 = (E9cet6 & A0j7z6[0]);
assign Yoaiw6 = (Slaiw6 & Elaiw6);
assign Elaiw6 = (Mpaiw6 & Tpaiw6);
assign Tpaiw6 = (Aqaiw6 & Hqaiw6);
assign Hqaiw6 = (Oqaiw6 & Vqaiw6);
assign Vqaiw6 = (~(Craiw6 | A0j7z6[7]));
assign Craiw6 = (A0j7z6[8] | A0j7z6[9]);
assign Oqaiw6 = (~(Jraiw6 | A0j7z6[4]));
assign Jraiw6 = (A0j7z6[5] | A0j7z6[6]);
assign Aqaiw6 = (Qraiw6 & Xraiw6);
assign Xraiw6 = (~(Esaiw6 | A0j7z6[23]));
assign Esaiw6 = (A0j7z6[2] | A0j7z6[3]);
assign Qraiw6 = (~(Lsaiw6 | A0j7z6[20]));
assign Lsaiw6 = (A0j7z6[21] | A0j7z6[22]);
assign Mpaiw6 = (Ssaiw6 & Zsaiw6);
assign Zsaiw6 = (Gtaiw6 & Ntaiw6);
assign Ntaiw6 = (~(Utaiw6 | A0j7z6[18]));
assign Utaiw6 = (A0j7z6[19] | A0j7z6[1]);
assign Gtaiw6 = (~(Buaiw6 | A0j7z6[15]));
assign Buaiw6 = (A0j7z6[16] | A0j7z6[17]);
assign Ssaiw6 = (Iuaiw6 & Puaiw6);
assign Puaiw6 = (~(Wuaiw6 | A0j7z6[12]));
assign Wuaiw6 = (A0j7z6[13] | A0j7z6[14]);
assign Iuaiw6 = (~(A0j7z6[10] | A0j7z6[11]));
assign Slaiw6 = (Dvaiw6 & Kvaiw6);
assign Kvaiw6 = (Rvaiw6 & Zlaiw6);
assign Zlaiw6 = (~(Yvaiw6 & Doaiw6));
assign Yvaiw6 = (L28iw6 & Q22nv6);
assign Q22nv6 = (~(Fwaiw6 & Mwaiw6));
assign Mwaiw6 = (Ie5iw6 & Dv3iw6);
assign Fwaiw6 = (Twaiw6 & Nq6iw6);
assign Rvaiw6 = (~(Axaiw6 & Hxaiw6));
assign Hxaiw6 = (As67z6 | Cndet6);
assign Dvaiw6 = (A8cet6 & Ldo7v6);
assign Rkc8v6 = (Oxaiw6 | AUXFAULT[31]);
assign Oxaiw6 = (Bwi7z6[31] & Vxaiw6);
assign Vxaiw6 = (~(Cyaiw6 & X0hov6));
assign Kkc8v6 = (Jyaiw6 | AUXFAULT[30]);
assign Jyaiw6 = (Bwi7z6[30] & Qyaiw6);
assign Qyaiw6 = (~(Cyaiw6 & Ro3iw6));
assign Dkc8v6 = (Xyaiw6 | AUXFAULT[29]);
assign Xyaiw6 = (Bwi7z6[29] & Ezaiw6);
assign Ezaiw6 = (~(Cyaiw6 & Zz3iw6));
assign Wjc8v6 = (Lzaiw6 | AUXFAULT[28]);
assign Lzaiw6 = (Bwi7z6[28] & Szaiw6);
assign Szaiw6 = (~(Cyaiw6 & W14iw6));
assign Pjc8v6 = (Zzaiw6 | AUXFAULT[27]);
assign Zzaiw6 = (Bwi7z6[27] & G0biw6);
assign G0biw6 = (~(Cyaiw6 & H44iw6));
assign Ijc8v6 = (N0biw6 | AUXFAULT[26]);
assign N0biw6 = (Bwi7z6[26] & U0biw6);
assign U0biw6 = (~(Cyaiw6 & E64iw6));
assign Bjc8v6 = (B1biw6 | AUXFAULT[25]);
assign B1biw6 = (Bwi7z6[25] & I1biw6);
assign I1biw6 = (~(Cyaiw6 & Iklov6));
assign Uic8v6 = (P1biw6 | AUXFAULT[24]);
assign P1biw6 = (Bwi7z6[24] & W1biw6);
assign W1biw6 = (~(Cyaiw6 & Wf4iw6));
assign Cyaiw6 = (~(D2biw6 | Dv3iw6));
assign Nic8v6 = (K2biw6 | AUXFAULT[23]);
assign K2biw6 = (Bwi7z6[23] & R2biw6);
assign R2biw6 = (~(Y2biw6 & Cx4iw6));
assign Gic8v6 = (F3biw6 | AUXFAULT[22]);
assign F3biw6 = (Bwi7z6[22] & M3biw6);
assign M3biw6 = (~(Y2biw6 & D85iw6));
assign Zhc8v6 = (T3biw6 | AUXFAULT[21]);
assign T3biw6 = (Bwi7z6[21] & A4biw6);
assign A4biw6 = (~(Y2biw6 & Ej5iw6));
assign Shc8v6 = (H4biw6 | AUXFAULT[20]);
assign H4biw6 = (Bwi7z6[20] & O4biw6);
assign O4biw6 = (~(Y2biw6 & Bl5iw6));
assign Lhc8v6 = (V4biw6 | AUXFAULT[19]);
assign V4biw6 = (Bwi7z6[19] & C5biw6);
assign C5biw6 = (~(Y2biw6 & Mn5iw6));
assign Ehc8v6 = (J5biw6 | AUXFAULT[18]);
assign J5biw6 = (Bwi7z6[18] & Q5biw6);
assign Q5biw6 = (~(Y2biw6 & Jp5iw6));
assign Xgc8v6 = (X5biw6 | AUXFAULT[17]);
assign X5biw6 = (Bwi7z6[17] & E6biw6);
assign E6biw6 = (~(Y2biw6 & Gr5iw6));
assign Qgc8v6 = (L6biw6 | AUXFAULT[16]);
assign L6biw6 = (Bwi7z6[16] & S6biw6);
assign S6biw6 = (~(Y2biw6 & Is5iw6));
assign Y2biw6 = (~(D2biw6 | Ie5iw6));
assign Jgc8v6 = (Z6biw6 | AUXFAULT[15]);
assign Z6biw6 = (Bwi7z6[15] & G7biw6);
assign G7biw6 = (~(N7biw6 & Z0iov6));
assign Cgc8v6 = (U7biw6 | AUXFAULT[14]);
assign U7biw6 = (Bwi7z6[14] & B8biw6);
assign B8biw6 = (~(N7biw6 & Bk6iw6));
assign Vfc8v6 = (I8biw6 | AUXFAULT[13]);
assign I8biw6 = (Bwi7z6[13] & P8biw6);
assign P8biw6 = (~(N7biw6 & Guhov6));
assign Ofc8v6 = (W8biw6 | AUXFAULT[12]);
assign W8biw6 = (Bwi7z6[12] & D9biw6);
assign D9biw6 = (~(N7biw6 & Emhov6));
assign Hfc8v6 = (K9biw6 | AUXFAULT[11]);
assign K9biw6 = (Bwi7z6[11] & R9biw6);
assign R9biw6 = (~(N7biw6 & Dz6iw6));
assign Afc8v6 = (Y9biw6 | AUXFAULT[10]);
assign Y9biw6 = (Bwi7z6[10] & Fabiw6);
assign Fabiw6 = (~(N7biw6 & H17iw6));
assign Tec8v6 = (Mabiw6 | AUXFAULT[9]);
assign Mabiw6 = (Bwi7z6[9] & Tabiw6);
assign Tabiw6 = (~(N7biw6 & J27iw6));
assign Mec8v6 = (Abbiw6 | AUXFAULT[8]);
assign Abbiw6 = (Bwi7z6[8] & Hbbiw6);
assign Hbbiw6 = (~(N7biw6 & U47iw6));
assign N7biw6 = (Obbiw6 & Bqi7z6[1]);
assign Obbiw6 = (!D2biw6);
assign Fec8v6 = (Vbbiw6 | AUXFAULT[7]);
assign Vbbiw6 = (Bwi7z6[7] & Ccbiw6);
assign Ccbiw6 = (~(Jcbiw6 & R62nv6));
assign Ydc8v6 = (Qcbiw6 | AUXFAULT[6]);
assign Qcbiw6 = (Bwi7z6[6] & Xcbiw6);
assign Xcbiw6 = (~(Jcbiw6 & K62nv6));
assign Rdc8v6 = (Edbiw6 | AUXFAULT[5]);
assign Edbiw6 = (Bwi7z6[5] & Ldbiw6);
assign Ldbiw6 = (~(Jcbiw6 & D62nv6));
assign Kdc8v6 = (Sdbiw6 | AUXFAULT[4]);
assign Sdbiw6 = (Bwi7z6[4] & Zdbiw6);
assign Zdbiw6 = (~(Jcbiw6 & W52nv6));
assign Ddc8v6 = (Gebiw6 | AUXFAULT[3]);
assign Gebiw6 = (Bwi7z6[3] & Nebiw6);
assign Nebiw6 = (~(Jcbiw6 & P52nv6));
assign Wcc8v6 = (Uebiw6 | AUXFAULT[2]);
assign Uebiw6 = (Bwi7z6[2] & Bfbiw6);
assign Bfbiw6 = (~(Jcbiw6 & I52nv6));
assign Pcc8v6 = (Ifbiw6 | AUXFAULT[1]);
assign Ifbiw6 = (Bwi7z6[1] & Pfbiw6);
assign Pfbiw6 = (~(Jcbiw6 & B52nv6));
assign Icc8v6 = (Wfbiw6 | AUXFAULT[0]);
assign Wfbiw6 = (Bwi7z6[0] & Dgbiw6);
assign Dgbiw6 = (~(Jcbiw6 & U42nv6));
assign Jcbiw6 = (~(D2biw6 | Twaiw6));
assign D2biw6 = (~(Kgbiw6 & L28iw6));
assign Bcc8v6 = (Rgbiw6 ? U42nv6 : Dri7z6[0]);
assign Ubc8v6 = (Rgbiw6 ? B52nv6 : Dri7z6[1]);
assign Nbc8v6 = (Rgbiw6 ? I52nv6 : Dri7z6[2]);
assign Gbc8v6 = (Rgbiw6 ? P52nv6 : Dri7z6[3]);
assign Zac8v6 = (Rgbiw6 ? W52nv6 : Dri7z6[4]);
assign Sac8v6 = (Rgbiw6 ? D62nv6 : Dri7z6[5]);
assign Lac8v6 = (Rgbiw6 ? K62nv6 : Dri7z6[6]);
assign Eac8v6 = (Rgbiw6 ? R62nv6 : Dri7z6[7]);
assign Rgbiw6 = (~(Kg4iw6 | Twaiw6));
assign Kg4iw6 = (~(Ygbiw6 & Toi7z6[3]));
assign Ygbiw6 = (~(N92iw6 | Toi7z6[2]));
assign X9c8v6 = (Fhbiw6 ? U42nv6 : Rbk7z6[0]);
assign Q9c8v6 = (Mhbiw6 ? U42nv6 : Zlk7z6[0]);
assign J9c8v6 = (Thbiw6 ? U42nv6 : Hwk7z6[0]);
assign C9c8v6 = (Aibiw6 ? U42nv6 : P6l7z6[0]);
assign V8c8v6 = (Hibiw6 ? U42nv6 : Xgl7z6[0]);
assign O8c8v6 = (Oibiw6 ? U42nv6 : Frl7z6[0]);
assign H8c8v6 = (Vibiw6 ? U42nv6 : N1m7z6[0]);
assign A8c8v6 = (Cjbiw6 ? U42nv6 : Vbm7z6[0]);
assign T7c8v6 = (Fhbiw6 ? B52nv6 : Rbk7z6[1]);
assign M7c8v6 = (Mhbiw6 ? B52nv6 : Zlk7z6[1]);
assign F7c8v6 = (Thbiw6 ? B52nv6 : Hwk7z6[1]);
assign Y6c8v6 = (Aibiw6 ? B52nv6 : P6l7z6[1]);
assign R6c8v6 = (Hibiw6 ? B52nv6 : Xgl7z6[1]);
assign K6c8v6 = (Oibiw6 ? B52nv6 : Frl7z6[1]);
assign D6c8v6 = (Vibiw6 ? B52nv6 : N1m7z6[1]);
assign W5c8v6 = (Cjbiw6 ? B52nv6 : Vbm7z6[1]);
assign P5c8v6 = (Fhbiw6 ? I52nv6 : Rbk7z6[2]);
assign I5c8v6 = (Mhbiw6 ? I52nv6 : Zlk7z6[2]);
assign B5c8v6 = (Thbiw6 ? I52nv6 : Hwk7z6[2]);
assign U4c8v6 = (Aibiw6 ? I52nv6 : P6l7z6[2]);
assign N4c8v6 = (Hibiw6 ? I52nv6 : Xgl7z6[2]);
assign G4c8v6 = (Oibiw6 ? I52nv6 : Frl7z6[2]);
assign Z3c8v6 = (Vibiw6 ? I52nv6 : N1m7z6[2]);
assign S3c8v6 = (Cjbiw6 ? I52nv6 : Vbm7z6[2]);
assign L3c8v6 = (Fhbiw6 ? P52nv6 : Rbk7z6[3]);
assign E3c8v6 = (Mhbiw6 ? P52nv6 : Zlk7z6[3]);
assign X2c8v6 = (Thbiw6 ? P52nv6 : Hwk7z6[3]);
assign Q2c8v6 = (Aibiw6 ? P52nv6 : P6l7z6[3]);
assign J2c8v6 = (Hibiw6 ? P52nv6 : Xgl7z6[3]);
assign C2c8v6 = (Oibiw6 ? P52nv6 : Frl7z6[3]);
assign V1c8v6 = (Vibiw6 ? P52nv6 : N1m7z6[3]);
assign O1c8v6 = (Cjbiw6 ? P52nv6 : Vbm7z6[3]);
assign H1c8v6 = (Fhbiw6 ? W52nv6 : Rbk7z6[4]);
assign A1c8v6 = (Mhbiw6 ? W52nv6 : Zlk7z6[4]);
assign T0c8v6 = (Thbiw6 ? W52nv6 : Hwk7z6[4]);
assign M0c8v6 = (Aibiw6 ? W52nv6 : P6l7z6[4]);
assign F0c8v6 = (Hibiw6 ? W52nv6 : Xgl7z6[4]);
assign Yzb8v6 = (Oibiw6 ? W52nv6 : Frl7z6[4]);
assign Rzb8v6 = (Vibiw6 ? W52nv6 : N1m7z6[4]);
assign Kzb8v6 = (Cjbiw6 ? W52nv6 : Vbm7z6[4]);
assign Dzb8v6 = (Fhbiw6 ? D62nv6 : Rbk7z6[5]);
assign Fhbiw6 = (Jjbiw6 & Qjbiw6);
assign Wyb8v6 = (Xjbiw6 ? D62nv6 : Dfk7z6[5]);
assign Pyb8v6 = (Mhbiw6 ? D62nv6 : Zlk7z6[5]);
assign Mhbiw6 = (Jjbiw6 & Ekbiw6);
assign Iyb8v6 = (Lkbiw6 ? D62nv6 : Lpk7z6[5]);
assign Byb8v6 = (Thbiw6 ? D62nv6 : Hwk7z6[5]);
assign Thbiw6 = (Jjbiw6 & Skbiw6);
assign Uxb8v6 = (Zkbiw6 ? D62nv6 : Tzk7z6[5]);
assign Nxb8v6 = (Aibiw6 ? D62nv6 : P6l7z6[5]);
assign Aibiw6 = (Jjbiw6 & Glbiw6);
assign Gxb8v6 = (Nlbiw6 ? D62nv6 : Bal7z6[5]);
assign Zwb8v6 = (Hibiw6 ? D62nv6 : Xgl7z6[5]);
assign Hibiw6 = (Jjbiw6 & Ulbiw6);
assign Swb8v6 = (Bmbiw6 ? D62nv6 : Jkl7z6[5]);
assign Lwb8v6 = (Oibiw6 ? D62nv6 : Frl7z6[5]);
assign Oibiw6 = (Jjbiw6 & Imbiw6);
assign Ewb8v6 = (Pmbiw6 ? D62nv6 : Rul7z6[5]);
assign Xvb8v6 = (Vibiw6 ? D62nv6 : N1m7z6[5]);
assign Vibiw6 = (Jjbiw6 & Wmbiw6);
assign Qvb8v6 = (Dnbiw6 ? D62nv6 : Z4m7z6[5]);
assign Jvb8v6 = (Cjbiw6 ? D62nv6 : Vbm7z6[5]);
assign Cjbiw6 = (Jjbiw6 & Knbiw6);
assign Jjbiw6 = (Hc3iw6 & Rnbiw6);
assign Cvb8v6 = (Ynbiw6 ? D62nv6 : Hfm7z6[5]);
assign Vub8v6 = (Xjbiw6 ? K62nv6 : Dfk7z6[6]);
assign Oub8v6 = (Lkbiw6 ? K62nv6 : Fobiw6);
assign Hub8v6 = (Zkbiw6 ? K62nv6 : Mobiw6);
assign Aub8v6 = (Nlbiw6 ? K62nv6 : Tobiw6);
assign Ttb8v6 = (Bmbiw6 ? K62nv6 : Jkl7z6[6]);
assign Mtb8v6 = (Pmbiw6 ? K62nv6 : Apbiw6);
assign Ftb8v6 = (Dnbiw6 ? K62nv6 : Hpbiw6);
assign Ysb8v6 = (Ynbiw6 ? K62nv6 : Opbiw6);
assign Rsb8v6 = (Xjbiw6 ? R62nv6 : Dfk7z6[7]);
assign Xjbiw6 = (~(Vpbiw6 | Cqbiw6));
assign Ksb8v6 = (Lkbiw6 ? R62nv6 : Jqbiw6);
assign Lkbiw6 = (~(Vpbiw6 | Qqbiw6));
assign Dsb8v6 = (Zkbiw6 ? R62nv6 : Xqbiw6);
assign Zkbiw6 = (~(Vpbiw6 | Erbiw6));
assign Wrb8v6 = (Nlbiw6 ? R62nv6 : Lrbiw6);
assign Nlbiw6 = (~(Vpbiw6 | Srbiw6));
assign Prb8v6 = (Bmbiw6 ? R62nv6 : Jkl7z6[7]);
assign Bmbiw6 = (~(Vpbiw6 | Zrbiw6));
assign Irb8v6 = (Pmbiw6 ? R62nv6 : Gsbiw6);
assign Pmbiw6 = (Nsbiw6 & Imbiw6);
assign Brb8v6 = (Dnbiw6 ? R62nv6 : Usbiw6);
assign Dnbiw6 = (Nsbiw6 & Wmbiw6);
assign Nsbiw6 = (!Vpbiw6);
assign Uqb8v6 = (Ynbiw6 ? R62nv6 : Btbiw6);
assign Ynbiw6 = (~(Vpbiw6 | Itbiw6));
assign Vpbiw6 = (~(Hc3iw6 & Ptbiw6));
assign Nqb8v6 = (Wtbiw6 ? Rbk7z6[6] : U47iw6);
assign Gqb8v6 = (Dubiw6 ? Dfk7z6[8] : U47iw6);
assign Zpb8v6 = (Kubiw6 ? Zlk7z6[6] : U47iw6);
assign Spb8v6 = (Rubiw6 ? Lpk7z6[8] : U47iw6);
assign Lpb8v6 = (Yubiw6 ? Hwk7z6[6] : U47iw6);
assign Epb8v6 = (Fvbiw6 ? Tzk7z6[8] : U47iw6);
assign Xob8v6 = (Mvbiw6 ? P6l7z6[6] : U47iw6);
assign Qob8v6 = (Tvbiw6 ? Bal7z6[8] : U47iw6);
assign Job8v6 = (Awbiw6 ? Xgl7z6[6] : U47iw6);
assign Cob8v6 = (Hwbiw6 ? Jkl7z6[8] : U47iw6);
assign Vnb8v6 = (Owbiw6 ? Frl7z6[6] : U47iw6);
assign Onb8v6 = (Vwbiw6 ? Rul7z6[8] : U47iw6);
assign Hnb8v6 = (Cxbiw6 ? N1m7z6[6] : U47iw6);
assign Anb8v6 = (Jxbiw6 ? Z4m7z6[8] : U47iw6);
assign Tmb8v6 = (Qxbiw6 ? U47iw6 : Vbm7z6[6]);
assign Mmb8v6 = (Xxbiw6 ? U47iw6 : Hfm7z6[8]);
assign Fmb8v6 = (Wtbiw6 ? Rbk7z6[7] : J27iw6);
assign Ylb8v6 = (Dubiw6 ? Dfk7z6[9] : J27iw6);
assign Rlb8v6 = (Kubiw6 ? Zlk7z6[7] : J27iw6);
assign Klb8v6 = (Rubiw6 ? Eybiw6 : J27iw6);
assign Dlb8v6 = (Yubiw6 ? Hwk7z6[7] : J27iw6);
assign Wkb8v6 = (Fvbiw6 ? Lybiw6 : J27iw6);
assign Pkb8v6 = (Mvbiw6 ? P6l7z6[7] : J27iw6);
assign Ikb8v6 = (Tvbiw6 ? Sybiw6 : J27iw6);
assign Bkb8v6 = (Awbiw6 ? Xgl7z6[7] : J27iw6);
assign Ujb8v6 = (Hwbiw6 ? Jkl7z6[9] : J27iw6);
assign Njb8v6 = (Owbiw6 ? Frl7z6[7] : J27iw6);
assign Gjb8v6 = (Vwbiw6 ? Zybiw6 : J27iw6);
assign Zib8v6 = (Cxbiw6 ? N1m7z6[7] : J27iw6);
assign Sib8v6 = (Jxbiw6 ? Gzbiw6 : J27iw6);
assign Lib8v6 = (Qxbiw6 ? J27iw6 : Vbm7z6[7]);
assign Eib8v6 = (Xxbiw6 ? J27iw6 : Nzbiw6);
assign Xhb8v6 = (Wtbiw6 ? Rbk7z6[8] : H17iw6);
assign Qhb8v6 = (Dubiw6 ? Dfk7z6[10] : H17iw6);
assign Jhb8v6 = (Kubiw6 ? Zlk7z6[8] : H17iw6);
assign Chb8v6 = (Rubiw6 ? Uzbiw6 : H17iw6);
assign Vgb8v6 = (Yubiw6 ? Hwk7z6[8] : H17iw6);
assign Ogb8v6 = (Fvbiw6 ? B0ciw6 : H17iw6);
assign Hgb8v6 = (Mvbiw6 ? P6l7z6[8] : H17iw6);
assign Agb8v6 = (Tvbiw6 ? I0ciw6 : H17iw6);
assign Tfb8v6 = (Awbiw6 ? Xgl7z6[8] : H17iw6);
assign Mfb8v6 = (Hwbiw6 ? Jkl7z6[10] : H17iw6);
assign Ffb8v6 = (Owbiw6 ? Frl7z6[8] : H17iw6);
assign Yeb8v6 = (Vwbiw6 ? P0ciw6 : H17iw6);
assign Reb8v6 = (Cxbiw6 ? N1m7z6[8] : H17iw6);
assign Keb8v6 = (Jxbiw6 ? W0ciw6 : H17iw6);
assign Deb8v6 = (Qxbiw6 ? H17iw6 : Vbm7z6[8]);
assign Wdb8v6 = (Xxbiw6 ? H17iw6 : D1ciw6);
assign Pdb8v6 = (Wtbiw6 ? Rbk7z6[9] : Dz6iw6);
assign Wtbiw6 = (!K1ciw6);
assign Idb8v6 = (Dubiw6 ? Dfk7z6[11] : Dz6iw6);
assign Bdb8v6 = (Kubiw6 ? Zlk7z6[9] : Dz6iw6);
assign Kubiw6 = (!R1ciw6);
assign Ucb8v6 = (Rubiw6 ? Y1ciw6 : Dz6iw6);
assign Ncb8v6 = (Yubiw6 ? Hwk7z6[9] : Dz6iw6);
assign Yubiw6 = (!F2ciw6);
assign Gcb8v6 = (Fvbiw6 ? M2ciw6 : Dz6iw6);
assign Zbb8v6 = (Mvbiw6 ? P6l7z6[9] : Dz6iw6);
assign Mvbiw6 = (!T2ciw6);
assign Sbb8v6 = (Tvbiw6 ? A3ciw6 : Dz6iw6);
assign Lbb8v6 = (Awbiw6 ? Xgl7z6[9] : Dz6iw6);
assign Awbiw6 = (!H3ciw6);
assign Ebb8v6 = (Hwbiw6 ? Jkl7z6[11] : Dz6iw6);
assign Xab8v6 = (Owbiw6 ? Frl7z6[9] : Dz6iw6);
assign Owbiw6 = (!O3ciw6);
assign Qab8v6 = (Vwbiw6 ? V3ciw6 : Dz6iw6);
assign Vwbiw6 = (!C4ciw6);
assign Jab8v6 = (Cxbiw6 ? N1m7z6[9] : Dz6iw6);
assign Cxbiw6 = (!J4ciw6);
assign Cab8v6 = (Jxbiw6 ? Q4ciw6 : Dz6iw6);
assign V9b8v6 = (Qxbiw6 ? Dz6iw6 : Vbm7z6[9]);
assign O9b8v6 = (Xxbiw6 ? Dz6iw6 : X4ciw6);
assign H9b8v6 = (K1ciw6 ? Emhov6 : Rbk7z6[10]);
assign A9b8v6 = (E5ciw6 ? Emhov6 : Dfk7z6[12]);
assign T8b8v6 = (R1ciw6 ? Emhov6 : Zlk7z6[10]);
assign M8b8v6 = (S5ciw6 ? Emhov6 : L5ciw6);
assign F8b8v6 = (F2ciw6 ? Emhov6 : Hwk7z6[10]);
assign Y7b8v6 = (G6ciw6 ? Emhov6 : Z5ciw6);
assign R7b8v6 = (T2ciw6 ? Emhov6 : P6l7z6[10]);
assign K7b8v6 = (U6ciw6 ? Emhov6 : N6ciw6);
assign D7b8v6 = (H3ciw6 ? Emhov6 : Xgl7z6[10]);
assign W6b8v6 = (B7ciw6 ? Emhov6 : Jkl7z6[12]);
assign P6b8v6 = (O3ciw6 ? Emhov6 : Frl7z6[10]);
assign I6b8v6 = (C4ciw6 ? Emhov6 : I7ciw6);
assign B6b8v6 = (J4ciw6 ? Emhov6 : N1m7z6[10]);
assign U5b8v6 = (W7ciw6 ? Emhov6 : P7ciw6);
assign N5b8v6 = (Qxbiw6 ? Emhov6 : Vbm7z6[10]);
assign G5b8v6 = (Xxbiw6 ? Emhov6 : D8ciw6);
assign Z4b8v6 = (K1ciw6 ? Guhov6 : Rbk7z6[11]);
assign S4b8v6 = (E5ciw6 ? Guhov6 : Dfk7z6[13]);
assign L4b8v6 = (R1ciw6 ? Guhov6 : Zlk7z6[11]);
assign E4b8v6 = (S5ciw6 ? Guhov6 : K8ciw6);
assign X3b8v6 = (F2ciw6 ? Guhov6 : Hwk7z6[11]);
assign Q3b8v6 = (G6ciw6 ? Guhov6 : R8ciw6);
assign J3b8v6 = (T2ciw6 ? Guhov6 : P6l7z6[11]);
assign C3b8v6 = (U6ciw6 ? Guhov6 : Y8ciw6);
assign V2b8v6 = (H3ciw6 ? Guhov6 : Xgl7z6[11]);
assign O2b8v6 = (B7ciw6 ? Guhov6 : Jkl7z6[13]);
assign H2b8v6 = (O3ciw6 ? Guhov6 : Frl7z6[11]);
assign A2b8v6 = (C4ciw6 ? Guhov6 : F9ciw6);
assign T1b8v6 = (J4ciw6 ? Guhov6 : N1m7z6[11]);
assign M1b8v6 = (W7ciw6 ? Guhov6 : M9ciw6);
assign F1b8v6 = (Qxbiw6 ? Guhov6 : Vbm7z6[11]);
assign Y0b8v6 = (Xxbiw6 ? Guhov6 : T9ciw6);
assign R0b8v6 = (K1ciw6 ? Bk6iw6 : Rbk7z6[12]);
assign K0b8v6 = (E5ciw6 ? Bk6iw6 : Dfk7z6[14]);
assign D0b8v6 = (R1ciw6 ? Bk6iw6 : Zlk7z6[12]);
assign Wza8v6 = (S5ciw6 ? Bk6iw6 : Aaciw6);
assign Pza8v6 = (F2ciw6 ? Bk6iw6 : Hwk7z6[12]);
assign Iza8v6 = (G6ciw6 ? Bk6iw6 : Haciw6);
assign Bza8v6 = (T2ciw6 ? Bk6iw6 : P6l7z6[12]);
assign Uya8v6 = (U6ciw6 ? Bk6iw6 : Oaciw6);
assign Nya8v6 = (H3ciw6 ? Bk6iw6 : Xgl7z6[12]);
assign Gya8v6 = (B7ciw6 ? Bk6iw6 : Jkl7z6[14]);
assign Zxa8v6 = (O3ciw6 ? Bk6iw6 : Frl7z6[12]);
assign Sxa8v6 = (C4ciw6 ? Bk6iw6 : Vaciw6);
assign Lxa8v6 = (J4ciw6 ? Bk6iw6 : N1m7z6[12]);
assign Exa8v6 = (W7ciw6 ? Bk6iw6 : Cbciw6);
assign Xwa8v6 = (Qxbiw6 ? Bk6iw6 : Vbm7z6[12]);
assign Qwa8v6 = (Xxbiw6 ? Bk6iw6 : Jbciw6);
assign Jwa8v6 = (K1ciw6 ? Z0iov6 : Rbk7z6[13]);
assign K1ciw6 = (~(Qbciw6 | Cqbiw6));
assign Cwa8v6 = (E5ciw6 ? Z0iov6 : Dfk7z6[15]);
assign Vva8v6 = (R1ciw6 ? Z0iov6 : Zlk7z6[13]);
assign R1ciw6 = (~(Qbciw6 | Qqbiw6));
assign Ova8v6 = (S5ciw6 ? Z0iov6 : Xbciw6);
assign Hva8v6 = (F2ciw6 ? Z0iov6 : Hwk7z6[13]);
assign F2ciw6 = (~(Qbciw6 | Erbiw6));
assign Ava8v6 = (G6ciw6 ? Z0iov6 : Ecciw6);
assign Tua8v6 = (T2ciw6 ? Z0iov6 : P6l7z6[13]);
assign T2ciw6 = (~(Qbciw6 | Srbiw6));
assign Mua8v6 = (U6ciw6 ? Z0iov6 : Lcciw6);
assign Fua8v6 = (H3ciw6 ? Z0iov6 : Xgl7z6[13]);
assign H3ciw6 = (~(Qbciw6 | Zrbiw6));
assign Yta8v6 = (B7ciw6 ? Z0iov6 : Jkl7z6[15]);
assign Rta8v6 = (O3ciw6 ? Z0iov6 : Frl7z6[13]);
assign O3ciw6 = (~(Qbciw6 | Scciw6));
assign Kta8v6 = (C4ciw6 ? Z0iov6 : Zcciw6);
assign Dta8v6 = (J4ciw6 ? Z0iov6 : N1m7z6[13]);
assign J4ciw6 = (~(Qbciw6 | Gdciw6));
assign Wsa8v6 = (W7ciw6 ? Z0iov6 : Ndciw6);
assign Psa8v6 = (Qxbiw6 ? Z0iov6 : Vbm7z6[13]);
assign Qxbiw6 = (~(Qbciw6 | Itbiw6));
assign Qbciw6 = (~(Pvj7z6[1] & Rnbiw6));
assign Isa8v6 = (Xxbiw6 ? Z0iov6 : Udciw6);
assign Bsa8v6 = (Beciw6 ? Is5iw6 : Rbk7z6[14]);
assign Ura8v6 = (Dubiw6 ? Dfk7z6[16] : Is5iw6);
assign Nra8v6 = (Ieciw6 ? Is5iw6 : Zlk7z6[14]);
assign Gra8v6 = (Rubiw6 ? Lpk7z6[16] : Is5iw6);
assign Zqa8v6 = (Peciw6 ? Is5iw6 : Hwk7z6[14]);
assign Sqa8v6 = (Fvbiw6 ? Tzk7z6[16] : Is5iw6);
assign Lqa8v6 = (Weciw6 ? Is5iw6 : P6l7z6[14]);
assign Eqa8v6 = (Tvbiw6 ? Bal7z6[16] : Is5iw6);
assign Xpa8v6 = (Dfciw6 ? Is5iw6 : Xgl7z6[14]);
assign Qpa8v6 = (Hwbiw6 ? Jkl7z6[16] : Is5iw6);
assign Jpa8v6 = (Kfciw6 ? Is5iw6 : Frl7z6[14]);
assign Cpa8v6 = (C4ciw6 ? Is5iw6 : Rul7z6[16]);
assign Voa8v6 = (Rfciw6 ? Is5iw6 : N1m7z6[14]);
assign Ooa8v6 = (Jxbiw6 ? Z4m7z6[16] : Is5iw6);
assign Hoa8v6 = (Yfciw6 ? Is5iw6 : Vbm7z6[14]);
assign Aoa8v6 = (Fgciw6 ? Hfm7z6[16] : Is5iw6);
assign Tna8v6 = (Beciw6 ? Gr5iw6 : Rbk7z6[15]);
assign Mna8v6 = (Dubiw6 ? Dfk7z6[17] : Gr5iw6);
assign Fna8v6 = (Ieciw6 ? Gr5iw6 : Zlk7z6[15]);
assign Yma8v6 = (Rubiw6 ? Mgciw6 : Gr5iw6);
assign Rma8v6 = (Peciw6 ? Gr5iw6 : Hwk7z6[15]);
assign Kma8v6 = (Fvbiw6 ? Tgciw6 : Gr5iw6);
assign Dma8v6 = (Weciw6 ? Gr5iw6 : P6l7z6[15]);
assign Wla8v6 = (Tvbiw6 ? Ahciw6 : Gr5iw6);
assign Pla8v6 = (Dfciw6 ? Gr5iw6 : Xgl7z6[15]);
assign Ila8v6 = (Hwbiw6 ? Jkl7z6[17] : Gr5iw6);
assign Bla8v6 = (Kfciw6 ? Gr5iw6 : Frl7z6[15]);
assign Uka8v6 = (C4ciw6 ? Gr5iw6 : Hhciw6);
assign Nka8v6 = (Rfciw6 ? Gr5iw6 : N1m7z6[15]);
assign Gka8v6 = (Jxbiw6 ? Ohciw6 : Gr5iw6);
assign Zja8v6 = (Yfciw6 ? Gr5iw6 : Vbm7z6[15]);
assign Sja8v6 = (Fgciw6 ? Vhciw6 : Gr5iw6);
assign Fgciw6 = (!Xxbiw6);
assign Lja8v6 = (Beciw6 ? Jp5iw6 : Rbk7z6[16]);
assign Eja8v6 = (Dubiw6 ? Dfk7z6[18] : Jp5iw6);
assign Xia8v6 = (Ieciw6 ? Jp5iw6 : Zlk7z6[16]);
assign Qia8v6 = (Rubiw6 ? Ciciw6 : Jp5iw6);
assign Jia8v6 = (Peciw6 ? Jp5iw6 : Hwk7z6[16]);
assign Cia8v6 = (Fvbiw6 ? Jiciw6 : Jp5iw6);
assign Vha8v6 = (Weciw6 ? Jp5iw6 : P6l7z6[16]);
assign Oha8v6 = (Tvbiw6 ? Qiciw6 : Jp5iw6);
assign Hha8v6 = (Dfciw6 ? Jp5iw6 : Xgl7z6[16]);
assign Aha8v6 = (Hwbiw6 ? Jkl7z6[18] : Jp5iw6);
assign Tga8v6 = (Kfciw6 ? Jp5iw6 : Frl7z6[16]);
assign Mga8v6 = (C4ciw6 ? Jp5iw6 : Xiciw6);
assign Fga8v6 = (Rfciw6 ? Jp5iw6 : N1m7z6[16]);
assign Yfa8v6 = (Jxbiw6 ? Ejciw6 : Jp5iw6);
assign Rfa8v6 = (Yfciw6 ? Jp5iw6 : Vbm7z6[16]);
assign Kfa8v6 = (Xxbiw6 ? Jp5iw6 : Ljciw6);
assign Dfa8v6 = (Beciw6 ? Mn5iw6 : Rbk7z6[17]);
assign Wea8v6 = (Dubiw6 ? Dfk7z6[19] : Mn5iw6);
assign Dubiw6 = (!E5ciw6);
assign Pea8v6 = (Ieciw6 ? Mn5iw6 : Zlk7z6[17]);
assign Iea8v6 = (Rubiw6 ? Sjciw6 : Mn5iw6);
assign Rubiw6 = (!S5ciw6);
assign Bea8v6 = (Peciw6 ? Mn5iw6 : Hwk7z6[17]);
assign Uda8v6 = (Fvbiw6 ? Zjciw6 : Mn5iw6);
assign Fvbiw6 = (!G6ciw6);
assign Nda8v6 = (Weciw6 ? Mn5iw6 : P6l7z6[17]);
assign Gda8v6 = (Tvbiw6 ? Gkciw6 : Mn5iw6);
assign Tvbiw6 = (!U6ciw6);
assign Zca8v6 = (Dfciw6 ? Mn5iw6 : Xgl7z6[17]);
assign Sca8v6 = (Hwbiw6 ? Jkl7z6[19] : Mn5iw6);
assign Hwbiw6 = (!B7ciw6);
assign Lca8v6 = (Kfciw6 ? Mn5iw6 : Frl7z6[17]);
assign Eca8v6 = (C4ciw6 ? Mn5iw6 : Nkciw6);
assign Xba8v6 = (Rfciw6 ? Mn5iw6 : N1m7z6[17]);
assign Qba8v6 = (Jxbiw6 ? Ukciw6 : Mn5iw6);
assign Jxbiw6 = (!W7ciw6);
assign Jba8v6 = (Yfciw6 ? Mn5iw6 : Vbm7z6[17]);
assign Cba8v6 = (Xxbiw6 ? Mn5iw6 : Blciw6);
assign Vaa8v6 = (Beciw6 ? Bl5iw6 : Rbk7z6[18]);
assign Oaa8v6 = (E5ciw6 ? Bl5iw6 : Dfk7z6[20]);
assign Haa8v6 = (Ieciw6 ? Bl5iw6 : Zlk7z6[18]);
assign Aaa8v6 = (S5ciw6 ? Bl5iw6 : Ilciw6);
assign T9a8v6 = (Peciw6 ? Bl5iw6 : Hwk7z6[18]);
assign M9a8v6 = (G6ciw6 ? Bl5iw6 : Plciw6);
assign F9a8v6 = (Weciw6 ? Bl5iw6 : P6l7z6[18]);
assign Y8a8v6 = (U6ciw6 ? Bl5iw6 : Wlciw6);
assign R8a8v6 = (Dfciw6 ? Bl5iw6 : Xgl7z6[18]);
assign K8a8v6 = (B7ciw6 ? Bl5iw6 : Jkl7z6[20]);
assign D8a8v6 = (Kfciw6 ? Bl5iw6 : Frl7z6[18]);
assign W7a8v6 = (C4ciw6 ? Bl5iw6 : Dmciw6);
assign P7a8v6 = (Rfciw6 ? Bl5iw6 : N1m7z6[18]);
assign I7a8v6 = (W7ciw6 ? Bl5iw6 : Kmciw6);
assign B7a8v6 = (Yfciw6 ? Bl5iw6 : Vbm7z6[18]);
assign U6a8v6 = (Xxbiw6 ? Bl5iw6 : Rmciw6);
assign N6a8v6 = (Beciw6 ? Ej5iw6 : Rbk7z6[19]);
assign Beciw6 = (~(Ymciw6 | Cqbiw6));
assign G6a8v6 = (E5ciw6 ? Ej5iw6 : Dfk7z6[21]);
assign Z5a8v6 = (Ieciw6 ? Ej5iw6 : Zlk7z6[19]);
assign Ieciw6 = (~(Ymciw6 | Qqbiw6));
assign S5a8v6 = (S5ciw6 ? Ej5iw6 : Fnciw6);
assign L5a8v6 = (Peciw6 ? Ej5iw6 : Hwk7z6[19]);
assign Peciw6 = (~(Ymciw6 | Erbiw6));
assign E5a8v6 = (G6ciw6 ? Ej5iw6 : Mnciw6);
assign X4a8v6 = (Weciw6 ? Ej5iw6 : P6l7z6[19]);
assign Weciw6 = (~(Ymciw6 | Srbiw6));
assign Q4a8v6 = (U6ciw6 ? Ej5iw6 : Tnciw6);
assign J4a8v6 = (Dfciw6 ? Ej5iw6 : Xgl7z6[19]);
assign Dfciw6 = (~(Ymciw6 | Zrbiw6));
assign C4a8v6 = (B7ciw6 ? Ej5iw6 : Jkl7z6[21]);
assign V3a8v6 = (Kfciw6 ? Ej5iw6 : Frl7z6[19]);
assign Kfciw6 = (~(Ymciw6 | Scciw6));
assign O3a8v6 = (C4ciw6 ? Ej5iw6 : Aociw6);
assign H3a8v6 = (Rfciw6 ? Ej5iw6 : N1m7z6[19]);
assign Rfciw6 = (~(Ymciw6 | Gdciw6));
assign Ymciw6 = (!Hociw6);
assign A3a8v6 = (W7ciw6 ? Ej5iw6 : Oociw6);
assign T2a8v6 = (Yfciw6 ? Ej5iw6 : Vbm7z6[19]);
assign Yfciw6 = (Hociw6 & Knbiw6);
assign Hociw6 = (Pvj7z6[2] & Rnbiw6);
assign Rnbiw6 = (!Vociw6);
assign M2a8v6 = (Xxbiw6 ? Ej5iw6 : Cpciw6);
assign F2a8v6 = (E5ciw6 ? D85iw6 : Dfk7z6[22]);
assign Y1a8v6 = (S5ciw6 ? D85iw6 : Jpciw6);
assign R1a8v6 = (G6ciw6 ? D85iw6 : Qpciw6);
assign K1a8v6 = (U6ciw6 ? D85iw6 : Xpciw6);
assign D1a8v6 = (B7ciw6 ? D85iw6 : Jkl7z6[22]);
assign W0a8v6 = (C4ciw6 ? D85iw6 : Eqciw6);
assign P0a8v6 = (W7ciw6 ? D85iw6 : Lqciw6);
assign I0a8v6 = (Xxbiw6 ? D85iw6 : Sqciw6);
assign B0a8v6 = (E5ciw6 ? Cx4iw6 : Dfk7z6[23]);
assign E5ciw6 = (~(Zqciw6 | Cqbiw6));
assign Uz98v6 = (S5ciw6 ? Cx4iw6 : Grciw6);
assign S5ciw6 = (~(Zqciw6 | Qqbiw6));
assign Nz98v6 = (G6ciw6 ? Cx4iw6 : Nrciw6);
assign G6ciw6 = (~(Zqciw6 | Erbiw6));
assign Gz98v6 = (U6ciw6 ? Cx4iw6 : Urciw6);
assign U6ciw6 = (~(Zqciw6 | Srbiw6));
assign Zy98v6 = (B7ciw6 ? Cx4iw6 : Jkl7z6[23]);
assign B7ciw6 = (~(Zqciw6 | Zrbiw6));
assign Sy98v6 = (C4ciw6 ? Cx4iw6 : Bsciw6);
assign C4ciw6 = (~(Zqciw6 | Scciw6));
assign Scciw6 = (!Imbiw6);
assign Ly98v6 = (W7ciw6 ? Cx4iw6 : Isciw6);
assign W7ciw6 = (~(Zqciw6 | Gdciw6));
assign Ey98v6 = (Xxbiw6 ? Cx4iw6 : Psciw6);
assign Xxbiw6 = (~(Zqciw6 | Itbiw6));
assign Zqciw6 = (~(Ptbiw6 & Cd3iw6));
assign Xx98v6 = (Wsciw6 ? Wf4iw6 : Rbk7z6[20]);
assign Qx98v6 = (Dtciw6 ? Wf4iw6 : Dfk7z6[24]);
assign Jx98v6 = (Ktciw6 ? Wf4iw6 : Zlk7z6[20]);
assign Cx98v6 = (Rtciw6 ? Wf4iw6 : Lpk7z6[24]);
assign Vw98v6 = (Ytciw6 ? Wf4iw6 : Hwk7z6[20]);
assign Ow98v6 = (Fuciw6 ? Wf4iw6 : Tzk7z6[24]);
assign Hw98v6 = (Muciw6 ? Wf4iw6 : P6l7z6[20]);
assign Aw98v6 = (Tuciw6 ? Wf4iw6 : Bal7z6[24]);
assign Tv98v6 = (Avciw6 ? Wf4iw6 : Xgl7z6[20]);
assign Mv98v6 = (Hvciw6 ? Wf4iw6 : Jkl7z6[24]);
assign Fv98v6 = (Ovciw6 ? Wf4iw6 : Frl7z6[20]);
assign Yu98v6 = (Vvciw6 ? Wf4iw6 : Rul7z6[24]);
assign Ru98v6 = (Cwciw6 ? Wf4iw6 : N1m7z6[20]);
assign Ku98v6 = (Jwciw6 ? Wf4iw6 : Z4m7z6[24]);
assign Du98v6 = (Qwciw6 ? Wf4iw6 : Vbm7z6[20]);
assign Wt98v6 = (Pklov6 ? Wf4iw6 : Xwciw6);
assign Pt98v6 = (Wsciw6 ? Iklov6 : Rbk7z6[21]);
assign It98v6 = (Dtciw6 ? Iklov6 : Dfk7z6[25]);
assign Bt98v6 = (Ktciw6 ? Iklov6 : Zlk7z6[21]);
assign Us98v6 = (Rtciw6 ? Iklov6 : Exciw6);
assign Ns98v6 = (Ytciw6 ? Iklov6 : Hwk7z6[21]);
assign Gs98v6 = (Fuciw6 ? Iklov6 : Lxciw6);
assign Zr98v6 = (Muciw6 ? Iklov6 : P6l7z6[21]);
assign Sr98v6 = (Tuciw6 ? Iklov6 : Sxciw6);
assign Lr98v6 = (Avciw6 ? Iklov6 : Xgl7z6[21]);
assign Er98v6 = (Hvciw6 ? Iklov6 : Jkl7z6[25]);
assign Xq98v6 = (Ovciw6 ? Iklov6 : Frl7z6[21]);
assign Qq98v6 = (Vvciw6 ? Iklov6 : Zxciw6);
assign Jq98v6 = (Cwciw6 ? Iklov6 : N1m7z6[21]);
assign Cq98v6 = (Jwciw6 ? Iklov6 : Gyciw6);
assign Vp98v6 = (Qwciw6 ? Iklov6 : Vbm7z6[21]);
assign Op98v6 = (Wsciw6 ? E64iw6 : Rbk7z6[22]);
assign Hp98v6 = (Dtciw6 ? E64iw6 : Dfk7z6[26]);
assign Ap98v6 = (Ktciw6 ? E64iw6 : Zlk7z6[22]);
assign To98v6 = (Rtciw6 ? E64iw6 : Nyciw6);
assign Mo98v6 = (Ytciw6 ? E64iw6 : Hwk7z6[22]);
assign Fo98v6 = (Fuciw6 ? E64iw6 : Uyciw6);
assign Yn98v6 = (Muciw6 ? E64iw6 : P6l7z6[22]);
assign Rn98v6 = (Tuciw6 ? E64iw6 : Bzciw6);
assign Kn98v6 = (Avciw6 ? E64iw6 : Xgl7z6[22]);
assign Dn98v6 = (Hvciw6 ? E64iw6 : Jkl7z6[26]);
assign Wm98v6 = (Ovciw6 ? E64iw6 : Frl7z6[22]);
assign Pm98v6 = (Vvciw6 ? E64iw6 : Izciw6);
assign Im98v6 = (Cwciw6 ? E64iw6 : N1m7z6[22]);
assign Bm98v6 = (Jwciw6 ? E64iw6 : Pzciw6);
assign Ul98v6 = (Qwciw6 ? E64iw6 : Vbm7z6[22]);
assign Nl98v6 = (Pklov6 ? E64iw6 : Wzciw6);
assign Gl98v6 = (Dtciw6 ? H44iw6 : Dfk7z6[27]);
assign Zk98v6 = (Rtciw6 ? H44iw6 : D0diw6);
assign Sk98v6 = (Fuciw6 ? H44iw6 : K0diw6);
assign Lk98v6 = (Tuciw6 ? H44iw6 : R0diw6);
assign Ek98v6 = (Hvciw6 ? H44iw6 : Jkl7z6[27]);
assign Xj98v6 = (Vvciw6 ? H44iw6 : Y0diw6);
assign Qj98v6 = (Jwciw6 ? H44iw6 : F1diw6);
assign Jj98v6 = (Pklov6 ? H44iw6 : M1diw6);
assign Cj98v6 = (Wsciw6 ? W14iw6 : Rbk7z6[23]);
assign Wsciw6 = (T1diw6 & Qjbiw6);
assign Qjbiw6 = (!Cqbiw6);
assign Vi98v6 = (Dtciw6 ? W14iw6 : Dfk7z6[28]);
assign Oi98v6 = (Ktciw6 ? W14iw6 : Zlk7z6[23]);
assign Ktciw6 = (T1diw6 & Ekbiw6);
assign Ekbiw6 = (!Qqbiw6);
assign Hi98v6 = (Rtciw6 ? W14iw6 : A2diw6);
assign Ai98v6 = (Ytciw6 ? W14iw6 : Hwk7z6[23]);
assign Ytciw6 = (T1diw6 & Skbiw6);
assign Skbiw6 = (!Erbiw6);
assign Th98v6 = (Fuciw6 ? W14iw6 : H2diw6);
assign Mh98v6 = (Muciw6 ? W14iw6 : P6l7z6[23]);
assign Muciw6 = (T1diw6 & Glbiw6);
assign Glbiw6 = (!Srbiw6);
assign Fh98v6 = (Tuciw6 ? W14iw6 : O2diw6);
assign Yg98v6 = (Avciw6 ? W14iw6 : Xgl7z6[23]);
assign Avciw6 = (T1diw6 & Ulbiw6);
assign Ulbiw6 = (!Zrbiw6);
assign Rg98v6 = (Hvciw6 ? W14iw6 : Jkl7z6[28]);
assign Kg98v6 = (Ovciw6 ? W14iw6 : Frl7z6[23]);
assign Ovciw6 = (T1diw6 & Imbiw6);
assign Dg98v6 = (Vvciw6 ? W14iw6 : V2diw6);
assign Wf98v6 = (Cwciw6 ? W14iw6 : N1m7z6[23]);
assign Cwciw6 = (~(C3diw6 | Gdciw6));
assign Pf98v6 = (Jwciw6 ? W14iw6 : J3diw6);
assign If98v6 = (Qwciw6 ? W14iw6 : Vbm7z6[23]);
assign Qwciw6 = (T1diw6 & Knbiw6);
assign T1diw6 = (!C3diw6);
assign C3diw6 = (Vc3iw6 | Vociw6);
assign Bf98v6 = (Pklov6 ? W14iw6 : Q3diw6);
assign Ue98v6 = (Dtciw6 ? Zz3iw6 : Dfk7z6[29]);
assign Ne98v6 = (Rtciw6 ? Zz3iw6 : X3diw6);
assign Ge98v6 = (Fuciw6 ? Zz3iw6 : E4diw6);
assign Zd98v6 = (Tuciw6 ? Zz3iw6 : L4diw6);
assign Sd98v6 = (Hvciw6 ? Zz3iw6 : Jkl7z6[29]);
assign Ld98v6 = (Vvciw6 ? Zz3iw6 : S4diw6);
assign Ed98v6 = (Jwciw6 ? Zz3iw6 : Z4diw6);
assign Xc98v6 = (Pklov6 ? Zz3iw6 : G5diw6);
assign Qc98v6 = (Dtciw6 ? Ro3iw6 : Dfk7z6[30]);
assign Jc98v6 = (Rtciw6 ? Ro3iw6 : N5diw6);
assign Cc98v6 = (Fuciw6 ? Ro3iw6 : U5diw6);
assign Vb98v6 = (Tuciw6 ? Ro3iw6 : B6diw6);
assign Ob98v6 = (Hvciw6 ? Ro3iw6 : Jkl7z6[30]);
assign Hb98v6 = (Vvciw6 ? Ro3iw6 : I6diw6);
assign Ab98v6 = (Jwciw6 ? Ro3iw6 : P6diw6);
assign Ta98v6 = (Pklov6 ? Ro3iw6 : W6diw6);
assign Ma98v6 = (Dtciw6 ? X0hov6 : Dfk7z6[31]);
assign Dtciw6 = (~(D7diw6 | Cqbiw6));
assign Cqbiw6 = (K7diw6 & R7diw6);
assign R7diw6 = (~(K49iw6 & Y7diw6));
assign K49iw6 = (L19iw6 & Orhov6);
assign K7diw6 = (~(Hyj7z6[0] & F8diw6));
assign Fa98v6 = (Rtciw6 ? X0hov6 : M8diw6);
assign Rtciw6 = (~(D7diw6 | Qqbiw6));
assign Qqbiw6 = (T8diw6 & A9diw6);
assign A9diw6 = (~(H9diw6 & Y7diw6));
assign T8diw6 = (~(Hyj7z6[1] & F8diw6));
assign M8diw6 = (!Yk87z6);
assign Y998v6 = (Fuciw6 ? X0hov6 : O9diw6);
assign Fuciw6 = (~(D7diw6 | Erbiw6));
assign Erbiw6 = (V9diw6 & Cadiw6);
assign Cadiw6 = (~(I39iw6 & Y7diw6));
assign I39iw6 = (Orhov6 & B52nv6);
assign V9diw6 = (~(Hyj7z6[2] & F8diw6));
assign O9diw6 = (!Sr87z6);
assign R998v6 = (Tuciw6 ? X0hov6 : Jadiw6);
assign Tuciw6 = (~(D7diw6 | Srbiw6));
assign Srbiw6 = (Qadiw6 & Xadiw6);
assign Xadiw6 = (~(Y7diw6 & Ebdiw6));
assign Y7diw6 = (~(I52nv6 | F8diw6));
assign Qadiw6 = (~(Hyj7z6[3] & F8diw6));
assign K998v6 = (Hvciw6 ? X0hov6 : Jkl7z6[31]);
assign Hvciw6 = (~(D7diw6 | Zrbiw6));
assign Zrbiw6 = (Lbdiw6 & Sbdiw6);
assign Sbdiw6 = (Zbdiw6 | B52nv6);
assign Lbdiw6 = (~(Hyj7z6[4] & F8diw6));
assign D998v6 = (Vvciw6 ? X0hov6 : Gcdiw6);
assign Vvciw6 = (Ncdiw6 & Imbiw6);
assign Imbiw6 = (Bddiw6 ? Ucdiw6 : Hyj7z6[5]);
assign Gcdiw6 = (!Ee87z6);
assign W898v6 = (Jwciw6 ? X0hov6 : Iddiw6);
assign Jwciw6 = (Ncdiw6 & Wmbiw6);
assign Wmbiw6 = (!Gdciw6);
assign Gdciw6 = (Pddiw6 & Wddiw6);
assign Wddiw6 = (Zbdiw6 | L19iw6);
assign Zbdiw6 = (~(Dediw6 & Bddiw6));
assign Dediw6 = (Orhov6 & I52nv6);
assign Pddiw6 = (~(Hyj7z6[6] & F8diw6));
assign Iddiw6 = (!K787z6);
assign P898v6 = (Pklov6 ? X0hov6 : Kediw6);
assign Pklov6 = (Ncdiw6 & Knbiw6);
assign Knbiw6 = (!Itbiw6);
assign Itbiw6 = (Bddiw6 ? Vz8iw6 : C09iw6);
assign Bddiw6 = (!F8diw6);
assign Vz8iw6 = (~(Ebdiw6 & I52nv6));
assign Ncdiw6 = (!D7diw6);
assign D7diw6 = (Vc3iw6 | Rediw6);
assign Vc3iw6 = (~(Pvj7z6[3] & Cd3iw6));
assign Kediw6 = (!Iw77z6);
assign I898v6 = (~(Yediw6 & Senet6));
assign Yediw6 = (Ffdiw6 & Mfdiw6);
assign Ffdiw6 = (Tfdiw6 | Gr2et6);
assign B898v6 = (Agdiw6 & Hgdiw6);
assign Hgdiw6 = (Ogdiw6 & Cmm7z6[0]);
assign Ogdiw6 = (Lgonv6 & Xc4iw6);
assign Agdiw6 = (Vgdiw6 & Pbhnv6);
assign Vgdiw6 = (Wbhnv6 & Vfmov6);
assign U798v6 = (Chdiw6 ? Dzget6 : Hjqnv6);
assign N798v6 = (Chdiw6 ? Qwget6 : Lhmov6);
assign G798v6 = (Chdiw6 ? V5k7z6[6] : X0k7z6[6]);
assign Z698v6 = (Chdiw6 ? V5k7z6[7] : X0k7z6[7]);
assign S698v6 = (Chdiw6 ? V5k7z6[8] : X0k7z6[8]);
assign L698v6 = (Chdiw6 ? V5k7z6[9] : X0k7z6[9]);
assign E698v6 = (Chdiw6 ? V5k7z6[10] : X0k7z6[10]);
assign X598v6 = (Chdiw6 ? V5k7z6[11] : X0k7z6[11]);
assign Q598v6 = (Chdiw6 ? V5k7z6[12] : X0k7z6[12]);
assign J598v6 = (Chdiw6 ? V5k7z6[13] : X0k7z6[13]);
assign C598v6 = (Chdiw6 ? V5k7z6[14] : X0k7z6[14]);
assign V498v6 = (Chdiw6 ? V5k7z6[15] : X0k7z6[15]);
assign O498v6 = (Chdiw6 ? V5k7z6[16] : X0k7z6[16]);
assign H498v6 = (Chdiw6 ? Jhdiw6 : X0k7z6[17]);
assign A498v6 = (Chdiw6 ? V5k7z6[18] : X0k7z6[18]);
assign T398v6 = (Chdiw6 ? V5k7z6[19] : X0k7z6[19]);
assign M398v6 = (Chdiw6 ? Qhdiw6 : X0k7z6[20]);
assign Qhdiw6 = (!Cj77z6);
assign F398v6 = (Chdiw6 ? V5k7z6[21] : X0k7z6[21]);
assign Y298v6 = (Chdiw6 ? V5k7z6[22] : X0k7z6[22]);
assign R298v6 = (Chdiw6 ? Xhdiw6 : X0k7z6[23]);
assign Xhdiw6 = (!Kj77z6);
assign K298v6 = (Chdiw6 ? V5k7z6[24] : X0k7z6[24]);
assign D298v6 = (Chdiw6 ? V5k7z6[25] : X0k7z6[25]);
assign W198v6 = (Chdiw6 ? Eidiw6 : X0k7z6[26]);
assign Eidiw6 = (!U297z6);
assign P198v6 = (Chdiw6 ? V5k7z6[27] : X0k7z6[27]);
assign I198v6 = (Chdiw6 ? V5k7z6[28] : X0k7z6[28]);
assign B198v6 = (Chdiw6 ? V5k7z6[29] : X0k7z6[29]);
assign Chdiw6 = (!Obo7v6);
assign U098v6 = (Obo7v6 ? X0k7z6[30] : V5k7z6[30]);
assign N098v6 = (Obo7v6 ? X0k7z6[31] : V5k7z6[31]);
assign G098v6 = (Obo7v6 ? X0k7z6[5] : V5k7z6[5]);
assign Zz88v6 = (Lidiw6 ? P9i7z6[9] : G4i7z6[9]);
assign Sz88v6 = (Lidiw6 ? P9i7z6[8] : G4i7z6[8]);
assign Lz88v6 = (Lidiw6 ? P9i7z6[7] : G4i7z6[7]);
assign Ez88v6 = (Lidiw6 ? P9i7z6[6] : G4i7z6[6]);
assign Xy88v6 = (Lidiw6 ? P9i7z6[5] : G4i7z6[5]);
assign Qy88v6 = (Lidiw6 ? P9i7z6[4] : G4i7z6[4]);
assign Jy88v6 = (Lidiw6 ? P9i7z6[3] : G4i7z6[3]);
assign Cy88v6 = (Lidiw6 ? P9i7z6[2] : G4i7z6[2]);
assign Vx88v6 = (Lidiw6 ? P9i7z6[1] : G4i7z6[1]);
assign Ox88v6 = (Sidiw6 ? G4i7z6[0] : P9i7z6[0]);
assign Hx88v6 = (Zidiw6 ? Wbhnv6 : Bbp7z6[0]);
assign Ax88v6 = (Zidiw6 ? Anehw6 : Bbp7z6[1]);
assign Tw88v6 = (Zidiw6 ? Cmm7z6[0] : Ncp7z6[0]);
assign Mw88v6 = (Zidiw6 ? Cmm7z6[1] : Ncp7z6[1]);
assign Fw88v6 = (Zidiw6 ? Lhmov6 : L42ft6);
assign Yv88v6 = (K94iw6 ? Ea2ft6 : Gjdiw6);
assign Rv88v6 = (~(Njdiw6 & Ujdiw6));
assign Ujdiw6 = (~(Bkdiw6 & Gr2et6));
assign Njdiw6 = (~(Ikdiw6 | Tfdiw6));
assign Ikdiw6 = (Ihnet6 & Ypinv6);
assign Kv88v6 = (~(Pkdiw6 & Wkdiw6));
assign Wkdiw6 = (~(Dldiw6 & Kldiw6));
assign Dldiw6 = (!Rldiw6);
assign Pkdiw6 = (~(Xnh7z6[0] & P1jhw6));
assign Dv88v6 = (~(Yldiw6 & Fmdiw6));
assign Fmdiw6 = (Rldiw6 | Kldiw6);
assign Rldiw6 = (~(Mmdiw6 & B1jhw6));
assign Mmdiw6 = (T3cdt6 & B2jnv6);
assign Yldiw6 = (~(Xnh7z6[1] & P1jhw6));
assign Wu88v6 = (~(Tmdiw6 & Andiw6));
assign Andiw6 = (~(Hndiw6 & B1jhw6));
assign B1jhw6 = (Ondiw6 & Vndiw6);
assign Vndiw6 = (Codiw6 & Fsmov6);
assign Ondiw6 = (Jodiw6 & Ii9ov6);
assign Jodiw6 = (!P1jhw6);
assign Hndiw6 = (Qodiw6 & Xodiw6);
assign Tmdiw6 = (~(Xnh7z6[2] & P1jhw6));
assign P1jhw6 = (~(O5a7z6 & Epdiw6));
assign Epdiw6 = (~(Lpdiw6 & Spdiw6));
assign Lpdiw6 = (~(Zpdiw6 & Codiw6));
assign Codiw6 = (Aeonv6 & Lxydt6);
assign Pu88v6 = (~(Ygh7v6 & Uimov6));
assign Iu88v6 = (Uimov6 ? Y9pet6 : Hjqnv6);
assign Bu88v6 = (~(Gqdiw6 & Nqdiw6));
assign Nqdiw6 = (~(Uqdiw6 & Ezphw6));
assign Ezphw6 = (Brdiw6 & Irdiw6);
assign Irdiw6 = (Prdiw6 & Wrdiw6);
assign Wrdiw6 = (B2jnv6 & Lhmov6);
assign Prdiw6 = (Zblov6 & Yhqnv6);
assign Brdiw6 = (Dsdiw6 & Ghonv6);
assign Ghonv6 = (!Bionv6);
assign Bionv6 = (~(Ksdiw6 & Rsdiw6));
assign Ksdiw6 = (Aeonv6 & Vb4iw6);
assign Dsdiw6 = (Qodiw6 & Tlmov6);
assign Uqdiw6 = (Lzphw6 & Ysdiw6);
assign Lzphw6 = (~(Cyphw6 | Ftdiw6));
assign Ftdiw6 = (~(Rj9ov6 | Hm1ov6));
assign Gqdiw6 = (~(Dkm7z6[0] & Zzphw6));
assign Zzphw6 = (!Rsdiw6);
assign Ut88v6 = (~(Mtdiw6 & Ttdiw6));
assign Ttdiw6 = (Audiw6 | Alonv6);
assign Alonv6 = (Hudiw6 & Oudiw6);
assign Oudiw6 = (~(Vudiw6 & Cvdiw6));
assign Cvdiw6 = (!Jvdiw6);
assign Hudiw6 = (~(Enonv6 & Qvdiw6));
assign Mtdiw6 = (~(Dq9ov6 & Ven7z6[2]));
assign Nt88v6 = (~(Xvdiw6 & Ewdiw6));
assign Ewdiw6 = (Audiw6 | Tkonv6);
assign Tkonv6 = (Lwdiw6 & Swdiw6);
assign Swdiw6 = (~(Vudiw6 & Zwdiw6));
assign Lwdiw6 = (~(Gxdiw6 & Enonv6));
assign Gxdiw6 = (!Nxdiw6);
assign Audiw6 = (!Hl9ov6);
assign Xvdiw6 = (~(Dq9ov6 & Ven7z6[1]));
assign Gt88v6 = (~(Uxdiw6 & Bydiw6));
assign Bydiw6 = (~(Hl9ov6 & Mkonv6));
assign Mkonv6 = (~(Iydiw6 & Pydiw6));
assign Pydiw6 = (~(Wydiw6 & Enonv6));
assign Wydiw6 = (Cmm7z6[1] & Dzdiw6);
assign Dzdiw6 = (~(Cmm7z6[0] & Ta4iw6));
assign Iydiw6 = (~(Vudiw6 & Kzdiw6));
assign Kzdiw6 = (~(Rzdiw6 & Yzdiw6));
assign Yzdiw6 = (~(Hub7z6[0] & Stpnv6));
assign Uxdiw6 = (~(Dq9ov6 & Ven7z6[0]));
assign Zs88v6 = (F0eiw6 ? Icn7z6[0] : X9yet6);
assign Ss88v6 = (F0eiw6 ? Icn7z6[1] : Icyet6);
assign Ls88v6 = (F0eiw6 ? Icn7z6[2] : T2zet6);
assign Es88v6 = (F0eiw6 ? Icn7z6[3] : S0zet6);
assign Xr88v6 = (F0eiw6 ? Icn7z6[4] : Ryyet6);
assign Qr88v6 = (F0eiw6 ? Icn7z6[5] : Hjn7z6[5]);
assign Jr88v6 = (F0eiw6 ? Icn7z6[6] : Hjn7z6[6]);
assign Cr88v6 = (F0eiw6 ? Icn7z6[7] : Hjn7z6[7]);
assign Vq88v6 = (F0eiw6 ? Icn7z6[8] : Hjn7z6[8]);
assign Oq88v6 = (F0eiw6 ? Icn7z6[9] : Hjn7z6[9]);
assign Hq88v6 = (F0eiw6 ? Icn7z6[10] : Hjn7z6[10]);
assign Aq88v6 = (F0eiw6 ? Icn7z6[11] : Hjn7z6[11]);
assign Tp88v6 = (F0eiw6 ? Icn7z6[12] : Hjn7z6[12]);
assign Mp88v6 = (F0eiw6 ? Icn7z6[13] : Hjn7z6[13]);
assign Fp88v6 = (F0eiw6 ? Icn7z6[14] : Hjn7z6[14]);
assign Yo88v6 = (F0eiw6 ? Icn7z6[15] : Hjn7z6[15]);
assign Ro88v6 = (F0eiw6 ? Icn7z6[16] : Hjn7z6[16]);
assign Ko88v6 = (F0eiw6 ? Icn7z6[17] : Hjn7z6[17]);
assign Do88v6 = (F0eiw6 ? Icn7z6[18] : Hjn7z6[18]);
assign Wn88v6 = (F0eiw6 ? Icn7z6[19] : Hjn7z6[19]);
assign Pn88v6 = (F0eiw6 ? Icn7z6[20] : Hjn7z6[20]);
assign In88v6 = (F0eiw6 ? Icn7z6[21] : Hjn7z6[21]);
assign Bn88v6 = (F0eiw6 ? Icn7z6[22] : Hjn7z6[22]);
assign Um88v6 = (F0eiw6 ? Icn7z6[23] : Hjn7z6[23]);
assign Nm88v6 = (F0eiw6 ? Icn7z6[24] : Hjn7z6[24]);
assign F0eiw6 = (!M0eiw6);
assign Gm88v6 = (M0eiw6 ? Hjn7z6[25] : Icn7z6[25]);
assign Zl88v6 = (M0eiw6 ? Hjn7z6[26] : Icn7z6[26]);
assign Sl88v6 = (M0eiw6 ? Hjn7z6[27] : Icn7z6[27]);
assign Ll88v6 = (M0eiw6 ? Hjn7z6[28] : Icn7z6[28]);
assign El88v6 = (M0eiw6 ? Hjn7z6[29] : Icn7z6[29]);
assign Xk88v6 = (M0eiw6 ? Hjn7z6[30] : Icn7z6[30]);
assign Qk88v6 = (M0eiw6 ? Hjn7z6[31] : Icn7z6[31]);
assign M0eiw6 = (T0eiw6 & N0qhw6);
assign T0eiw6 = (~(A1eiw6 & H1eiw6));
assign H1eiw6 = (X02iw6 & O1eiw6);
assign A1eiw6 = (V1eiw6 & C2eiw6);
assign C2eiw6 = (~(J2eiw6 & Q2eiw6));
assign Q2eiw6 = (~(N22iw6 & Kjonv6));
assign Jk88v6 = (~(X2eiw6 & E3eiw6));
assign E3eiw6 = (~(Hl9ov6 & L3eiw6));
assign Hl9ov6 = (~(U22iw6 | Dq9ov6));
assign X2eiw6 = (~(Dq9ov6 & Qln7z6[0]));
assign Dq9ov6 = (~(U22iw6 | S3eiw6));
assign U22iw6 = (!Jalov6);
assign Ck88v6 = (~(Z3eiw6 & G4eiw6));
assign G4eiw6 = (~(Teyet6 & N4eiw6));
assign Z3eiw6 = (U4eiw6 | N4eiw6);
assign N4eiw6 = (~(O1eiw6 & B5eiw6));
assign B5eiw6 = (~(I5eiw6 & P5eiw6));
assign P5eiw6 = (~(S12iw6 | A4qhw6));
assign I5eiw6 = (~(X02iw6 | N22iw6));
assign U4eiw6 = (W5eiw6 | D6eiw6);
assign Vj88v6 = (Uimov6 ? X7pet6 : Yhqnv6);
assign Oj88v6 = (Uimov6 ? W5pet6 : Pgqnv6);
assign Hj88v6 = (Uimov6 ? V3pet6 : Gfqnv6);
assign Uimov6 = (!Sblov6);
assign Aj88v6 = (Sblov6 ? Qdqnv6 : U1pet6);
assign Ti88v6 = (~(K6eiw6 & R6eiw6));
assign R6eiw6 = (~(P39iw6 & Ebdiw6));
assign K6eiw6 = (~(J09iw6 & Hyj7z6[3]));
assign Mi88v6 = (~(Y6eiw6 & F7eiw6));
assign F7eiw6 = (~(H9diw6 & P39iw6));
assign P39iw6 = (~(I52nv6 | J09iw6));
assign H9diw6 = (L19iw6 & U42nv6);
assign Y6eiw6 = (~(J09iw6 & Hyj7z6[1]));
assign J09iw6 = (!N29iw6);
assign Fi88v6 = (N29iw6 ? Ucdiw6 : Hyj7z6[5]);
assign N29iw6 = (~(M7eiw6 & F8diw6));
assign F8diw6 = (~(T7eiw6 & A8eiw6));
assign A8eiw6 = (Ptbiw6 & W52nv6);
assign T7eiw6 = (H8eiw6 & Pohov6);
assign M7eiw6 = (~(O8eiw6 & V8eiw6));
assign V8eiw6 = (C9eiw6 & J9eiw6);
assign J9eiw6 = (~(Dtj7z6[2] | Dtj7z6[5]));
assign C9eiw6 = (Hc3iw6 & Q9eiw6);
assign Hc3iw6 = (Pvj7z6[0] & Cd3iw6);
assign Cd3iw6 = (Rediw6 | H8eiw6);
assign H8eiw6 = (X9eiw6 & Eaeiw6);
assign Eaeiw6 = (Laeiw6 & Pvj7z6[1]);
assign Laeiw6 = (Pvj7z6[0] & Hkget6);
assign X9eiw6 = (Pvj7z6[3] & Pvj7z6[2]);
assign O8eiw6 = (Saeiw6 & Zaeiw6);
assign Saeiw6 = (Gbeiw6 & Nbeiw6);
assign Yh88v6 = (~(Ubeiw6 & Bceiw6));
assign Bceiw6 = (~(Ohj7z6[0] & Iceiw6));
assign Iceiw6 = (~(Qn7iw6 & U42nv6));
assign Qn7iw6 = (~(Mh4iw6 | Twaiw6));
assign Mh4iw6 = (~(Pceiw6 & Wceiw6));
assign Ubeiw6 = (~(Ip8iw6 & U42nv6));
assign Ip8iw6 = (Jz2iw6 & Bqi7z6[0]);
assign Jz2iw6 = (Ddeiw6 & Wceiw6);
assign Rh88v6 = (~(Kdeiw6 & Rdeiw6));
assign Rdeiw6 = (~(Ohj7z6[32] & Ydeiw6));
assign Ydeiw6 = (~(So7iw6 & U42nv6));
assign So7iw6 = (~(Oi4iw6 | Twaiw6));
assign Oi4iw6 = (~(Feeiw6 & Wceiw6));
assign Kdeiw6 = (~(Kq8iw6 & U42nv6));
assign Kq8iw6 = (Ay2iw6 & Bqi7z6[0]);
assign Ay2iw6 = (Meeiw6 & Wceiw6);
assign Wceiw6 = (Teeiw6 & Afeiw6);
assign Afeiw6 = (~(Hfeiw6 | Toi7z6[9]));
assign Kh88v6 = (Vfeiw6 ? Ofeiw6 : Klo7z6[0]);
assign Dh88v6 = (~(Cgeiw6 & Jgeiw6));
assign Jgeiw6 = (~(Qgeiw6 & Xgeiw6));
assign Cgeiw6 = (~(Klo7z6[6] & Eheiw6));
assign Wg88v6 = (~(Lheiw6 & Sheiw6));
assign Sheiw6 = (~(Xgeiw6 & N13iw6));
assign Lheiw6 = (~(Eheiw6 & Klo7z6[5]));
assign Pg88v6 = (~(Zheiw6 & Gieiw6));
assign Gieiw6 = (~(Nieiw6 & Xgeiw6));
assign Xgeiw6 = (G13iw6 & Vfeiw6);
assign G13iw6 = (Uieiw6 & Bjeiw6);
assign Bjeiw6 = (Ijeiw6 & Pjeiw6);
assign Ijeiw6 = (Wjeiw6 & Dkeiw6);
assign Uieiw6 = (Kkeiw6 & Rkeiw6);
assign Nieiw6 = (~(N13iw6 | Qgeiw6));
assign Qgeiw6 = (Ykeiw6 & Fleiw6);
assign Fleiw6 = (X72iw6 & E82iw6);
assign Ykeiw6 = (~(Mleiw6 | V62iw6));
assign N13iw6 = (Tleiw6 & Ameiw6);
assign Ameiw6 = (~(Hmeiw6 | Omeiw6));
assign Omeiw6 = (!J72iw6);
assign Tleiw6 = (Vmeiw6 & Cneiw6);
assign Zheiw6 = (~(Klo7z6[4] & Eheiw6));
assign Ig88v6 = (Vfeiw6 ? Jneiw6 : Klo7z6[3]);
assign Vfeiw6 = (!Eheiw6);
assign Bg88v6 = (Eheiw6 ? Klo7z6[2] : Yelov6);
assign Uf88v6 = (Eheiw6 ? Klo7z6[1] : Fflov6);
assign Eheiw6 = (C63iw6 & Qneiw6);
assign Qneiw6 = (~(Xneiw6 & Vd2iw6));
assign Nf88v6 = (~(Eoeiw6 & Loeiw6));
assign Loeiw6 = (~(Soeiw6 & D42iw6));
assign Eoeiw6 = (~(D02ft6 & Pdlov6));
assign Gf88v6 = (Zoeiw6 ? Z4p7z6[1] : L82iw6);
assign Ze88v6 = (Zoeiw6 ? Z4p7z6[2] : E82iw6);
assign Se88v6 = (Zoeiw6 ? Z4p7z6[3] : X72iw6);
assign Le88v6 = (!Gpeiw6);
assign Gpeiw6 = (Zoeiw6 ? Upeiw6 : Npeiw6);
assign Zoeiw6 = (!Soeiw6);
assign Npeiw6 = (~(Bqeiw6 & Iqeiw6));
assign Bqeiw6 = (Cneiw6 & Pqeiw6);
assign Pqeiw6 = (~(X72iw6 & Wqeiw6));
assign Wqeiw6 = (L82iw6 | E82iw6);
assign Ee88v6 = (Soeiw6 ? Dreiw6 : Z4p7z6[5]);
assign Dreiw6 = (Kreiw6 & Rreiw6);
assign Rreiw6 = (J72iw6 & V62iw6);
assign Kreiw6 = (~(Hmeiw6 | Cneiw6));
assign Cneiw6 = (!Q72iw6);
assign Hmeiw6 = (~(Yreiw6 & Fseiw6));
assign Fseiw6 = (A62iw6 & O62iw6);
assign Yreiw6 = (T43iw6 & C72iw6);
assign T43iw6 = (~(Mseiw6 & Tseiw6));
assign Tseiw6 = (!X72iw6);
assign Mseiw6 = (!E82iw6);
assign Xd88v6 = (Soeiw6 ? S82iw6 : Z4p7z6[0]);
assign Soeiw6 = (~(Ateiw6 | Da3iw6));
assign Ateiw6 = (!Yelov6);
assign Yelov6 = (Hteiw6 & Rkeiw6);
assign Hteiw6 = (Oteiw6 & Dkeiw6);
assign Qd88v6 = (Vteiw6 ? Nmq7z6[3] : L82iw6);
assign Jd88v6 = (Vteiw6 ? Nmq7z6[4] : E82iw6);
assign Cd88v6 = (Vteiw6 ? Nmq7z6[5] : X72iw6);
assign Vc88v6 = (Vteiw6 ? Nmq7z6[6] : Q72iw6);
assign Oc88v6 = (Vteiw6 ? Cueiw6 : D42iw6);
assign Hc88v6 = (!Jueiw6);
assign Jueiw6 = (Vteiw6 ? Xueiw6 : Queiw6);
assign Queiw6 = (Iqeiw6 & Eveiw6);
assign Eveiw6 = (~(Q72iw6 & X72iw6));
assign Ac88v6 = (!Lveiw6);
assign Lveiw6 = (Vteiw6 ? Zveiw6 : Sveiw6);
assign Vteiw6 = (!Zdo7v6);
assign Sveiw6 = (Mleiw6 | Vmeiw6);
assign Vmeiw6 = (!V62iw6);
assign Mleiw6 = (~(Gweiw6 & Nweiw6));
assign Nweiw6 = (Uweiw6 & O62iw6);
assign Uweiw6 = (Q72iw6 & J72iw6);
assign Gweiw6 = (C72iw6 & A62iw6);
assign Tb88v6 = (Zdo7v6 ? S82iw6 : Bxeiw6);
assign Mb88v6 = (Ixeiw6 & Pxeiw6);
assign Pxeiw6 = (~(Wxeiw6 | Sgp7z6[2]));
assign Ixeiw6 = (Sgp7z6[3] & HTMDHBURST[0]);
assign Fb88v6 = (Ypinv6 ? Kg5ft6 : Dyeiw6);
assign Dyeiw6 = (Kyeiw6 & Ryeiw6);
assign Kyeiw6 = (~(Yyeiw6 & Fzeiw6));
assign Fzeiw6 = (~(Sgp7z6[1] & Mzeiw6));
assign Yyeiw6 = (~(Tzeiw6 & A0fiw6));
assign Ya88v6 = (Ypinv6 ? Dw4ft6 : H0fiw6);
assign H0fiw6 = (O0fiw6 & V0fiw6);
assign O0fiw6 = (~(C1fiw6 & J1fiw6));
assign J1fiw6 = (Q1fiw6 | X1fiw6);
assign C1fiw6 = (~(E2fiw6 & L2fiw6));
assign Ra88v6 = (K94iw6 ? Fy4ft6 : S2fiw6);
assign Ka88v6 = (Z2fiw6 ? Zdp7z6[1] : Gpgnv6);
assign Z2fiw6 = (Kygnv6 & B1rnv6);
assign Da88v6 = (~(G3fiw6 & N3fiw6));
assign N3fiw6 = (~(U3fiw6 & Zidiw6));
assign U3fiw6 = (Jx5ov6 & Zc5ft6);
assign Jx5ov6 = (!B4fiw6);
assign G3fiw6 = (~(B82ft6 & K94iw6));
assign W988v6 = (~(I4fiw6 & P4fiw6));
assign P4fiw6 = (~(W4fiw6 & Zidiw6));
assign W4fiw6 = (Hw5ov6 & Xn5ft6);
assign Hw5ov6 = (!D5fiw6);
assign I4fiw6 = (~(Y52ft6 & K94iw6));
assign P988v6 = (K5fiw6 ? Zdp7z6[3] : V1gnv6);
assign K5fiw6 = (Kygnv6 & U0rnv6);
assign V1gnv6 = (R5fiw6 & Y5fiw6);
assign Y5fiw6 = (F6fiw6 & D5fiw6);
assign R5fiw6 = (M6fiw6 & T6fiw6);
assign I988v6 = (~(A7fiw6 & H7fiw6));
assign H7fiw6 = (~(O7fiw6 & U9p7z6[0]));
assign A7fiw6 = (V7fiw6 & C8fiw6);
assign C8fiw6 = (~(L84ft6 & J8fiw6));
assign V7fiw6 = (Q8fiw6 | Orhov6);
assign B988v6 = (~(X8fiw6 & E9fiw6));
assign E9fiw6 = (~(O7fiw6 & U9p7z6[1]));
assign X8fiw6 = (L9fiw6 & S9fiw6);
assign S9fiw6 = (~(A74ft6 & J8fiw6));
assign L9fiw6 = (Q8fiw6 | L19iw6);
assign U888v6 = (~(Z9fiw6 & Gafiw6));
assign Gafiw6 = (~(O7fiw6 & U9p7z6[2]));
assign Z9fiw6 = (Nafiw6 & Uafiw6);
assign Uafiw6 = (~(P54ft6 & J8fiw6));
assign Nafiw6 = (Q8fiw6 | Fhrnv6);
assign N888v6 = (~(Bbfiw6 & Ibfiw6));
assign Ibfiw6 = (Q8fiw6 | Pohov6);
assign Bbfiw6 = (Pbfiw6 & Wbfiw6);
assign Wbfiw6 = (~(E44ft6 & J8fiw6));
assign Pbfiw6 = (~(O7fiw6 & U9p7z6[3]));
assign G888v6 = (~(Dcfiw6 & Kcfiw6));
assign Kcfiw6 = (Q8fiw6 | Zaeiw6);
assign Dcfiw6 = (Rcfiw6 & Ycfiw6);
assign Ycfiw6 = (~(T24ft6 & J8fiw6));
assign Rcfiw6 = (~(O7fiw6 & U9p7z6[4]));
assign Z788v6 = (~(Fdfiw6 & Mdfiw6));
assign Mdfiw6 = (Q8fiw6 | Tdfiw6);
assign Fdfiw6 = (Aefiw6 & Hefiw6);
assign Hefiw6 = (~(I14ft6 & J8fiw6));
assign Aefiw6 = (~(O7fiw6 & U9p7z6[5]));
assign S788v6 = (~(Oefiw6 & Vefiw6));
assign Vefiw6 = (Q8fiw6 | Gbeiw6);
assign Oefiw6 = (Cffiw6 & Jffiw6);
assign Jffiw6 = (~(Xz3ft6 & J8fiw6));
assign Cffiw6 = (~(O7fiw6 & U9p7z6[6]));
assign L788v6 = (~(Qffiw6 & Xffiw6));
assign Xffiw6 = (Q8fiw6 | Egfiw6);
assign Qffiw6 = (Lgfiw6 & Sgfiw6);
assign Sgfiw6 = (~(My3ft6 & J8fiw6));
assign Lgfiw6 = (~(O7fiw6 & U9p7z6[7]));
assign E788v6 = (~(Zgfiw6 & Ghfiw6));
assign Ghfiw6 = (Q8fiw6 | Nhfiw6);
assign Zgfiw6 = (Uhfiw6 & Bifiw6);
assign Bifiw6 = (~(Bx3ft6 & J8fiw6));
assign Uhfiw6 = (~(O7fiw6 & U9p7z6[8]));
assign X688v6 = (~(Iifiw6 & Pifiw6));
assign Pifiw6 = (Q8fiw6 | Wifiw6);
assign Iifiw6 = (Djfiw6 & Kjfiw6);
assign Kjfiw6 = (~(Qv3ft6 & J8fiw6));
assign Djfiw6 = (~(O7fiw6 & U9p7z6[9]));
assign Q688v6 = (~(Rjfiw6 & Yjfiw6));
assign Yjfiw6 = (Q8fiw6 | Fkfiw6);
assign Rjfiw6 = (Mkfiw6 & Tkfiw6);
assign Tkfiw6 = (~(Fu3ft6 & J8fiw6));
assign Mkfiw6 = (~(O7fiw6 & U9p7z6[10]));
assign J688v6 = (~(Alfiw6 & Hlfiw6));
assign Hlfiw6 = (Q8fiw6 | Olfiw6);
assign Alfiw6 = (Vlfiw6 & Cmfiw6);
assign Cmfiw6 = (~(Us3ft6 & J8fiw6));
assign Vlfiw6 = (~(O7fiw6 & U9p7z6[11]));
assign C688v6 = (~(Jmfiw6 & Qmfiw6));
assign Qmfiw6 = (Q8fiw6 | Xmfiw6);
assign Jmfiw6 = (Enfiw6 & Lnfiw6);
assign Lnfiw6 = (~(Jr3ft6 & J8fiw6));
assign Enfiw6 = (~(O7fiw6 & U9p7z6[12]));
assign V588v6 = (~(Snfiw6 & Znfiw6));
assign Znfiw6 = (Q8fiw6 | Gofiw6);
assign Snfiw6 = (Nofiw6 & Uofiw6);
assign Uofiw6 = (~(Yp3ft6 & J8fiw6));
assign Nofiw6 = (~(O7fiw6 & U9p7z6[13]));
assign O588v6 = (~(Bpfiw6 & Ipfiw6));
assign Ipfiw6 = (Q8fiw6 | Ppfiw6);
assign Bpfiw6 = (Wpfiw6 & Dqfiw6);
assign Dqfiw6 = (~(No3ft6 & J8fiw6));
assign Wpfiw6 = (~(O7fiw6 & U9p7z6[14]));
assign H588v6 = (~(Kqfiw6 & Rqfiw6));
assign Rqfiw6 = (Q8fiw6 | Yqfiw6);
assign Kqfiw6 = (Frfiw6 & Mrfiw6);
assign Mrfiw6 = (~(Cn3ft6 & J8fiw6));
assign Frfiw6 = (~(O7fiw6 & U9p7z6[15]));
assign A588v6 = (~(Trfiw6 & Asfiw6));
assign Asfiw6 = (Q8fiw6 | Hsfiw6);
assign Trfiw6 = (Osfiw6 & Vsfiw6);
assign Vsfiw6 = (~(Rl3ft6 & J8fiw6));
assign Osfiw6 = (~(O7fiw6 & U9p7z6[16]));
assign T488v6 = (~(Ctfiw6 & Jtfiw6));
assign Jtfiw6 = (Q8fiw6 | Oyhov6);
assign Ctfiw6 = (Qtfiw6 & Xtfiw6);
assign Xtfiw6 = (~(Gk3ft6 & J8fiw6));
assign Qtfiw6 = (~(O7fiw6 & U9p7z6[17]));
assign M488v6 = (~(Eufiw6 & Lufiw6));
assign Lufiw6 = (Q8fiw6 | Sufiw6);
assign Eufiw6 = (Zufiw6 & Gvfiw6);
assign Gvfiw6 = (~(Vi3ft6 & J8fiw6));
assign Zufiw6 = (~(O7fiw6 & U9p7z6[18]));
assign F488v6 = (~(Nvfiw6 & Uvfiw6));
assign Uvfiw6 = (Q8fiw6 | Bwfiw6);
assign Nvfiw6 = (Iwfiw6 & Pwfiw6);
assign Pwfiw6 = (~(Kh3ft6 & J8fiw6));
assign Iwfiw6 = (~(O7fiw6 & U9p7z6[19]));
assign Y388v6 = (~(Wwfiw6 & Dxfiw6));
assign Dxfiw6 = (Q8fiw6 | Kxfiw6);
assign Wwfiw6 = (Rxfiw6 & Yxfiw6);
assign Yxfiw6 = (~(Zf3ft6 & J8fiw6));
assign Rxfiw6 = (~(O7fiw6 & U9p7z6[20]));
assign R388v6 = (~(Fyfiw6 & Myfiw6));
assign Myfiw6 = (Q8fiw6 | Tyfiw6);
assign Fyfiw6 = (Azfiw6 & Hzfiw6);
assign Hzfiw6 = (~(Oe3ft6 & J8fiw6));
assign Azfiw6 = (~(O7fiw6 & U9p7z6[21]));
assign K388v6 = (~(Ozfiw6 & Vzfiw6));
assign Vzfiw6 = (Q8fiw6 | C0giw6);
assign Ozfiw6 = (J0giw6 & Q0giw6);
assign Q0giw6 = (~(Dd3ft6 & J8fiw6));
assign J0giw6 = (~(O7fiw6 & U9p7z6[22]));
assign D388v6 = (~(X0giw6 & E1giw6));
assign E1giw6 = (Q8fiw6 | L1giw6);
assign X0giw6 = (S1giw6 & Z1giw6);
assign Z1giw6 = (~(Sb3ft6 & J8fiw6));
assign S1giw6 = (~(O7fiw6 & U9p7z6[23]));
assign W288v6 = (~(G2giw6 & N2giw6));
assign N2giw6 = (Q8fiw6 | U2giw6);
assign G2giw6 = (B3giw6 & I3giw6);
assign I3giw6 = (~(Ha3ft6 & J8fiw6));
assign B3giw6 = (~(O7fiw6 & U9p7z6[24]));
assign P288v6 = (~(P3giw6 & W3giw6));
assign W3giw6 = (Q8fiw6 | D4giw6);
assign P3giw6 = (K4giw6 & R4giw6);
assign R4giw6 = (~(W83ft6 & J8fiw6));
assign K4giw6 = (~(O7fiw6 & U9p7z6[25]));
assign I288v6 = (~(Y4giw6 & F5giw6));
assign F5giw6 = (Q8fiw6 | M5giw6);
assign Y4giw6 = (T5giw6 & A6giw6);
assign A6giw6 = (~(L73ft6 & J8fiw6));
assign T5giw6 = (~(O7fiw6 & U9p7z6[26]));
assign B288v6 = (~(H6giw6 & O6giw6));
assign O6giw6 = (Q8fiw6 | V6giw6);
assign H6giw6 = (C7giw6 & J7giw6);
assign J7giw6 = (~(A63ft6 & J8fiw6));
assign C7giw6 = (~(O7fiw6 & U9p7z6[27]));
assign U188v6 = (~(Q7giw6 & X7giw6));
assign X7giw6 = (Q8fiw6 | E8giw6);
assign Q7giw6 = (L8giw6 & S8giw6);
assign S8giw6 = (~(P43ft6 & J8fiw6));
assign L8giw6 = (~(O7fiw6 & U9p7z6[28]));
assign N188v6 = (~(Z8giw6 & G9giw6));
assign G9giw6 = (Q8fiw6 | N9giw6);
assign Z8giw6 = (U9giw6 & Bagiw6);
assign Bagiw6 = (~(E33ft6 & J8fiw6));
assign U9giw6 = (~(O7fiw6 & U9p7z6[29]));
assign G188v6 = (~(Iagiw6 & Pagiw6));
assign Pagiw6 = (Q8fiw6 | Wagiw6);
assign Iagiw6 = (Dbgiw6 & Kbgiw6);
assign Kbgiw6 = (~(T13ft6 & J8fiw6));
assign Dbgiw6 = (~(O7fiw6 & U9p7z6[30]));
assign Z088v6 = (~(Rbgiw6 & Ybgiw6));
assign Ybgiw6 = (Q8fiw6 | Fcgiw6);
assign Rbgiw6 = (Mcgiw6 & Tcgiw6);
assign Tcgiw6 = (~(I03ft6 & J8fiw6));
assign J8fiw6 = (Adgiw6 & Q8fiw6);
assign Adgiw6 = (!O7fiw6);
assign Mcgiw6 = (~(O7fiw6 & U9p7z6[31]));
assign S088v6 = (~(Hdgiw6 & Odgiw6));
assign Odgiw6 = (~(Vdgiw6 & Zidiw6));
assign Zidiw6 = (~(Cegiw6 | Kygnv6));
assign Vdgiw6 = (Cx5ov6 & Fs4ft6);
assign Hdgiw6 = (~(Hc2ft6 & K94iw6));
assign L088v6 = (~(Jegiw6 & Qegiw6));
assign Qegiw6 = (~(Xegiw6 & U42nv6));
assign Jegiw6 = (Tbq7z6[0] ? Lfgiw6 : Efgiw6);
assign E088v6 = (~(Sfgiw6 & Zfgiw6));
assign Zfgiw6 = (~(Xegiw6 & B52nv6));
assign Sfgiw6 = (Tbq7z6[1] ? Nggiw6 : Gggiw6);
assign Gggiw6 = (~(Uggiw6 & Tbq7z6[0]));
assign Xz78v6 = (~(Bhgiw6 & Ihgiw6));
assign Ihgiw6 = (Phgiw6 | Fhrnv6);
assign Bhgiw6 = (Tbq7z6[2] ? Digiw6 : Whgiw6);
assign Digiw6 = (Nggiw6 & Kigiw6);
assign Kigiw6 = (Efgiw6 | Tbq7z6[1]);
assign Nggiw6 = (Lfgiw6 & Rigiw6);
assign Rigiw6 = (Efgiw6 | Tbq7z6[0]);
assign Whgiw6 = (~(Yigiw6 & Uggiw6));
assign Qz78v6 = (~(Fjgiw6 & Mjgiw6));
assign Mjgiw6 = (~(Xegiw6 & P52nv6));
assign Fjgiw6 = (Tbq7z6[3] ? Akgiw6 : Tjgiw6);
assign Tjgiw6 = (~(Hkgiw6 & Uggiw6));
assign Jz78v6 = (~(Okgiw6 & Vkgiw6));
assign Vkgiw6 = (Phgiw6 | Zaeiw6);
assign Okgiw6 = (Tbq7z6[4] ? Jlgiw6 : Clgiw6);
assign Jlgiw6 = (Akgiw6 & Qlgiw6);
assign Qlgiw6 = (Efgiw6 | Tbq7z6[3]);
assign Akgiw6 = (Lfgiw6 & Xlgiw6);
assign Xlgiw6 = (Efgiw6 | Hkgiw6);
assign Clgiw6 = (~(Emgiw6 & Hkgiw6));
assign Emgiw6 = (Uggiw6 & Tbq7z6[3]);
assign Cz78v6 = (~(Lmgiw6 & Smgiw6));
assign Smgiw6 = (~(Xegiw6 & D62nv6));
assign Lmgiw6 = (Tbq7z6[5] ? Gngiw6 : Zmgiw6);
assign Zmgiw6 = (~(Nngiw6 & Uggiw6));
assign Vy78v6 = (~(Ungiw6 & Bogiw6));
assign Bogiw6 = (~(Xegiw6 & K62nv6));
assign Xegiw6 = (!Phgiw6);
assign Ungiw6 = (Tbq7z6[6] ? Pogiw6 : Iogiw6);
assign Oy78v6 = (~(Wogiw6 & Dpgiw6));
assign Dpgiw6 = (Phgiw6 | Egfiw6);
assign Wogiw6 = (Tbq7z6[7] ? Rpgiw6 : Kpgiw6);
assign Rpgiw6 = (Pogiw6 & Ypgiw6);
assign Ypgiw6 = (~(Uggiw6 & Fqgiw6));
assign Pogiw6 = (Gngiw6 & Mqgiw6);
assign Mqgiw6 = (Efgiw6 | Tbq7z6[5]);
assign Gngiw6 = (Lfgiw6 & Tqgiw6);
assign Tqgiw6 = (Efgiw6 | Nngiw6);
assign Kpgiw6 = (Iogiw6 | Fqgiw6);
assign Fqgiw6 = (!Tbq7z6[6]);
assign Iogiw6 = (~(Argiw6 & Nngiw6));
assign Argiw6 = (Uggiw6 & Tbq7z6[5]);
assign Uggiw6 = (!Efgiw6);
assign Efgiw6 = (~(Hrgiw6 & Orgiw6));
assign Hrgiw6 = (Lfgiw6 & Phgiw6);
assign Lfgiw6 = (Vrgiw6 | Csgiw6);
assign Vrgiw6 = (~(Orgiw6 & Phgiw6));
assign Phgiw6 = (~(Jsgiw6 & Qsgiw6));
assign Orgiw6 = (~(Xsgiw6 & Etgiw6));
assign Xsgiw6 = (Ltgiw6 & Ej5iw6);
assign Ltgiw6 = (~(Xkq7z6[21] & HTMDHBURST[0]));
assign Hy78v6 = (~(Stgiw6 & Ztgiw6));
assign Ztgiw6 = (~(Gugiw6 & U42nv6));
assign Stgiw6 = (Kfq7z6[0] ? Uugiw6 : Nugiw6);
assign Ay78v6 = (~(Bvgiw6 & Ivgiw6));
assign Ivgiw6 = (~(Gugiw6 & B52nv6));
assign Bvgiw6 = (Kfq7z6[1] ? Wvgiw6 : Pvgiw6);
assign Pvgiw6 = (~(Dwgiw6 & Kfq7z6[0]));
assign Tx78v6 = (~(Kwgiw6 & Rwgiw6));
assign Rwgiw6 = (Ywgiw6 | Fhrnv6);
assign Kwgiw6 = (Kfq7z6[2] ? Mxgiw6 : Fxgiw6);
assign Mxgiw6 = (Wvgiw6 & Txgiw6);
assign Txgiw6 = (Nugiw6 | Kfq7z6[1]);
assign Wvgiw6 = (Uugiw6 & Aygiw6);
assign Aygiw6 = (Nugiw6 | Kfq7z6[0]);
assign Fxgiw6 = (~(Hygiw6 & Dwgiw6));
assign Mx78v6 = (~(Oygiw6 & Vygiw6));
assign Vygiw6 = (~(Gugiw6 & P52nv6));
assign Oygiw6 = (Kfq7z6[3] ? Jzgiw6 : Czgiw6);
assign Czgiw6 = (~(Qzgiw6 & Dwgiw6));
assign Fx78v6 = (~(Xzgiw6 & E0hiw6));
assign E0hiw6 = (Ywgiw6 | Zaeiw6);
assign Xzgiw6 = (Kfq7z6[4] ? S0hiw6 : L0hiw6);
assign S0hiw6 = (Jzgiw6 & Z0hiw6);
assign Z0hiw6 = (Nugiw6 | Kfq7z6[3]);
assign Jzgiw6 = (Uugiw6 & G1hiw6);
assign G1hiw6 = (Nugiw6 | Qzgiw6);
assign L0hiw6 = (~(N1hiw6 & Qzgiw6));
assign N1hiw6 = (Dwgiw6 & Kfq7z6[3]);
assign Yw78v6 = (~(U1hiw6 & B2hiw6));
assign B2hiw6 = (~(Gugiw6 & D62nv6));
assign U1hiw6 = (Kfq7z6[5] ? P2hiw6 : I2hiw6);
assign I2hiw6 = (~(W2hiw6 & Dwgiw6));
assign Rw78v6 = (~(D3hiw6 & K3hiw6));
assign K3hiw6 = (~(Gugiw6 & K62nv6));
assign Gugiw6 = (!Ywgiw6);
assign D3hiw6 = (Kfq7z6[6] ? Y3hiw6 : R3hiw6);
assign Kw78v6 = (~(F4hiw6 & M4hiw6));
assign M4hiw6 = (Ywgiw6 | Egfiw6);
assign F4hiw6 = (Kfq7z6[7] ? A5hiw6 : T4hiw6);
assign A5hiw6 = (Y3hiw6 & H5hiw6);
assign H5hiw6 = (~(Dwgiw6 & O5hiw6));
assign Y3hiw6 = (P2hiw6 & V5hiw6);
assign V5hiw6 = (Nugiw6 | Kfq7z6[5]);
assign P2hiw6 = (Uugiw6 & C6hiw6);
assign C6hiw6 = (Nugiw6 | W2hiw6);
assign T4hiw6 = (R3hiw6 | O5hiw6);
assign O5hiw6 = (!Kfq7z6[6]);
assign R3hiw6 = (~(J6hiw6 & W2hiw6));
assign J6hiw6 = (Dwgiw6 & Kfq7z6[5]);
assign Dwgiw6 = (!Nugiw6);
assign Nugiw6 = (~(Q6hiw6 & X6hiw6));
assign Q6hiw6 = (Uugiw6 & Ywgiw6);
assign Uugiw6 = (E7hiw6 | L7hiw6);
assign E7hiw6 = (~(X6hiw6 & Ywgiw6));
assign Ywgiw6 = (~(Jsgiw6 & S7hiw6));
assign X6hiw6 = (~(Z7hiw6 & Etgiw6));
assign Z7hiw6 = (G8hiw6 & Mn5iw6);
assign G8hiw6 = (~(Xkq7z6[19] & HTMDHBURST[0]));
assign Dw78v6 = (~(N8hiw6 & U8hiw6));
assign U8hiw6 = (~(B9hiw6 & I9hiw6));
assign I9hiw6 = (P9hiw6 & W9hiw6);
assign W9hiw6 = (W5q7z6[1] | W5q7z6[0]);
assign P9hiw6 = (~(Txadt6 | Gw2ft6));
assign B9hiw6 = (Dahiw6 & Qb4ft6);
assign Dahiw6 = (A9i8v6 & HTMDHBURST[0]);
assign N8hiw6 = (~(Kahiw6 & Rahiw6));
assign Rahiw6 = (Yahiw6 & Fbhiw6);
assign Fbhiw6 = (Hu2ft6 ^ Mbhiw6);
assign Yahiw6 = (Tbhiw6 & Zb1nv6);
assign Tbhiw6 = (~(Gw2ft6 & O7fiw6));
assign Kahiw6 = (Qb4ft6 & HTMDHBURST[0]);
assign Wv78v6 = (~(Achiw6 & Hchiw6));
assign Hchiw6 = (Ochiw6 & Vchiw6);
assign Ochiw6 = (~(Cdhiw6 & Y7q7z6[0]));
assign Achiw6 = (Jdhiw6 & Qdhiw6);
assign Qdhiw6 = (~(W3q7z6[0] & Xdhiw6));
assign Jdhiw6 = (~(Eehiw6 & X9q7z6[0]));
assign Pv78v6 = (~(Lehiw6 & Sehiw6));
assign Sehiw6 = (W3q7z6[1] ? Zehiw6 : Vchiw6);
assign Lehiw6 = (Gfhiw6 & Nfhiw6);
assign Nfhiw6 = (~(Cdhiw6 & Y7q7z6[1]));
assign Gfhiw6 = (~(Eehiw6 & X9q7z6[1]));
assign Iv78v6 = (~(Ufhiw6 & Bghiw6));
assign Bghiw6 = (W3q7z6[2] ? Pghiw6 : Ighiw6);
assign Ighiw6 = (Vchiw6 | W3q7z6[1]);
assign Vchiw6 = (~(Wghiw6 & Dhhiw6));
assign Dhhiw6 = (~(Khhiw6 | W3q7z6[0]));
assign Ufhiw6 = (Rhhiw6 & Yhhiw6);
assign Yhhiw6 = (~(Cdhiw6 & Y7q7z6[2]));
assign Rhhiw6 = (~(Eehiw6 & X9q7z6[2]));
assign Bv78v6 = (~(Fihiw6 & Mihiw6));
assign Mihiw6 = (~(Eehiw6 & X9q7z6[3]));
assign Fihiw6 = (Tihiw6 & Ajhiw6);
assign Ajhiw6 = (~(W3q7z6[3] & Hjhiw6));
assign Hjhiw6 = (~(Pghiw6 & Ojhiw6));
assign Ojhiw6 = (~(W3q7z6[2] & Vjhiw6));
assign Pghiw6 = (Zehiw6 & Ckhiw6);
assign Ckhiw6 = (~(W3q7z6[1] & Vjhiw6));
assign Zehiw6 = (Jkhiw6 & Qkhiw6);
assign Qkhiw6 = (~(W3q7z6[0] & Vjhiw6));
assign Tihiw6 = (~(Cdhiw6 & Y7q7z6[3]));
assign Cdhiw6 = (Wghiw6 & Khhiw6);
assign Wghiw6 = (Jkhiw6 & Vjhiw6);
assign Jkhiw6 = (!Xdhiw6);
assign Xdhiw6 = (~(Eehiw6 | Xkhiw6));
assign Eehiw6 = (!Vjhiw6);
assign Vjhiw6 = (~(Etgiw6 & Elhiw6));
assign Elhiw6 = (~(Llhiw6 & Slhiw6));
assign Slhiw6 = (~(Zlhiw6 & Gmhiw6));
assign Zlhiw6 = (~(Xmfiw6 & Nmhiw6));
assign Nmhiw6 = (C0giw6 | Xkq7z6[22]);
assign Llhiw6 = (Umhiw6 | HTMDHBURST[0]);
assign Uu78v6 = (Inhiw6 ? Cu5ft6 : Bnhiw6);
assign Nu78v6 = (~(Pnhiw6 & Wnhiw6));
assign Wnhiw6 = (~(W2adt6 & Dohiw6));
assign Dohiw6 = (D16ft6 | Kohiw6);
assign Kohiw6 = (~(Sdo7v6 | K2adt6));
assign Pnhiw6 = (~(Sdo7v6 & D42iw6));
assign Gu78v6 = (!Rohiw6);
assign Rohiw6 = (Mphiw6 ? Fphiw6 : Yohiw6);
assign Fphiw6 = (~(W2adt6 & Tphiw6));
assign Tphiw6 = (!K2adt6);
assign Zt78v6 = (W5fov6 ? Pjb7z6[2] : S82iw6);
assign St78v6 = (W5fov6 ? Pjb7z6[18] : Aqhiw6);
assign Lt78v6 = (W5fov6 ? Pjb7z6[17] : Hqhiw6);
assign Et78v6 = (!Oqhiw6);
assign Oqhiw6 = (W5fov6 ? Crhiw6 : Vqhiw6);
assign Xs78v6 = (W5fov6 ? Pjb7z6[15] : Wjeiw6);
assign Qs78v6 = (W5fov6 ? Pjb7z6[14] : Pjeiw6);
assign Js78v6 = (W5fov6 ? Pjb7z6[13] : Dkeiw6);
assign Cs78v6 = (W5fov6 ? Pjb7z6[12] : Jrhiw6);
assign Vr78v6 = (Xrhiw6 ? Qrhiw6 : Jke7v6);
assign Qrhiw6 = (~(K2adt6 | W2adt6));
assign Or78v6 = (W5fov6 ? Pjb7z6[11] : A62iw6);
assign Hr78v6 = (W5fov6 ? Pjb7z6[10] : O62iw6);
assign Ar78v6 = (W5fov6 ? Pjb7z6[9] : V62iw6);
assign Tq78v6 = (W5fov6 ? Pjb7z6[8] : C72iw6);
assign Mq78v6 = (W5fov6 ? Pjb7z6[7] : J72iw6);
assign Fq78v6 = (W5fov6 ? Pjb7z6[6] : Q72iw6);
assign Yp78v6 = (W5fov6 ? Pjb7z6[5] : X72iw6);
assign W5fov6 = (!Sdo7v6);
assign Rp78v6 = (Sdo7v6 ? E82iw6 : Pjb7z6[4]);
assign Kp78v6 = (Sdo7v6 ? L82iw6 : Pjb7z6[3]);
assign Dp78v6 = (Lshiw6 ? Eshiw6 : Xu67v6);
assign Lshiw6 = (Sshiw6 & L877v6);
assign Sshiw6 = (Zshiw6 & Gthiw6);
assign Wo78v6 = (Nthiw6 ? U42nv6 : Iy1nz6[0]);
assign Po78v6 = (Nthiw6 ? P52nv6 : Gie7v6);
assign Io78v6 = (Nthiw6 ? B52nv6 : Iy1nz6[1]);
assign Nthiw6 = (Uthiw6 & Buhiw6);
assign Uthiw6 = (Iuhiw6 & Puhiw6);
assign Bo78v6 = (Wuhiw6 ? Pk1nz6[0] : U42nv6);
assign Un78v6 = (~(Nyd7v6 ^ Wuhiw6));
assign Nn78v6 = (Wuhiw6 ? Pk1nz6[12] : Emhov6);
assign Gn78v6 = (Wuhiw6 ? Pk1nz6[11] : Dz6iw6);
assign Zm78v6 = (Wuhiw6 ? Pk1nz6[10] : H17iw6);
assign Sm78v6 = (Wuhiw6 ? Pk1nz6[9] : J27iw6);
assign Lm78v6 = (Wuhiw6 ? Pk1nz6[8] : U47iw6);
assign Wuhiw6 = (!Dvhiw6);
assign Em78v6 = (Dvhiw6 ? R62nv6 : Pk1nz6[7]);
assign Xl78v6 = (Dvhiw6 ? K62nv6 : Pk1nz6[6]);
assign Ql78v6 = (Dvhiw6 ? D62nv6 : Pk1nz6[5]);
assign Jl78v6 = (Dvhiw6 ? W52nv6 : Pk1nz6[4]);
assign Cl78v6 = (Dvhiw6 ? P52nv6 : Pk1nz6[3]);
assign Vk78v6 = (Dvhiw6 ? I52nv6 : Pk1nz6[2]);
assign Ok78v6 = (Dvhiw6 ? B52nv6 : Pk1nz6[1]);
assign Dvhiw6 = (Kvhiw6 & Rvhiw6);
assign Kvhiw6 = (Yvhiw6 & Iuhiw6);
assign Hk78v6 = (Fwhiw6 ? Nl1nz6[0] : U42nv6);
assign Ak78v6 = (Fwhiw6 ? Nl1nz6[1] : B52nv6);
assign Fwhiw6 = (~(Rvhiw6 & Mwhiw6));
assign Tj78v6 = (~(Twhiw6 & Axhiw6));
assign Axhiw6 = (~(Hxhiw6 & Oxhiw6));
assign Oxhiw6 = (Vxhiw6 & Cyhiw6);
assign Cyhiw6 = (Jyhiw6 & Qyhiw6);
assign Qyhiw6 = (~(Td2nz6[8] | Td2nz6[9]));
assign Jyhiw6 = (~(Td2nz6[6] | Td2nz6[7]));
assign Vxhiw6 = (Xyhiw6 & Ezhiw6);
assign Xyhiw6 = (~(Td2nz6[4] | Td2nz6[5]));
assign Hxhiw6 = (Lzhiw6 & Szhiw6);
assign Szhiw6 = (Zzhiw6 & G0iiw6);
assign Zzhiw6 = (~(Td2nz6[1] | Td2nz6[2]));
assign Lzhiw6 = (N0iiw6 & U0iiw6);
assign N0iiw6 = (~(Td2nz6[10] | Td2nz6[11]));
assign Mj78v6 = (~(B1iiw6 & I1iiw6));
assign I1iiw6 = (~(Tpf7v6 & P1iiw6));
assign B1iiw6 = (~(W1iiw6 & Td2nz6[0]));
assign Fj78v6 = (~(D2iiw6 & K2iiw6));
assign K2iiw6 = (~(Jof7v6 & P1iiw6));
assign D2iiw6 = (~(W1iiw6 & Td2nz6[1]));
assign Yi78v6 = (~(R2iiw6 & Y2iiw6));
assign Y2iiw6 = (~(Zmf7v6 & P1iiw6));
assign R2iiw6 = (~(W1iiw6 & Td2nz6[2]));
assign Ri78v6 = (~(F3iiw6 & M3iiw6));
assign M3iiw6 = (~(Plf7v6 & P1iiw6));
assign F3iiw6 = (~(W1iiw6 & Td2nz6[3]));
assign Ki78v6 = (~(T3iiw6 & A4iiw6));
assign A4iiw6 = (~(Fkf7v6 & P1iiw6));
assign T3iiw6 = (~(W1iiw6 & Td2nz6[4]));
assign Di78v6 = (~(H4iiw6 & O4iiw6));
assign O4iiw6 = (~(Vif7v6 & P1iiw6));
assign H4iiw6 = (~(W1iiw6 & Td2nz6[5]));
assign Wh78v6 = (~(V4iiw6 & C5iiw6));
assign C5iiw6 = (~(Lhf7v6 & P1iiw6));
assign V4iiw6 = (~(W1iiw6 & Td2nz6[6]));
assign Ph78v6 = (~(J5iiw6 & Q5iiw6));
assign Q5iiw6 = (~(Bgf7v6 & P1iiw6));
assign J5iiw6 = (~(W1iiw6 & Td2nz6[7]));
assign Ih78v6 = (~(X5iiw6 & E6iiw6));
assign E6iiw6 = (~(Ref7v6 & P1iiw6));
assign X5iiw6 = (~(W1iiw6 & Td2nz6[8]));
assign Bh78v6 = (~(L6iiw6 & S6iiw6));
assign S6iiw6 = (~(Hdf7v6 & P1iiw6));
assign L6iiw6 = (~(W1iiw6 & Td2nz6[9]));
assign Ug78v6 = (~(Z6iiw6 & G7iiw6));
assign G7iiw6 = (~(Xbf7v6 & P1iiw6));
assign Z6iiw6 = (~(W1iiw6 & Td2nz6[10]));
assign Ng78v6 = (~(N7iiw6 & U7iiw6));
assign U7iiw6 = (~(Naf7v6 & P1iiw6));
assign N7iiw6 = (~(W1iiw6 & Td2nz6[11]));
assign Gg78v6 = (~(B8iiw6 & I8iiw6));
assign I8iiw6 = (~(D9f7v6 & P1iiw6));
assign P1iiw6 = (P8iiw6 & W8iiw6);
assign P8iiw6 = (D9iiw6 & K9iiw6);
assign K9iiw6 = (!W1iiw6);
assign D9iiw6 = (~(R9iiw6 & Y9iiw6));
assign Y9iiw6 = (Faiiw6 & Maiiw6);
assign Maiiw6 = (Taiiw6 & Abiiw6);
assign Abiiw6 = (Hbiiw6 & Obiiw6);
assign Obiiw6 = (Pk1nz6[0] ^ U0iiw6);
assign U0iiw6 = (!Td2nz6[0]);
assign Hbiiw6 = (~(Pk1nz6[10] ^ Td2nz6[10]));
assign Taiiw6 = (Vbiiw6 & Cciiw6);
assign Cciiw6 = (~(Pk1nz6[11] ^ Td2nz6[11]));
assign Vbiiw6 = (Pk1nz6[12] ^ G0iiw6);
assign G0iiw6 = (!Td2nz6[12]);
assign Faiiw6 = (Jciiw6 & Qciiw6);
assign Qciiw6 = (~(Pk1nz6[2] ^ Td2nz6[2]));
assign Jciiw6 = (Xciiw6 & Ediiw6);
assign Ediiw6 = (Pk1nz6[3] ^ Ezhiw6);
assign Ezhiw6 = (!Td2nz6[3]);
assign Xciiw6 = (~(Pk1nz6[1] ^ Td2nz6[1]));
assign R9iiw6 = (Ldiiw6 & Sdiiw6);
assign Sdiiw6 = (Zdiiw6 & Geiiw6);
assign Geiiw6 = (~(Pk1nz6[5] ^ Td2nz6[5]));
assign Zdiiw6 = (Neiiw6 & Ueiiw6);
assign Ueiiw6 = (~(Pk1nz6[6] ^ Td2nz6[6]));
assign Neiiw6 = (~(Pk1nz6[4] ^ Td2nz6[4]));
assign Ldiiw6 = (Bfiiw6 & Ifiiw6);
assign Ifiiw6 = (~(Pk1nz6[8] ^ Td2nz6[8]));
assign Bfiiw6 = (Pfiiw6 & Wfiiw6);
assign Wfiiw6 = (~(Pk1nz6[9] ^ Td2nz6[9]));
assign Pfiiw6 = (~(Pk1nz6[7] ^ Td2nz6[7]));
assign B8iiw6 = (~(W1iiw6 & Td2nz6[12]));
assign W1iiw6 = (Dgiiw6 & W8iiw6);
assign W8iiw6 = (Fhh7v6 ^ Drf7v6);
assign Dgiiw6 = (M81nv6 & Vuf7v6);
assign Zf78v6 = (Kgiiw6 ? B52nv6 : Lge7v6);
assign Kgiiw6 = (Buhiw6 & Rgiiw6);
assign Buhiw6 = (Rvhiw6 & J02nz6[2]);
assign Sf78v6 = (Ygiiw6 ? U42nv6 : Hce7v6);
assign Ygiiw6 = (Fhiiw6 & Rvhiw6);
assign Fhiiw6 = (Mhiiw6 & Thiiw6);
assign Lf78v6 = (Aiiiw6 ? Eee7v6 : U42nv6);
assign Ef78v6 = (Aiiiw6 ? Hae7v6 : B52nv6);
assign Aiiiw6 = (~(Rvhiw6 & Hiiiw6));
assign Xe78v6 = (~(Oiiiw6 & Viiiw6));
assign Viiiw6 = (~(Jw1nz6[0] & Cjiiw6));
assign Cjiiw6 = (~(Jjiiw6 & U42nv6));
assign Oiiiw6 = (~(Qjiiw6 & U42nv6));
assign Qe78v6 = (~(Xjiiw6 & Ekiiw6));
assign Ekiiw6 = (~(Jw1nz6[1] & Lkiiw6));
assign Lkiiw6 = (~(Jjiiw6 & B52nv6));
assign Xjiiw6 = (~(Qjiiw6 & B52nv6));
assign Je78v6 = (~(Skiiw6 & Zkiiw6));
assign Zkiiw6 = (~(Jw1nz6[2] & Gliiw6));
assign Gliiw6 = (~(Jjiiw6 & I52nv6));
assign Skiiw6 = (~(Qjiiw6 & I52nv6));
assign Ce78v6 = (~(Nliiw6 & Uliiw6));
assign Uliiw6 = (~(Jw1nz6[3] & Bmiiw6));
assign Bmiiw6 = (~(Jjiiw6 & P52nv6));
assign Nliiw6 = (~(Qjiiw6 & P52nv6));
assign Qjiiw6 = (Jjiiw6 & Imiiw6);
assign Jjiiw6 = (Rvhiw6 & Pmiiw6);
assign Rvhiw6 = (Wmiiw6 & Xrhiw6);
assign Xrhiw6 = (Dniiw6 & Kniiw6);
assign Wmiiw6 = (K2adt6 & W2adt6);
assign Vd78v6 = (~(Rniiw6 & Yniiw6));
assign Yniiw6 = (~(Xc5ov6 & Sk5ov6));
assign Sk5ov6 = (!Foiiw6);
assign Foiiw6 = (U81nz6[2] ? Toiiw6 : Moiiw6);
assign Toiiw6 = (Nl5ov6 & Ld5ov6);
assign Moiiw6 = (~(Ul5ov6 & Nl5ov6));
assign Xc5ov6 = (Apiiw6 & Cc5ov6);
assign Rniiw6 = (~(U81nz6[2] & Sd5ov6));
assign Sd5ov6 = (!Apiiw6);
assign Od78v6 = (~(Hpiiw6 & Opiiw6));
assign Opiiw6 = (~(Vpiiw6 & Hcget6));
assign Vpiiw6 = (U3cet6 & Cqiiw6);
assign Hpiiw6 = (~(Jd47v6 & Jqiiw6));
assign Jqiiw6 = (Hcget6 | Qqiiw6);
assign Qqiiw6 = (K3jnv6 & Byeov6);
assign Hd78v6 = (~(Xqiiw6 & Eriiw6));
assign Eriiw6 = (~(Fjb7z6[0] & Lriiw6));
assign Xqiiw6 = (~(Sriiw6 & Zriiw6));
assign Ad78v6 = (~(Gsiiw6 & Nsiiw6));
assign Nsiiw6 = (~(Oc47v6 & Usiiw6));
assign Tc78v6 = (~(Btiiw6 & Itiiw6));
assign Itiiw6 = (~(O1fov6 & RXEV));
assign Btiiw6 = (~(Ei77z6 & V1fov6));
assign Mc78v6 = (~(Ptiiw6 & Wtiiw6));
assign Wtiiw6 = (~(INTISR[62] & O1fov6));
assign Ptiiw6 = (~(C797z6 & V1fov6));
assign Fc78v6 = (~(Duiiw6 & Kuiiw6));
assign Kuiiw6 = (~(INTISR[61] & O1fov6));
assign Duiiw6 = (~(K797z6 & V1fov6));
assign Yb78v6 = (~(Ruiiw6 & Yuiiw6));
assign Yuiiw6 = (~(INTISR[60] & O1fov6));
assign Ruiiw6 = (~(S797z6 & V1fov6));
assign Rb78v6 = (~(Fviiw6 & Mviiw6));
assign Mviiw6 = (~(INTISR[59] & O1fov6));
assign Fviiw6 = (~(A897z6 & V1fov6));
assign Kb78v6 = (~(Tviiw6 & Awiiw6));
assign Awiiw6 = (~(INTISR[58] & O1fov6));
assign Tviiw6 = (~(I897z6 & V1fov6));
assign Db78v6 = (~(Hwiiw6 & Owiiw6));
assign Owiiw6 = (~(INTISR[57] & O1fov6));
assign Hwiiw6 = (~(Q897z6 & V1fov6));
assign Wa78v6 = (~(Vwiiw6 & Cxiiw6));
assign Cxiiw6 = (~(INTISR[56] & O1fov6));
assign Vwiiw6 = (~(Y897z6 & V1fov6));
assign Pa78v6 = (~(Jxiiw6 & Qxiiw6));
assign Qxiiw6 = (~(INTISR[55] & O1fov6));
assign Jxiiw6 = (~(G997z6 & V1fov6));
assign Ia78v6 = (~(Xxiiw6 & Eyiiw6));
assign Eyiiw6 = (~(INTISR[54] & O1fov6));
assign Xxiiw6 = (~(O997z6 & V1fov6));
assign Ba78v6 = (~(Lyiiw6 & Syiiw6));
assign Syiiw6 = (~(INTISR[53] & O1fov6));
assign Lyiiw6 = (~(W997z6 & V1fov6));
assign U978v6 = (~(Zyiiw6 & Gziiw6));
assign Gziiw6 = (~(INTISR[52] & O1fov6));
assign Zyiiw6 = (~(Ea97z6 & V1fov6));
assign N978v6 = (~(Nziiw6 & Uziiw6));
assign Uziiw6 = (~(INTISR[51] & O1fov6));
assign Nziiw6 = (~(Ma97z6 & V1fov6));
assign G978v6 = (~(B0jiw6 & I0jiw6));
assign I0jiw6 = (~(INTISR[50] & O1fov6));
assign B0jiw6 = (~(Ua97z6 & V1fov6));
assign Z878v6 = (~(P0jiw6 & W0jiw6));
assign W0jiw6 = (~(INTISR[49] & O1fov6));
assign P0jiw6 = (~(Cb97z6 & V1fov6));
assign S878v6 = (~(D1jiw6 & K1jiw6));
assign K1jiw6 = (~(INTISR[48] & O1fov6));
assign D1jiw6 = (~(Kb97z6 & V1fov6));
assign L878v6 = (~(R1jiw6 & Y1jiw6));
assign Y1jiw6 = (~(INTISR[47] & O1fov6));
assign R1jiw6 = (~(Sb97z6 & V1fov6));
assign E878v6 = (~(F2jiw6 & M2jiw6));
assign M2jiw6 = (~(INTISR[46] & O1fov6));
assign F2jiw6 = (~(Ac97z6 & V1fov6));
assign X778v6 = (~(T2jiw6 & A3jiw6));
assign A3jiw6 = (~(INTISR[45] & O1fov6));
assign T2jiw6 = (~(Ic97z6 & V1fov6));
assign Q778v6 = (~(H3jiw6 & O3jiw6));
assign O3jiw6 = (~(INTISR[44] & O1fov6));
assign H3jiw6 = (~(Qc97z6 & V1fov6));
assign J778v6 = (~(V3jiw6 & C4jiw6));
assign C4jiw6 = (~(INTISR[43] & O1fov6));
assign V3jiw6 = (~(Yc97z6 & V1fov6));
assign C778v6 = (~(J4jiw6 & Q4jiw6));
assign Q4jiw6 = (~(INTISR[42] & O1fov6));
assign J4jiw6 = (~(Gd97z6 & V1fov6));
assign V678v6 = (~(X4jiw6 & E5jiw6));
assign E5jiw6 = (~(INTISR[41] & O1fov6));
assign X4jiw6 = (~(Od97z6 & V1fov6));
assign O678v6 = (~(L5jiw6 & S5jiw6));
assign S5jiw6 = (~(INTISR[40] & O1fov6));
assign L5jiw6 = (~(Wd97z6 & V1fov6));
assign H678v6 = (~(Z5jiw6 & G6jiw6));
assign G6jiw6 = (~(INTISR[39] & O1fov6));
assign Z5jiw6 = (~(Ee97z6 & V1fov6));
assign A678v6 = (~(N6jiw6 & U6jiw6));
assign U6jiw6 = (~(INTISR[38] & O1fov6));
assign N6jiw6 = (~(Me97z6 & V1fov6));
assign T578v6 = (~(B7jiw6 & I7jiw6));
assign I7jiw6 = (~(INTISR[37] & O1fov6));
assign B7jiw6 = (~(Ue97z6 & V1fov6));
assign M578v6 = (~(P7jiw6 & W7jiw6));
assign W7jiw6 = (~(INTISR[36] & O1fov6));
assign P7jiw6 = (~(Cf97z6 & V1fov6));
assign F578v6 = (~(D8jiw6 & K8jiw6));
assign K8jiw6 = (~(INTISR[35] & O1fov6));
assign D8jiw6 = (~(Kf97z6 & V1fov6));
assign Y478v6 = (~(R8jiw6 & Y8jiw6));
assign Y8jiw6 = (~(INTISR[34] & O1fov6));
assign R8jiw6 = (~(Sf97z6 & V1fov6));
assign R478v6 = (~(F9jiw6 & M9jiw6));
assign M9jiw6 = (~(INTISR[33] & O1fov6));
assign F9jiw6 = (~(Ag97z6 & V1fov6));
assign K478v6 = (~(T9jiw6 & Aajiw6));
assign Aajiw6 = (~(INTISR[32] & O1fov6));
assign T9jiw6 = (~(Ig97z6 & V1fov6));
assign D478v6 = (~(Hajiw6 & Oajiw6));
assign Oajiw6 = (~(INTISR[31] & O1fov6));
assign Hajiw6 = (~(Qg97z6 & V1fov6));
assign W378v6 = (~(Vajiw6 & Cbjiw6));
assign Cbjiw6 = (~(INTISR[30] & O1fov6));
assign Vajiw6 = (~(Yg97z6 & V1fov6));
assign P378v6 = (~(Jbjiw6 & Qbjiw6));
assign Qbjiw6 = (~(INTISR[29] & O1fov6));
assign Jbjiw6 = (~(Gh97z6 & V1fov6));
assign I378v6 = (~(Xbjiw6 & Ecjiw6));
assign Ecjiw6 = (~(INTISR[28] & O1fov6));
assign Xbjiw6 = (~(Oh97z6 & V1fov6));
assign B378v6 = (~(Lcjiw6 & Scjiw6));
assign Scjiw6 = (~(INTISR[27] & O1fov6));
assign Lcjiw6 = (~(Wh97z6 & V1fov6));
assign U278v6 = (~(Zcjiw6 & Gdjiw6));
assign Gdjiw6 = (~(INTISR[26] & O1fov6));
assign Zcjiw6 = (~(Ei97z6 & V1fov6));
assign N278v6 = (~(Ndjiw6 & Udjiw6));
assign Udjiw6 = (~(INTISR[25] & O1fov6));
assign Ndjiw6 = (~(Mi97z6 & V1fov6));
assign G278v6 = (~(Bejiw6 & Iejiw6));
assign Iejiw6 = (~(INTISR[24] & O1fov6));
assign Bejiw6 = (~(Ui97z6 & V1fov6));
assign Z178v6 = (~(Pejiw6 & Wejiw6));
assign Wejiw6 = (~(INTISR[23] & O1fov6));
assign Pejiw6 = (~(Cj97z6 & V1fov6));
assign S178v6 = (~(Dfjiw6 & Kfjiw6));
assign Kfjiw6 = (~(INTISR[22] & O1fov6));
assign Dfjiw6 = (~(Kj97z6 & V1fov6));
assign L178v6 = (~(Rfjiw6 & Yfjiw6));
assign Yfjiw6 = (~(INTISR[21] & O1fov6));
assign Rfjiw6 = (~(Sj97z6 & V1fov6));
assign E178v6 = (~(Fgjiw6 & Mgjiw6));
assign Mgjiw6 = (~(INTISR[20] & O1fov6));
assign Fgjiw6 = (~(Ak97z6 & V1fov6));
assign X078v6 = (~(Tgjiw6 & Ahjiw6));
assign Ahjiw6 = (~(INTISR[19] & O1fov6));
assign Tgjiw6 = (~(Ik97z6 & V1fov6));
assign Q078v6 = (~(Hhjiw6 & Ohjiw6));
assign Ohjiw6 = (~(INTISR[18] & O1fov6));
assign Hhjiw6 = (~(Qk97z6 & V1fov6));
assign J078v6 = (~(Vhjiw6 & Cijiw6));
assign Cijiw6 = (~(INTISR[17] & O1fov6));
assign Vhjiw6 = (~(Yk97z6 & V1fov6));
assign C078v6 = (~(Jijiw6 & Qijiw6));
assign Qijiw6 = (~(INTISR[16] & O1fov6));
assign Jijiw6 = (~(Gl97z6 & V1fov6));
assign Vz68v6 = (~(Xijiw6 & Ejjiw6));
assign Ejjiw6 = (~(INTISR[15] & O1fov6));
assign Xijiw6 = (~(Ol97z6 & V1fov6));
assign Oz68v6 = (~(Ljjiw6 & Sjjiw6));
assign Sjjiw6 = (~(INTISR[14] & O1fov6));
assign Ljjiw6 = (~(Wl97z6 & V1fov6));
assign Hz68v6 = (~(Zjjiw6 & Gkjiw6));
assign Gkjiw6 = (~(INTISR[13] & O1fov6));
assign Zjjiw6 = (~(Em97z6 & V1fov6));
assign Az68v6 = (~(Nkjiw6 & Ukjiw6));
assign Ukjiw6 = (~(INTISR[12] & O1fov6));
assign Nkjiw6 = (~(Mm97z6 & V1fov6));
assign Ty68v6 = (~(Bljiw6 & Iljiw6));
assign Iljiw6 = (~(INTISR[11] & O1fov6));
assign Bljiw6 = (~(Um97z6 & V1fov6));
assign My68v6 = (~(Pljiw6 & Wljiw6));
assign Wljiw6 = (~(INTISR[10] & O1fov6));
assign Pljiw6 = (~(Cn97z6 & V1fov6));
assign Fy68v6 = (~(Dmjiw6 & Kmjiw6));
assign Kmjiw6 = (~(INTISR[9] & O1fov6));
assign Dmjiw6 = (~(Kn97z6 & V1fov6));
assign Yx68v6 = (~(Rmjiw6 & Ymjiw6));
assign Ymjiw6 = (~(INTISR[8] & O1fov6));
assign Rmjiw6 = (~(Sn97z6 & V1fov6));
assign Rx68v6 = (~(Fnjiw6 & Mnjiw6));
assign Mnjiw6 = (~(INTISR[7] & O1fov6));
assign Fnjiw6 = (~(Ao97z6 & V1fov6));
assign Kx68v6 = (~(Tnjiw6 & Aojiw6));
assign Aojiw6 = (~(INTISR[6] & O1fov6));
assign Tnjiw6 = (~(Io97z6 & V1fov6));
assign Dx68v6 = (~(Hojiw6 & Oojiw6));
assign Oojiw6 = (~(INTISR[5] & O1fov6));
assign Hojiw6 = (~(Qo97z6 & V1fov6));
assign Ww68v6 = (~(Vojiw6 & Cpjiw6));
assign Cpjiw6 = (~(INTISR[4] & O1fov6));
assign Vojiw6 = (~(Yo97z6 & V1fov6));
assign Pw68v6 = (~(Jpjiw6 & Qpjiw6));
assign Qpjiw6 = (~(INTISR[3] & O1fov6));
assign Jpjiw6 = (~(Gp97z6 & V1fov6));
assign Iw68v6 = (~(Xpjiw6 & Eqjiw6));
assign Eqjiw6 = (~(INTISR[2] & O1fov6));
assign Xpjiw6 = (~(Op97z6 & V1fov6));
assign Bw68v6 = (~(Lqjiw6 & Sqjiw6));
assign Sqjiw6 = (~(INTISR[1] & O1fov6));
assign Lqjiw6 = (~(Wp97z6 & V1fov6));
assign Uv68v6 = (~(Zqjiw6 & Grjiw6));
assign Grjiw6 = (~(INTISR[0] & O1fov6));
assign Zqjiw6 = (~(Eq97z6 & V1fov6));
assign Nv68v6 = (~(Nrjiw6 & Urjiw6));
assign Urjiw6 = (~(EDBGRQ & O1fov6));
assign Nrjiw6 = (~(Mq97z6 & V1fov6));
assign Gv68v6 = (~(Bsjiw6 & Isjiw6));
assign Isjiw6 = (~(INTNMI & O1fov6));
assign O1fov6 = (Psjiw6 & Usiiw6);
assign Bsjiw6 = (~(Uq97z6 & V1fov6));
assign V1fov6 = (~(M6bdt6 & Psjiw6));
assign Psjiw6 = (Oc47v6 | Sriiw6);
assign Zu68v6 = (~(Wsjiw6 & Dtjiw6));
assign Wsjiw6 = (G7bdt6 & U42nv6);
assign Su68v6 = (Dtjiw6 ? I52nv6 : SYSRESETREQ);
assign Lu68v6 = (Dtjiw6 ? H17iw6 : Hsi7z6[2]);
assign Eu68v6 = (Dtjiw6 ? J27iw6 : Hsi7z6[1]);
assign Xt68v6 = (Dtjiw6 ? U47iw6 : Hsi7z6[0]);
assign Qt68v6 = (Ktjiw6 ? Z0iov6 : Pnb7z6[15]);
assign Jt68v6 = (Ktjiw6 ? U47iw6 : Qti7z6[8]);
assign Ct68v6 = (Ktjiw6 ? J27iw6 : Qti7z6[9]);
assign Vs68v6 = (Ktjiw6 ? H17iw6 : Pnb7z6[10]);
assign Os68v6 = (Ktjiw6 ? Dz6iw6 : Pnb7z6[11]);
assign Hs68v6 = (Ktjiw6 ? Emhov6 : Pnb7z6[12]);
assign As68v6 = (Ktjiw6 ? Guhov6 : Pnb7z6[13]);
assign Tr68v6 = (Ktjiw6 ? Bk6iw6 : Pnb7z6[14]);
assign Ktjiw6 = (Rtjiw6 & Bqi7z6[1]);
assign Mr68v6 = (Ytjiw6 ? Cx4iw6 : Pnb7z6[23]);
assign Fr68v6 = (Ytjiw6 ? Is5iw6 : Pnb7z6[16]);
assign Yq68v6 = (Ytjiw6 ? Gr5iw6 : Pnb7z6[17]);
assign Rq68v6 = (Ytjiw6 ? Jp5iw6 : Pnb7z6[18]);
assign Kq68v6 = (Ytjiw6 ? Mn5iw6 : Pnb7z6[19]);
assign Dq68v6 = (Ytjiw6 ? Bl5iw6 : Pnb7z6[20]);
assign Wp68v6 = (Ytjiw6 ? Ej5iw6 : Pnb7z6[21]);
assign Pp68v6 = (Ytjiw6 ? D85iw6 : Pnb7z6[22]);
assign Ytjiw6 = (Rtjiw6 & Bqi7z6[2]);
assign Ip68v6 = (Fujiw6 ? X0hov6 : Pnb7z6[31]);
assign Bp68v6 = (Fujiw6 ? Wf4iw6 : Pnb7z6[24]);
assign Uo68v6 = (Fujiw6 ? Iklov6 : Pnb7z6[25]);
assign No68v6 = (Fujiw6 ? E64iw6 : Pnb7z6[26]);
assign Go68v6 = (Fujiw6 ? H44iw6 : Pnb7z6[27]);
assign Zn68v6 = (Fujiw6 ? W14iw6 : Pnb7z6[28]);
assign Sn68v6 = (Fujiw6 ? Zz3iw6 : Pnb7z6[29]);
assign Ln68v6 = (Fujiw6 ? Ro3iw6 : Pnb7z6[30]);
assign Fujiw6 = (Rtjiw6 & Bqi7z6[3]);
assign En68v6 = (~(Mujiw6 & Tujiw6));
assign Tujiw6 = (~(Qti7z6[7] & Avjiw6));
assign Avjiw6 = (~(Rtjiw6 & Bqi7z6[0]));
assign Mujiw6 = (~(Rtjiw6 & O87iw6));
assign Rtjiw6 = (Hvjiw6 & T68iw6);
assign Xm68v6 = (!Ovjiw6);
assign Ovjiw6 = (Kdmov6 ? I497z6 : Vvjiw6);
assign Qm68v6 = (~(Cwjiw6 & Jwjiw6));
assign Jwjiw6 = (~(Qwjiw6 & Ysdiw6));
assign Cwjiw6 = (~(Kdmov6 & Rnm7z6[0]));
assign Jm68v6 = (~(Xwjiw6 & Exjiw6));
assign Exjiw6 = (~(Lxjiw6 & Qwjiw6));
assign Xwjiw6 = (~(Kdmov6 & Rnm7z6[1]));
assign Cm68v6 = (~(Sxjiw6 & Zxjiw6));
assign Zxjiw6 = (~(Qwjiw6 & Gyjiw6));
assign Qwjiw6 = (Vvjiw6 & Mdonv6);
assign Vvjiw6 = (Nyjiw6 & Uyjiw6);
assign Uyjiw6 = (~(Bzjiw6 & I2yet6));
assign Nyjiw6 = (Izjiw6 & Sgonv6);
assign Izjiw6 = (~(Lgonv6 & Zgonv6));
assign Sxjiw6 = (~(Kdmov6 & Rnm7z6[2]));
assign Kdmov6 = (!Mdonv6);
assign Vl68v6 = (Jalov6 & Pzjiw6);
assign Pzjiw6 = (~(Wzjiw6 & D0kiw6));
assign D0kiw6 = (~(K0kiw6 & Woyet6));
assign K0kiw6 = (R0kiw6 & Y0kiw6);
assign R0kiw6 = (~(F1kiw6 & Znn7z6[0]));
assign F1kiw6 = (!M1kiw6);
assign Wzjiw6 = (~(T1kiw6 & A2kiw6));
assign T1kiw6 = (~(H2kiw6 | M4xnv6));
assign Jalov6 = (~(L1bdt6 | Qteet6));
assign Ol68v6 = (~(O2kiw6 & V2kiw6));
assign V2kiw6 = (~(C3kiw6 & J3kiw6));
assign C3kiw6 = (Ebdiw6 & Q3kiw6);
assign O2kiw6 = (~(Zy1ft6 & X3kiw6));
assign X3kiw6 = (~(E4kiw6 & J3kiw6));
assign E4kiw6 = (Q3kiw6 & B52nv6);
assign Hl68v6 = (L4kiw6 ? K62nv6 : Ugtet6);
assign Al68v6 = (L4kiw6 ? R62nv6 : Tetet6);
assign Tk68v6 = (L4kiw6 ? U47iw6 : Sctet6);
assign Mk68v6 = (L4kiw6 ? J27iw6 : Ratet6);
assign Fk68v6 = (L4kiw6 ? H17iw6 : Q8tet6);
assign Yj68v6 = (L4kiw6 ? Dz6iw6 : P6tet6);
assign Rj68v6 = (L4kiw6 ? Emhov6 : O4tet6);
assign Kj68v6 = (L4kiw6 ? Guhov6 : N2tet6);
assign Dj68v6 = (L4kiw6 ? Bk6iw6 : M0tet6);
assign Wi68v6 = (L4kiw6 ? Z0iov6 : Lyset6);
assign Pi68v6 = (L4kiw6 ? Is5iw6 : Kwset6);
assign Ii68v6 = (L4kiw6 ? Gr5iw6 : Juset6);
assign Bi68v6 = (L4kiw6 ? Jp5iw6 : Isset6);
assign Uh68v6 = (L4kiw6 ? Mn5iw6 : Hqset6);
assign Nh68v6 = (L4kiw6 ? Bl5iw6 : Goset6);
assign Gh68v6 = (L4kiw6 ? Ej5iw6 : Fmset6);
assign Zg68v6 = (L4kiw6 ? D85iw6 : Ekset6);
assign Sg68v6 = (L4kiw6 ? Cx4iw6 : Diset6);
assign Lg68v6 = (L4kiw6 ? Wf4iw6 : Cgset6);
assign Eg68v6 = (L4kiw6 ? Iklov6 : Beset6);
assign Xf68v6 = (L4kiw6 ? E64iw6 : Acset6);
assign Qf68v6 = (L4kiw6 ? H44iw6 : Z9set6);
assign Jf68v6 = (L4kiw6 ? W14iw6 : Y7set6);
assign Cf68v6 = (L4kiw6 ? D62nv6 : Vitet6);
assign L4kiw6 = (J3kiw6 & S4kiw6);
assign Ve68v6 = (Z4kiw6 ? P52nv6 : W3p7z6[3]);
assign Oe68v6 = (Z4kiw6 ? W52nv6 : W3p7z6[4]);
assign He68v6 = (Z4kiw6 ? D62nv6 : W3p7z6[5]);
assign Ae68v6 = (Z4kiw6 ? K62nv6 : W3p7z6[6]);
assign Td68v6 = (Z4kiw6 ? R62nv6 : W3p7z6[7]);
assign Md68v6 = (Z4kiw6 ? U47iw6 : W3p7z6[8]);
assign Fd68v6 = (Z4kiw6 ? J27iw6 : W3p7z6[9]);
assign Yc68v6 = (Z4kiw6 ? H17iw6 : W3p7z6[10]);
assign Rc68v6 = (Z4kiw6 ? Dz6iw6 : W3p7z6[11]);
assign Kc68v6 = (Z4kiw6 ? Emhov6 : W3p7z6[12]);
assign Dc68v6 = (Z4kiw6 ? Guhov6 : W3p7z6[13]);
assign Wb68v6 = (Z4kiw6 ? Bk6iw6 : W3p7z6[14]);
assign Pb68v6 = (Z4kiw6 ? Z0iov6 : W3p7z6[15]);
assign Ib68v6 = (Z4kiw6 ? Is5iw6 : W3p7z6[16]);
assign Bb68v6 = (Z4kiw6 ? Gr5iw6 : W3p7z6[17]);
assign Ua68v6 = (Z4kiw6 ? Jp5iw6 : W3p7z6[18]);
assign Na68v6 = (Z4kiw6 ? Mn5iw6 : W3p7z6[19]);
assign Ga68v6 = (Z4kiw6 ? Bl5iw6 : W3p7z6[20]);
assign Z968v6 = (Z4kiw6 ? Ej5iw6 : W3p7z6[21]);
assign S968v6 = (Z4kiw6 ? D85iw6 : W3p7z6[22]);
assign L968v6 = (Z4kiw6 ? Cx4iw6 : W3p7z6[23]);
assign E968v6 = (Z4kiw6 ? Wf4iw6 : W3p7z6[24]);
assign X868v6 = (Z4kiw6 ? Iklov6 : W3p7z6[25]);
assign Q868v6 = (Z4kiw6 ? E64iw6 : W3p7z6[26]);
assign J868v6 = (Z4kiw6 ? H44iw6 : W3p7z6[27]);
assign C868v6 = (Z4kiw6 ? W14iw6 : W3p7z6[28]);
assign V768v6 = (Z4kiw6 ? Ro3iw6 : Nw1ft6);
assign O768v6 = (Z4kiw6 ? X0hov6 : Tx1ft6);
assign H768v6 = (Z4kiw6 ? I52nv6 : W3p7z6[2]);
assign A768v6 = (Z4kiw6 ? U42nv6 : Iv1ft6);
assign Z4kiw6 = (J3kiw6 & G5kiw6);
assign T668v6 = (N5kiw6 ? P52nv6 : T2p7z6[3]);
assign M668v6 = (N5kiw6 ? W52nv6 : T2p7z6[4]);
assign F668v6 = (N5kiw6 ? D62nv6 : T2p7z6[5]);
assign Y568v6 = (N5kiw6 ? K62nv6 : T2p7z6[6]);
assign R568v6 = (N5kiw6 ? R62nv6 : T2p7z6[7]);
assign K568v6 = (N5kiw6 ? U47iw6 : T2p7z6[8]);
assign D568v6 = (N5kiw6 ? J27iw6 : T2p7z6[9]);
assign W468v6 = (N5kiw6 ? H17iw6 : T2p7z6[10]);
assign P468v6 = (N5kiw6 ? Dz6iw6 : T2p7z6[11]);
assign I468v6 = (N5kiw6 ? Emhov6 : T2p7z6[12]);
assign B468v6 = (N5kiw6 ? Guhov6 : T2p7z6[13]);
assign U368v6 = (N5kiw6 ? Bk6iw6 : T2p7z6[14]);
assign N368v6 = (N5kiw6 ? Z0iov6 : T2p7z6[15]);
assign G368v6 = (N5kiw6 ? Is5iw6 : T2p7z6[16]);
assign Z268v6 = (N5kiw6 ? Gr5iw6 : T2p7z6[17]);
assign S268v6 = (N5kiw6 ? Jp5iw6 : T2p7z6[18]);
assign L268v6 = (N5kiw6 ? Mn5iw6 : T2p7z6[19]);
assign E268v6 = (N5kiw6 ? Bl5iw6 : T2p7z6[20]);
assign X168v6 = (N5kiw6 ? Ej5iw6 : T2p7z6[21]);
assign Q168v6 = (N5kiw6 ? D85iw6 : T2p7z6[22]);
assign J168v6 = (N5kiw6 ? Cx4iw6 : T2p7z6[23]);
assign C168v6 = (N5kiw6 ? Wf4iw6 : T2p7z6[24]);
assign V068v6 = (N5kiw6 ? Iklov6 : T2p7z6[25]);
assign O068v6 = (N5kiw6 ? E64iw6 : T2p7z6[26]);
assign H068v6 = (N5kiw6 ? H44iw6 : T2p7z6[27]);
assign A068v6 = (N5kiw6 ? W14iw6 : T2p7z6[28]);
assign Tz58v6 = (N5kiw6 ? Ro3iw6 : Ws1ft6);
assign Mz58v6 = (N5kiw6 ? X0hov6 : Cu1ft6);
assign Fz58v6 = (N5kiw6 ? I52nv6 : T2p7z6[2]);
assign Yy58v6 = (N5kiw6 ? U42nv6 : Rr1ft6);
assign N5kiw6 = (J3kiw6 & U5kiw6);
assign Ry58v6 = (B6kiw6 ? P52nv6 : A0p7z6[1]);
assign Ky58v6 = (B6kiw6 ? W52nv6 : A0p7z6[2]);
assign Dy58v6 = (B6kiw6 ? D62nv6 : A0p7z6[3]);
assign Wx58v6 = (B6kiw6 ? K62nv6 : A0p7z6[4]);
assign Px58v6 = (B6kiw6 ? R62nv6 : A0p7z6[5]);
assign Ix58v6 = (B6kiw6 ? U47iw6 : A0p7z6[6]);
assign Bx58v6 = (B6kiw6 ? J27iw6 : A0p7z6[7]);
assign Uw58v6 = (B6kiw6 ? H17iw6 : A0p7z6[8]);
assign Nw58v6 = (B6kiw6 ? Dz6iw6 : A0p7z6[9]);
assign Gw58v6 = (B6kiw6 ? Emhov6 : A0p7z6[10]);
assign Zv58v6 = (B6kiw6 ? Guhov6 : A0p7z6[11]);
assign Sv58v6 = (B6kiw6 ? Bk6iw6 : A0p7z6[12]);
assign Lv58v6 = (B6kiw6 ? Z0iov6 : A0p7z6[13]);
assign Ev58v6 = (B6kiw6 ? Is5iw6 : A0p7z6[14]);
assign Xu58v6 = (B6kiw6 ? Gr5iw6 : A0p7z6[15]);
assign Qu58v6 = (B6kiw6 ? Jp5iw6 : A0p7z6[16]);
assign Ju58v6 = (B6kiw6 ? Mn5iw6 : A0p7z6[17]);
assign Cu58v6 = (B6kiw6 ? Bl5iw6 : A0p7z6[18]);
assign Vt58v6 = (B6kiw6 ? Ej5iw6 : A0p7z6[19]);
assign Ot58v6 = (B6kiw6 ? D85iw6 : A0p7z6[20]);
assign Ht58v6 = (B6kiw6 ? Cx4iw6 : A0p7z6[21]);
assign At58v6 = (B6kiw6 ? Wf4iw6 : A0p7z6[22]);
assign Ts58v6 = (B6kiw6 ? Iklov6 : A0p7z6[23]);
assign Ms58v6 = (B6kiw6 ? E64iw6 : A0p7z6[24]);
assign Fs58v6 = (B6kiw6 ? H44iw6 : A0p7z6[25]);
assign Yr58v6 = (B6kiw6 ? W14iw6 : A0p7z6[26]);
assign Rr58v6 = (B6kiw6 ? Ro3iw6 : I1p7z6[0]);
assign Kr58v6 = (B6kiw6 ? X0hov6 : I1p7z6[1]);
assign Dr58v6 = (B6kiw6 ? I52nv6 : A0p7z6[0]);
assign Wq58v6 = (B6kiw6 ? U42nv6 : Hq1ft6);
assign B6kiw6 = (J3kiw6 & I6kiw6);
assign Pq58v6 = (P6kiw6 ? P52nv6 : Hxo7z6[1]);
assign Iq58v6 = (P6kiw6 ? W52nv6 : Hxo7z6[2]);
assign Bq58v6 = (P6kiw6 ? D62nv6 : Hxo7z6[3]);
assign Up58v6 = (P6kiw6 ? K62nv6 : Hxo7z6[4]);
assign Np58v6 = (P6kiw6 ? R62nv6 : Hxo7z6[5]);
assign Gp58v6 = (P6kiw6 ? U47iw6 : Hxo7z6[6]);
assign Zo58v6 = (P6kiw6 ? J27iw6 : Hxo7z6[7]);
assign So58v6 = (P6kiw6 ? H17iw6 : Hxo7z6[8]);
assign Lo58v6 = (P6kiw6 ? Dz6iw6 : Hxo7z6[9]);
assign Eo58v6 = (P6kiw6 ? Emhov6 : Hxo7z6[10]);
assign Xn58v6 = (P6kiw6 ? Guhov6 : Hxo7z6[11]);
assign Qn58v6 = (P6kiw6 ? Bk6iw6 : Hxo7z6[12]);
assign Jn58v6 = (P6kiw6 ? Z0iov6 : Hxo7z6[13]);
assign Cn58v6 = (P6kiw6 ? Is5iw6 : Hxo7z6[14]);
assign Vm58v6 = (P6kiw6 ? Gr5iw6 : Hxo7z6[15]);
assign Om58v6 = (P6kiw6 ? Jp5iw6 : Hxo7z6[16]);
assign Hm58v6 = (P6kiw6 ? Mn5iw6 : Hxo7z6[17]);
assign Am58v6 = (P6kiw6 ? Bl5iw6 : Hxo7z6[18]);
assign Tl58v6 = (P6kiw6 ? Ej5iw6 : Hxo7z6[19]);
assign Ml58v6 = (P6kiw6 ? D85iw6 : Hxo7z6[20]);
assign Fl58v6 = (P6kiw6 ? Cx4iw6 : Hxo7z6[21]);
assign Yk58v6 = (P6kiw6 ? Wf4iw6 : Hxo7z6[22]);
assign Rk58v6 = (P6kiw6 ? Iklov6 : Hxo7z6[23]);
assign Kk58v6 = (P6kiw6 ? E64iw6 : Hxo7z6[24]);
assign Dk58v6 = (P6kiw6 ? H44iw6 : Hxo7z6[25]);
assign Wj58v6 = (P6kiw6 ? W14iw6 : Hxo7z6[26]);
assign Pj58v6 = (P6kiw6 ? Ro3iw6 : Pyo7z6[0]);
assign Ij58v6 = (P6kiw6 ? X0hov6 : Pyo7z6[1]);
assign Bj58v6 = (P6kiw6 ? I52nv6 : Hxo7z6[0]);
assign Ui58v6 = (P6kiw6 ? U42nv6 : Xo1ft6);
assign P6kiw6 = (J3kiw6 & W6kiw6);
assign Ni58v6 = (D7kiw6 ? P52nv6 : Ouo7z6[1]);
assign Gi58v6 = (D7kiw6 ? W52nv6 : Ouo7z6[2]);
assign Zh58v6 = (D7kiw6 ? D62nv6 : Ouo7z6[3]);
assign Sh58v6 = (D7kiw6 ? K62nv6 : Ouo7z6[4]);
assign Lh58v6 = (D7kiw6 ? R62nv6 : Ouo7z6[5]);
assign Eh58v6 = (D7kiw6 ? U47iw6 : Ouo7z6[6]);
assign Xg58v6 = (D7kiw6 ? J27iw6 : Ouo7z6[7]);
assign Qg58v6 = (D7kiw6 ? H17iw6 : Ouo7z6[8]);
assign Jg58v6 = (D7kiw6 ? Dz6iw6 : Ouo7z6[9]);
assign Cg58v6 = (D7kiw6 ? Emhov6 : Ouo7z6[10]);
assign Vf58v6 = (D7kiw6 ? Guhov6 : Ouo7z6[11]);
assign Of58v6 = (D7kiw6 ? Bk6iw6 : Ouo7z6[12]);
assign Hf58v6 = (D7kiw6 ? Z0iov6 : Ouo7z6[13]);
assign Af58v6 = (D7kiw6 ? Is5iw6 : Ouo7z6[14]);
assign Te58v6 = (D7kiw6 ? Gr5iw6 : Ouo7z6[15]);
assign Me58v6 = (D7kiw6 ? Jp5iw6 : Ouo7z6[16]);
assign Fe58v6 = (D7kiw6 ? Mn5iw6 : Ouo7z6[17]);
assign Yd58v6 = (D7kiw6 ? Bl5iw6 : Ouo7z6[18]);
assign Rd58v6 = (D7kiw6 ? Ej5iw6 : Ouo7z6[19]);
assign Kd58v6 = (D7kiw6 ? D85iw6 : Ouo7z6[20]);
assign Dd58v6 = (D7kiw6 ? Cx4iw6 : Ouo7z6[21]);
assign Wc58v6 = (D7kiw6 ? Wf4iw6 : Ouo7z6[22]);
assign Pc58v6 = (D7kiw6 ? Iklov6 : Ouo7z6[23]);
assign Ic58v6 = (D7kiw6 ? E64iw6 : Ouo7z6[24]);
assign Bc58v6 = (D7kiw6 ? H44iw6 : Ouo7z6[25]);
assign Ub58v6 = (D7kiw6 ? W14iw6 : Ouo7z6[26]);
assign Nb58v6 = (D7kiw6 ? Ro3iw6 : Wvo7z6[0]);
assign Gb58v6 = (D7kiw6 ? X0hov6 : Wvo7z6[1]);
assign Za58v6 = (D7kiw6 ? I52nv6 : Ouo7z6[0]);
assign Sa58v6 = (D7kiw6 ? U42nv6 : Nn1ft6);
assign D7kiw6 = (J3kiw6 & K7kiw6);
assign La58v6 = (R7kiw6 ? P52nv6 : Vro7z6[1]);
assign Ea58v6 = (R7kiw6 ? W52nv6 : Vro7z6[2]);
assign X958v6 = (R7kiw6 ? D62nv6 : Vro7z6[3]);
assign Q958v6 = (R7kiw6 ? K62nv6 : Vro7z6[4]);
assign J958v6 = (R7kiw6 ? R62nv6 : Vro7z6[5]);
assign C958v6 = (R7kiw6 ? U47iw6 : Vro7z6[6]);
assign V858v6 = (R7kiw6 ? J27iw6 : Vro7z6[7]);
assign O858v6 = (R7kiw6 ? H17iw6 : Vro7z6[8]);
assign H858v6 = (R7kiw6 ? Dz6iw6 : Vro7z6[9]);
assign A858v6 = (R7kiw6 ? Emhov6 : Vro7z6[10]);
assign T758v6 = (R7kiw6 ? Guhov6 : Vro7z6[11]);
assign M758v6 = (R7kiw6 ? Bk6iw6 : Vro7z6[12]);
assign F758v6 = (R7kiw6 ? Z0iov6 : Vro7z6[13]);
assign Y658v6 = (R7kiw6 ? Is5iw6 : Vro7z6[14]);
assign R658v6 = (R7kiw6 ? Gr5iw6 : Vro7z6[15]);
assign K658v6 = (R7kiw6 ? Jp5iw6 : Vro7z6[16]);
assign D658v6 = (R7kiw6 ? Mn5iw6 : Vro7z6[17]);
assign W558v6 = (R7kiw6 ? Bl5iw6 : Vro7z6[18]);
assign P558v6 = (R7kiw6 ? Ej5iw6 : Vro7z6[19]);
assign I558v6 = (R7kiw6 ? D85iw6 : Vro7z6[20]);
assign B558v6 = (R7kiw6 ? Cx4iw6 : Vro7z6[21]);
assign U458v6 = (R7kiw6 ? Wf4iw6 : Vro7z6[22]);
assign N458v6 = (R7kiw6 ? Iklov6 : Vro7z6[23]);
assign G458v6 = (R7kiw6 ? E64iw6 : Vro7z6[24]);
assign Z358v6 = (R7kiw6 ? H44iw6 : Vro7z6[25]);
assign S358v6 = (R7kiw6 ? W14iw6 : Vro7z6[26]);
assign L358v6 = (R7kiw6 ? Ro3iw6 : Dto7z6[0]);
assign E358v6 = (R7kiw6 ? X0hov6 : Dto7z6[1]);
assign X258v6 = (R7kiw6 ? I52nv6 : Vro7z6[0]);
assign Q258v6 = (R7kiw6 ? U42nv6 : Dm1ft6);
assign R7kiw6 = (J3kiw6 & Y7kiw6);
assign J258v6 = (F8kiw6 ? P52nv6 : Nqo7z6[1]);
assign C258v6 = (F8kiw6 ? W52nv6 : Nqo7z6[2]);
assign V158v6 = (F8kiw6 ? D62nv6 : Nqo7z6[3]);
assign O158v6 = (F8kiw6 ? K62nv6 : Nqo7z6[4]);
assign H158v6 = (F8kiw6 ? R62nv6 : Nqo7z6[5]);
assign A158v6 = (F8kiw6 ? U47iw6 : Nqo7z6[6]);
assign T058v6 = (F8kiw6 ? J27iw6 : Nqo7z6[7]);
assign M058v6 = (F8kiw6 ? H17iw6 : Nqo7z6[8]);
assign F058v6 = (F8kiw6 ? Dz6iw6 : Nqo7z6[9]);
assign Yz48v6 = (F8kiw6 ? Emhov6 : Nqo7z6[10]);
assign Rz48v6 = (F8kiw6 ? Guhov6 : Nqo7z6[11]);
assign Kz48v6 = (F8kiw6 ? Bk6iw6 : Nqo7z6[12]);
assign Dz48v6 = (F8kiw6 ? Z0iov6 : Nqo7z6[13]);
assign Wy48v6 = (F8kiw6 ? Is5iw6 : Nqo7z6[14]);
assign Py48v6 = (F8kiw6 ? Gr5iw6 : Nqo7z6[15]);
assign Iy48v6 = (F8kiw6 ? Jp5iw6 : Nqo7z6[16]);
assign By48v6 = (F8kiw6 ? Mn5iw6 : Nqo7z6[17]);
assign Ux48v6 = (F8kiw6 ? Bl5iw6 : Nqo7z6[18]);
assign Nx48v6 = (F8kiw6 ? Ej5iw6 : Nqo7z6[19]);
assign Gx48v6 = (F8kiw6 ? D85iw6 : Nqo7z6[20]);
assign Zw48v6 = (F8kiw6 ? Cx4iw6 : Nqo7z6[21]);
assign Sw48v6 = (F8kiw6 ? Wf4iw6 : Nqo7z6[22]);
assign Lw48v6 = (F8kiw6 ? Iklov6 : Nqo7z6[23]);
assign Ew48v6 = (F8kiw6 ? E64iw6 : Nqo7z6[24]);
assign Xv48v6 = (F8kiw6 ? H44iw6 : Nqo7z6[25]);
assign Qv48v6 = (F8kiw6 ? W14iw6 : Nqo7z6[26]);
assign Jv48v6 = (F8kiw6 ? I52nv6 : Nqo7z6[0]);
assign Cv48v6 = (F8kiw6 ? U42nv6 : Tk1ft6);
assign F8kiw6 = (J3kiw6 & M8kiw6);
assign Vu48v6 = (T8kiw6 ? Fpo7z6[1] : P52nv6);
assign Ou48v6 = (T8kiw6 ? Fpo7z6[2] : W52nv6);
assign Hu48v6 = (T8kiw6 ? Fpo7z6[3] : D62nv6);
assign Au48v6 = (T8kiw6 ? Fpo7z6[4] : K62nv6);
assign Tt48v6 = (T8kiw6 ? Fpo7z6[5] : R62nv6);
assign Mt48v6 = (T8kiw6 ? Fpo7z6[6] : U47iw6);
assign Ft48v6 = (T8kiw6 ? Fpo7z6[7] : J27iw6);
assign Ys48v6 = (T8kiw6 ? Fpo7z6[8] : H17iw6);
assign Rs48v6 = (T8kiw6 ? Fpo7z6[9] : Dz6iw6);
assign Ks48v6 = (T8kiw6 ? Fpo7z6[10] : Emhov6);
assign Ds48v6 = (T8kiw6 ? Fpo7z6[11] : Guhov6);
assign Wr48v6 = (T8kiw6 ? Fpo7z6[12] : Bk6iw6);
assign Pr48v6 = (T8kiw6 ? Fpo7z6[13] : Z0iov6);
assign Ir48v6 = (T8kiw6 ? Fpo7z6[14] : Is5iw6);
assign Br48v6 = (T8kiw6 ? Fpo7z6[15] : Gr5iw6);
assign Uq48v6 = (T8kiw6 ? Fpo7z6[16] : Jp5iw6);
assign Nq48v6 = (T8kiw6 ? Fpo7z6[17] : Mn5iw6);
assign Gq48v6 = (T8kiw6 ? Fpo7z6[18] : Bl5iw6);
assign Zp48v6 = (T8kiw6 ? Fpo7z6[19] : Ej5iw6);
assign Sp48v6 = (T8kiw6 ? Fpo7z6[20] : D85iw6);
assign Lp48v6 = (T8kiw6 ? Fpo7z6[21] : Cx4iw6);
assign T8kiw6 = (!A9kiw6);
assign Ep48v6 = (A9kiw6 ? Wf4iw6 : Fpo7z6[22]);
assign Xo48v6 = (A9kiw6 ? Iklov6 : Fpo7z6[23]);
assign Qo48v6 = (A9kiw6 ? E64iw6 : Fpo7z6[24]);
assign Jo48v6 = (A9kiw6 ? H44iw6 : Fpo7z6[25]);
assign Co48v6 = (A9kiw6 ? W14iw6 : Fpo7z6[26]);
assign Vn48v6 = (A9kiw6 ? I52nv6 : Fpo7z6[0]);
assign On48v6 = (A9kiw6 ? U42nv6 : Jj1ft6);
assign A9kiw6 = (J3kiw6 & H9kiw6);
assign J3kiw6 = (O9kiw6 & V9kiw6);
assign V9kiw6 = (M1kiw6 & Vd2iw6);
assign M1kiw6 = (Cakiw6 | Znn7z6[1]);
assign O9kiw6 = (D02ft6 & Jakiw6);
assign Jakiw6 = (~(Qakiw6 & Znn7z6[1]));
assign Hn48v6 = (~(Rconv6 & Xakiw6));
assign Xakiw6 = (~(Ebkiw6 & Lbkiw6));
assign Ebkiw6 = (Sbkiw6 & Kconv6);
assign Sbkiw6 = (~(Dconv6 & Wp9ov6));
assign An48v6 = (M4xnv6 ? Ryadt6 : Zbkiw6);
assign Zbkiw6 = (~(H2kiw6 | A2kiw6));
assign A2kiw6 = (~(Fr9ov6 | Gckiw6));
assign Fr9ov6 = (~(Nckiw6 & Uckiw6));
assign Uckiw6 = (Bdkiw6 & Idkiw6);
assign Idkiw6 = (~(Pdkiw6 & Pyo7z6[0]));
assign Bdkiw6 = (Wdkiw6 & Dekiw6);
assign Dekiw6 = (~(Kekiw6 & I1p7z6[0]));
assign Wdkiw6 = (~(Rekiw6 & Ws1ft6));
assign Nckiw6 = (Yekiw6 & Ffkiw6);
assign Ffkiw6 = (~(Mfkiw6 & Nw1ft6));
assign Yekiw6 = (Tfkiw6 & Agkiw6);
assign Agkiw6 = (~(Hgkiw6 & Wvo7z6[0]));
assign Tfkiw6 = (~(Ogkiw6 & Dto7z6[0]));
assign Tm48v6 = (Mr9ov6 ? Hrb7z6[1] : Gckiw6);
assign Gckiw6 = (~(Vgkiw6 & Chkiw6));
assign Chkiw6 = (Jhkiw6 & Qhkiw6);
assign Qhkiw6 = (~(Pdkiw6 & Pyo7z6[1]));
assign Jhkiw6 = (Xhkiw6 & Eikiw6);
assign Eikiw6 = (~(Kekiw6 & I1p7z6[1]));
assign Xhkiw6 = (~(Rekiw6 & Cu1ft6));
assign Vgkiw6 = (Likiw6 & Sikiw6);
assign Sikiw6 = (~(Mfkiw6 & Tx1ft6));
assign Likiw6 = (Zikiw6 & Gjkiw6);
assign Gjkiw6 = (~(Hgkiw6 & Wvo7z6[1]));
assign Zikiw6 = (~(Ogkiw6 & Dto7z6[1]));
assign Mm48v6 = (Rconv6 ? Njkiw6 : Kqm7z6[0]);
assign Fm48v6 = (Rconv6 ? Ujkiw6 : Kqm7z6[1]);
assign Ujkiw6 = (~(Bkkiw6 | Njkiw6));
assign Yl48v6 = (Rconv6 ? Bkkiw6 : Kqm7z6[2]);
assign Rl48v6 = (Pkkiw6 ? Geynv6 : Ikkiw6);
assign Ikkiw6 = (!Y877z6);
assign Kl48v6 = (Pkkiw6 ? Viynv6 : Wkkiw6);
assign Wkkiw6 = (!S777z6);
assign Dl48v6 = (Klkiw6 ? Viynv6 : Dlkiw6);
assign Dlkiw6 = (!I877z6);
assign Wk48v6 = (Pkkiw6 ? Knynv6 : Rlkiw6);
assign Rlkiw6 = (!M677z6);
assign Pk48v6 = (Klkiw6 ? Knynv6 : Ylkiw6);
assign Ylkiw6 = (!C777z6);
assign Ik48v6 = (Pkkiw6 ? Zrynv6 : Fmkiw6);
assign Fmkiw6 = (!G577z6);
assign Bk48v6 = (Klkiw6 ? Zrynv6 : Mmkiw6);
assign Mmkiw6 = (!W577z6);
assign Uj48v6 = (Pkkiw6 ? Owynv6 : Tmkiw6);
assign Tmkiw6 = (!A477z6);
assign Nj48v6 = (Klkiw6 ? Owynv6 : Ankiw6);
assign Ankiw6 = (!Q477z6);
assign Gj48v6 = (Pkkiw6 ? D1znv6 : Hnkiw6);
assign Hnkiw6 = (!U277z6);
assign Zi48v6 = (Klkiw6 ? D1znv6 : Onkiw6);
assign Onkiw6 = (!K377z6);
assign Si48v6 = (Pkkiw6 ? S5znv6 : Vnkiw6);
assign Vnkiw6 = (!O177z6);
assign Li48v6 = (Klkiw6 ? S5znv6 : Cokiw6);
assign Cokiw6 = (!E277z6);
assign Ei48v6 = (Pkkiw6 ? N1xnv6 : Jokiw6);
assign Jokiw6 = (!I077z6);
assign Xh48v6 = (Klkiw6 ? N1xnv6 : Qokiw6);
assign Qokiw6 = (!Y077z6);
assign Qh48v6 = (Pkkiw6 ? Eexnv6 : Xokiw6);
assign Xokiw6 = (!Cz67z6);
assign Jh48v6 = (Klkiw6 ? Eexnv6 : Epkiw6);
assign Epkiw6 = (!Sz67z6);
assign Ch48v6 = (Pkkiw6 ? Tixnv6 : Lpkiw6);
assign Lpkiw6 = (!Wx67z6);
assign Vg48v6 = (Klkiw6 ? Tixnv6 : Spkiw6);
assign Spkiw6 = (!My67z6);
assign Og48v6 = (!Zpkiw6);
assign Zpkiw6 = (Pkkiw6 ? Gqkiw6 : Qw67z6);
assign Hg48v6 = (!Nqkiw6);
assign Nqkiw6 = (Klkiw6 ? Gqkiw6 : Gx67z6);
assign Gqkiw6 = (!Inxnv6);
assign Ag48v6 = (!Uqkiw6);
assign Uqkiw6 = (Pkkiw6 ? Brkiw6 : Kv67z6);
assign Tf48v6 = (!Irkiw6);
assign Irkiw6 = (Klkiw6 ? Brkiw6 : Aw67z6);
assign Brkiw6 = (!Xrxnv6);
assign Mf48v6 = (!Prkiw6);
assign Prkiw6 = (Tqoov6 ? Eu67z6 : Wrkiw6);
assign Ff48v6 = (!Dskiw6);
assign Dskiw6 = (As9ov6 ? Uu67z6 : Wrkiw6);
assign Wrkiw6 = (!Mwxnv6);
assign Ye48v6 = (!Kskiw6);
assign Kskiw6 = (Tqoov6 ? Ys67z6 : Rskiw6);
assign Re48v6 = (!Yskiw6);
assign Yskiw6 = (As9ov6 ? Ot67z6 : Rskiw6);
assign Rskiw6 = (!B1ynv6);
assign Ke48v6 = (!Ftkiw6);
assign Ftkiw6 = (Pkkiw6 ? Mtkiw6 : O977z6);
assign De48v6 = (!Ttkiw6);
assign Ttkiw6 = (Klkiw6 ? Mtkiw6 : Ea77z6);
assign Mtkiw6 = (!Kaxnv6);
assign Wd48v6 = (Aukiw6 & Tlmov6);
assign Pd48v6 = (Hukiw6 & Oukiw6);
assign Oukiw6 = (O5a7z6 & Vukiw6);
assign Vukiw6 = (~(Cvkiw6 & Jvkiw6));
assign Jvkiw6 = (~(Qvkiw6 & Hmmov6));
assign Hmmov6 = (!Ihnet6);
assign Cvkiw6 = (Xvkiw6 & Mlmov6);
assign Hukiw6 = (~(Tr8iw6 | Whhov6));
assign Id48v6 = (Ewkiw6 & Tlmov6);
assign Bd48v6 = (Lwkiw6 & Ewkiw6);
assign Uc48v6 = (Swkiw6 & Ewkiw6);
assign Ewkiw6 = (Zwkiw6 & Ihnet6);
assign Zwkiw6 = (O5a7z6 & Gimov6);
assign Nc48v6 = (Lwkiw6 & Aukiw6);
assign Lwkiw6 = (Ow2et6 & Whhov6);
assign Gc48v6 = (Swkiw6 & Aukiw6);
assign Aukiw6 = (Gxkiw6 & Nxkiw6);
assign Nxkiw6 = (Xvkiw6 & Gimov6);
assign Gimov6 = (!Pl7et6);
assign Gxkiw6 = (A0onv6 & O5a7z6);
assign Swkiw6 = (Whhov6 & Uxkiw6);
assign Zb48v6 = (~(Fsfov6 & Bykiw6));
assign Bykiw6 = (~(Cmbdt6 & Iykiw6));
assign Iykiw6 = (F02nv6 | Z2onv6);
assign Z2onv6 = (Vs9ov6 & Kkmhw6);
assign Sb48v6 = (Pykiw6 & Wykiw6);
assign Wykiw6 = (Tlmov6 & O5a7z6);
assign Pykiw6 = (~(Xvkiw6 | Qvkiw6));
assign Xvkiw6 = (Flmov6 | Uxkiw6);
assign Uxkiw6 = (!Ow2et6);
assign Flmov6 = (~(Xnh7z6[2] & Dzkiw6));
assign Lb48v6 = (~(Kzkiw6 & Rzkiw6));
assign Rzkiw6 = (Yzkiw6 | Orhov6);
assign Kzkiw6 = (Hhq7z6[0] ? M0liw6 : F0liw6);
assign Eb48v6 = (~(T0liw6 & A1liw6));
assign A1liw6 = (Yzkiw6 | L19iw6);
assign T0liw6 = (Hhq7z6[1] ? O1liw6 : H1liw6);
assign H1liw6 = (~(V1liw6 & Hhq7z6[0]));
assign Xa48v6 = (~(C2liw6 & J2liw6));
assign J2liw6 = (Yzkiw6 | Fhrnv6);
assign C2liw6 = (Hhq7z6[2] ? X2liw6 : Q2liw6);
assign X2liw6 = (O1liw6 & E3liw6);
assign E3liw6 = (F0liw6 | Hhq7z6[1]);
assign O1liw6 = (M0liw6 & L3liw6);
assign L3liw6 = (F0liw6 | Hhq7z6[0]);
assign Q2liw6 = (~(S3liw6 & V1liw6));
assign Qa48v6 = (~(Z3liw6 & G4liw6));
assign G4liw6 = (Yzkiw6 | Pohov6);
assign Z3liw6 = (B5liw6 ? U4liw6 : N4liw6);
assign U4liw6 = (~(I5liw6 & V1liw6));
assign Ja48v6 = (~(P5liw6 & W5liw6));
assign W5liw6 = (Yzkiw6 | Zaeiw6);
assign P5liw6 = (Hhq7z6[4] ? K6liw6 : D6liw6);
assign K6liw6 = (N4liw6 & R6liw6);
assign R6liw6 = (~(V1liw6 & B5liw6));
assign B5liw6 = (!Hhq7z6[3]);
assign N4liw6 = (M0liw6 & Y6liw6);
assign Y6liw6 = (F0liw6 | I5liw6);
assign D6liw6 = (~(F7liw6 & I5liw6));
assign F7liw6 = (V1liw6 & Hhq7z6[3]);
assign Ca48v6 = (~(M7liw6 & T7liw6));
assign T7liw6 = (Yzkiw6 | Tdfiw6);
assign M7liw6 = (Hhq7z6[5] ? H8liw6 : A8liw6);
assign A8liw6 = (O8liw6 | F0liw6);
assign V948v6 = (~(V8liw6 & C9liw6));
assign C9liw6 = (Yzkiw6 | Gbeiw6);
assign V8liw6 = (Hhq7z6[6] ? Q9liw6 : J9liw6);
assign O948v6 = (~(X9liw6 & Ealiw6));
assign Ealiw6 = (Yzkiw6 | Egfiw6);
assign X9liw6 = (Hhq7z6[7] ? Saliw6 : Laliw6);
assign Saliw6 = (Q9liw6 & Zaliw6);
assign Zaliw6 = (~(V1liw6 & Gbliw6));
assign Q9liw6 = (H8liw6 & Nbliw6);
assign Nbliw6 = (F0liw6 | Hhq7z6[5]);
assign H8liw6 = (M0liw6 & Ubliw6);
assign Ubliw6 = (~(V1liw6 & O8liw6));
assign Laliw6 = (J9liw6 | Gbliw6);
assign Gbliw6 = (!Hhq7z6[6]);
assign J9liw6 = (Bcliw6 | O8liw6);
assign Bcliw6 = (~(V1liw6 & Hhq7z6[5]));
assign V1liw6 = (!F0liw6);
assign F0liw6 = (~(Icliw6 & Pcliw6));
assign Icliw6 = (M0liw6 & Yzkiw6);
assign M0liw6 = (~(Wcliw6 & Pcliw6));
assign Pcliw6 = (~(Ddliw6 & Etgiw6));
assign Ddliw6 = (Kdliw6 & Jp5iw6);
assign Kdliw6 = (~(Xkq7z6[18] & HTMDHBURST[0]));
assign Wcliw6 = (Yzkiw6 & Rdliw6);
assign Yzkiw6 = (~(Jsgiw6 & Ydliw6));
assign H948v6 = (Teliw6 ? Meliw6 : Feliw6);
assign Meliw6 = (Dtadt6 & Tnzdt6);
assign Feliw6 = (Afliw6 & Ku7et6);
assign Afliw6 = (U28et6 & Lo1ov6);
assign A948v6 = (Lo1ov6 & Hfliw6);
assign Lo1ov6 = (Tlmov6 | Kslov6);
assign T848v6 = (Ofliw6 & Vfliw6);
assign Vfliw6 = (~(Cgliw6 | Zofov6));
assign Zofov6 = (Yfadt6 & Qg2nv6);
assign Cgliw6 = (~(Sh2nv6 & Jgliw6));
assign Ofliw6 = (Kslov6 & Kihov6);
assign M848v6 = (Qgliw6 & Jgliw6);
assign Qgliw6 = (~(Kslov6 & Kihov6));
assign F848v6 = (Xgliw6 & Jgliw6);
assign Xgliw6 = (~(Vsgov6 & Sh2nv6));
assign Y748v6 = (Lhliw6 ? Tjr7z6[1] : Ehliw6);
assign R748v6 = (Lhliw6 ? Tjr7z6[0] : W3wnv6);
assign K748v6 = (~(Shliw6 & Zhliw6));
assign Zhliw6 = (Qxjov6 | Giliw6);
assign Shliw6 = (Niliw6 & Uiliw6);
assign Uiliw6 = (~(Bjliw6 & P2j7z6[1]));
assign Niliw6 = (~(Qmb7z6[1] & Jxjov6));
assign D748v6 = (~(Ijliw6 & Pjliw6));
assign Pjliw6 = (Qxjov6 | Wjliw6);
assign Ijliw6 = (Dkliw6 & Kkliw6);
assign Kkliw6 = (~(Bjliw6 & P2j7z6[2]));
assign Dkliw6 = (~(Qmb7z6[2] & Jxjov6));
assign W648v6 = (~(Rkliw6 & Ykliw6));
assign Ykliw6 = (Qxjov6 | Flliw6);
assign Rkliw6 = (Mlliw6 & Tlliw6);
assign Tlliw6 = (~(Bjliw6 & P2j7z6[3]));
assign Mlliw6 = (~(Qmb7z6[3] & Jxjov6));
assign P648v6 = (~(Amliw6 & Hmliw6));
assign Hmliw6 = (Qxjov6 | Omliw6);
assign Amliw6 = (Vmliw6 & Cnliw6);
assign Cnliw6 = (~(Bjliw6 & P2j7z6[4]));
assign Vmliw6 = (~(Qmb7z6[4] & Jxjov6));
assign I648v6 = (~(Jnliw6 & Qnliw6));
assign Qnliw6 = (Qxjov6 | Xnliw6);
assign Jnliw6 = (Eoliw6 & Loliw6);
assign Loliw6 = (~(Bjliw6 & P2j7z6[5]));
assign Eoliw6 = (~(Qmb7z6[5] & Jxjov6));
assign B648v6 = (~(Soliw6 & Zoliw6));
assign Zoliw6 = (Qxjov6 | Gpliw6);
assign Soliw6 = (Npliw6 & Upliw6);
assign Upliw6 = (~(Bjliw6 & P2j7z6[6]));
assign Npliw6 = (~(Qmb7z6[6] & Jxjov6));
assign U548v6 = (~(Bqliw6 & Iqliw6));
assign Iqliw6 = (~(Qmb7z6[7] & Jxjov6));
assign Bqliw6 = (Qxjov6 | Pqliw6);
assign N548v6 = (~(Wqliw6 & Drliw6));
assign Drliw6 = (Qxjov6 | Krliw6);
assign Wqliw6 = (Rrliw6 & Yrliw6);
assign Yrliw6 = (~(Bjliw6 & P2j7z6[0]));
assign Bjliw6 = (~(Ga3nv6 | Fsliw6));
assign Rrliw6 = (~(Qmb7z6[0] & Jxjov6));
assign Jxjov6 = (Msliw6 & Qxjov6);
assign Qxjov6 = (~(Tsliw6 & Kslov6));
assign Tsliw6 = (~(Fsliw6 | Lcadt6));
assign Msliw6 = (U4fov6 & Ga3nv6);
assign G548v6 = (~(Atliw6 & Htliw6));
assign Htliw6 = (~(G5j7z6[0] & Otliw6));
assign Otliw6 = (~(Vtliw6 & Culiw6));
assign Z448v6 = (!Juliw6);
assign Juliw6 = (M6j7z6[0] ? Xuliw6 : Quliw6);
assign Xuliw6 = (~(Evliw6 & Atliw6));
assign Atliw6 = (~(Lvliw6 & Svliw6));
assign Lvliw6 = (~(Zvliw6 | G5j7z6[0]));
assign Evliw6 = (~(Gwliw6 & U42nv6));
assign Quliw6 = (Nwliw6 & Uwliw6);
assign Uwliw6 = (~(Bxliw6 & U42nv6));
assign Nwliw6 = (~(Qkj7z6[0] | Ixliw6));
assign Ixliw6 = (Pxliw6 & Tib7z6[0]);
assign Pxliw6 = (~(Jqj7z6[9] & G5j7z6[0]));
assign S448v6 = (~(Wxliw6 & Dyliw6));
assign Dyliw6 = (~(G5j7z6[2] & Kyliw6));
assign Kyliw6 = (~(Vtliw6 & Ryliw6));
assign L448v6 = (!Yyliw6);
assign Yyliw6 = (M6j7z6[2] ? Mzliw6 : Fzliw6);
assign Mzliw6 = (~(Wxliw6 & Tzliw6));
assign Tzliw6 = (~(Gwliw6 & I52nv6));
assign Wxliw6 = (~(A0miw6 & H0miw6));
assign A0miw6 = (~(Rxgov6 | G5j7z6[2]));
assign Fzliw6 = (O0miw6 & V0miw6);
assign V0miw6 = (~(Bxliw6 & I52nv6));
assign O0miw6 = (~(Qkj7z6[2] | C1miw6));
assign C1miw6 = (J1miw6 & Tib7z6[2]);
assign J1miw6 = (~(Jqj7z6[11] & G5j7z6[2]));
assign E448v6 = (~(Q1miw6 & X1miw6));
assign X1miw6 = (~(G5j7z6[4] & E2miw6));
assign E2miw6 = (~(Vtliw6 & L2miw6));
assign X348v6 = (!S2miw6);
assign S2miw6 = (M6j7z6[4] ? G3miw6 : Z2miw6);
assign G3miw6 = (~(N3miw6 & Q1miw6));
assign Q1miw6 = (~(U3miw6 & H0miw6));
assign U3miw6 = (Uuhov6 & B4miw6);
assign N3miw6 = (~(Gwliw6 & W52nv6));
assign Z2miw6 = (I4miw6 & P4miw6);
assign P4miw6 = (~(Bxliw6 & W52nv6));
assign I4miw6 = (~(Qkj7z6[4] | W4miw6));
assign W4miw6 = (D5miw6 & Tib7z6[4]);
assign D5miw6 = (~(Jqj7z6[13] & G5j7z6[4]));
assign Q348v6 = (~(K5miw6 & R5miw6));
assign R5miw6 = (~(G5j7z6[6] & Y5miw6));
assign Y5miw6 = (~(Vtliw6 & F6miw6));
assign J348v6 = (!M6miw6);
assign M6miw6 = (M6j7z6[6] ? A7miw6 : T6miw6);
assign A7miw6 = (~(K5miw6 & H7miw6));
assign H7miw6 = (~(Gwliw6 & K62nv6));
assign K5miw6 = (~(O7miw6 & H0miw6));
assign O7miw6 = (Gnhov6 & V7miw6);
assign T6miw6 = (C8miw6 & J8miw6);
assign J8miw6 = (~(Bxliw6 & K62nv6));
assign C8miw6 = (~(Qkj7z6[6] | Q8miw6));
assign Q8miw6 = (X8miw6 & Tib7z6[6]);
assign X8miw6 = (~(Jqj7z6[15] & G5j7z6[6]));
assign C348v6 = (~(E9miw6 & L9miw6));
assign L9miw6 = (~(G5j7z6[16] & S9miw6));
assign E9miw6 = (Z9miw6 & Gamiw6);
assign Z9miw6 = (Namiw6 | Fsliw6);
assign V248v6 = (!Uamiw6);
assign Uamiw6 = (M6j7z6[16] ? Ibmiw6 : Bbmiw6);
assign Ibmiw6 = (~(Pbmiw6 & Gamiw6));
assign Gamiw6 = (~(Wbmiw6 & Svliw6));
assign Wbmiw6 = (Dcmiw6 & Cu2nv6);
assign Cu2nv6 = (!G5j7z6[16]);
assign Pbmiw6 = (~(Kcmiw6 & Is5iw6));
assign Bbmiw6 = (Rcmiw6 & Ycmiw6);
assign Ycmiw6 = (~(Fdmiw6 & Is5iw6));
assign Rcmiw6 = (~(Qkj7z6[16] | Mdmiw6));
assign Mdmiw6 = (Tdmiw6 & Tib7z6[16]);
assign Tdmiw6 = (~(Jqj7z6[25] & G5j7z6[16]));
assign O248v6 = (~(Aemiw6 & Hemiw6));
assign Hemiw6 = (~(Oemiw6 & G5j7z6[18]));
assign Oemiw6 = (Vemiw6 & U4fov6);
assign Vemiw6 = (~(Cfmiw6 & Jfmiw6));
assign H248v6 = (!Qfmiw6);
assign Qfmiw6 = (M6j7z6[18] ? Egmiw6 : Xfmiw6);
assign Egmiw6 = (~(Aemiw6 & Lgmiw6));
assign Lgmiw6 = (~(Kcmiw6 & Jp5iw6));
assign Aemiw6 = (~(Sgmiw6 & Dcmiw6));
assign Sgmiw6 = (~(Rxgov6 | G5j7z6[18]));
assign Xfmiw6 = (Zgmiw6 & Ghmiw6);
assign Ghmiw6 = (~(Fdmiw6 & Jp5iw6));
assign Zgmiw6 = (~(Qkj7z6[18] | Nhmiw6));
assign Nhmiw6 = (Uhmiw6 & Tib7z6[18]);
assign Uhmiw6 = (~(Jqj7z6[27] & G5j7z6[18]));
assign A248v6 = (~(Bimiw6 & Iimiw6));
assign Iimiw6 = (~(G5j7z6[20] & Pimiw6));
assign Pimiw6 = (~(Wimiw6 & L2miw6));
assign T148v6 = (!Djmiw6);
assign Djmiw6 = (M6j7z6[20] ? Rjmiw6 : Kjmiw6);
assign Rjmiw6 = (~(Yjmiw6 & Bimiw6));
assign Bimiw6 = (~(Fkmiw6 & Dcmiw6));
assign Fkmiw6 = (Uuhov6 & Mkmiw6);
assign Yjmiw6 = (~(Kcmiw6 & Bl5iw6));
assign Kjmiw6 = (Tkmiw6 & Almiw6);
assign Almiw6 = (~(Fdmiw6 & Bl5iw6));
assign Tkmiw6 = (~(Qkj7z6[20] | Hlmiw6));
assign Hlmiw6 = (Olmiw6 & Tib7z6[20]);
assign Olmiw6 = (~(Jqj7z6[29] & G5j7z6[20]));
assign M148v6 = (~(Vlmiw6 & Cmmiw6));
assign Cmmiw6 = (~(Jmmiw6 & G5j7z6[22]));
assign Jmmiw6 = (Qmmiw6 & U4fov6);
assign Qmmiw6 = (~(Cfmiw6 & Rphov6));
assign F148v6 = (!Xmmiw6);
assign Xmmiw6 = (M6j7z6[22] ? Lnmiw6 : Enmiw6);
assign Lnmiw6 = (~(Vlmiw6 & Snmiw6));
assign Snmiw6 = (~(Kcmiw6 & D85iw6));
assign Vlmiw6 = (~(Znmiw6 & Dcmiw6));
assign Znmiw6 = (Gnhov6 & Gomiw6);
assign Enmiw6 = (Nomiw6 & Uomiw6);
assign Uomiw6 = (~(Fdmiw6 & D85iw6));
assign Nomiw6 = (~(Qkj7z6[22] | Bpmiw6));
assign Bpmiw6 = (Ipmiw6 & Tib7z6[22]);
assign Ipmiw6 = (~(Jqj7z6[31] & G5j7z6[22]));
assign Y048v6 = (~(Ppmiw6 & Wpmiw6));
assign Wpmiw6 = (~(G5j7z6[32] & Dqmiw6));
assign Dqmiw6 = (~(Kqmiw6 & Culiw6));
assign Culiw6 = (~(Rqmiw6 & U4fov6));
assign R048v6 = (!Yqmiw6);
assign Yqmiw6 = (M6j7z6[32] ? Mrmiw6 : Frmiw6);
assign Mrmiw6 = (~(Trmiw6 & Ppmiw6));
assign Ppmiw6 = (~(Asmiw6 & Svliw6));
assign Asmiw6 = (A5iov6 & Hsmiw6);
assign Trmiw6 = (~(Osmiw6 & U42nv6));
assign Frmiw6 = (Vsmiw6 & Ctmiw6);
assign Ctmiw6 = (~(Jtmiw6 & U42nv6));
assign Vsmiw6 = (~(Qkj7z6[32] | Qtmiw6));
assign Qtmiw6 = (Xtmiw6 & Tib7z6[32]);
assign Xtmiw6 = (~(Jqj7z6[41] & G5j7z6[32]));
assign K048v6 = (~(Eumiw6 & Lumiw6));
assign Lumiw6 = (~(G5j7z6[34] & Sumiw6));
assign Sumiw6 = (~(D3iov6 & Ryliw6));
assign Ryliw6 = (~(U4fov6 & Zumiw6));
assign D048v6 = (!Gvmiw6);
assign Gvmiw6 = (M6j7z6[34] ? Uvmiw6 : Nvmiw6);
assign Uvmiw6 = (~(Eumiw6 & Bwmiw6));
assign Bwmiw6 = (~(Osmiw6 & I52nv6));
assign Eumiw6 = (~(Iwmiw6 & A5iov6));
assign Iwmiw6 = (~(Rxgov6 | G5j7z6[34]));
assign Nvmiw6 = (Pwmiw6 & Wwmiw6);
assign Wwmiw6 = (~(Jtmiw6 & I52nv6));
assign Pwmiw6 = (~(Qkj7z6[34] | Dxmiw6));
assign Dxmiw6 = (Kxmiw6 & Tib7z6[34]);
assign Kxmiw6 = (~(Jqj7z6[43] & G5j7z6[34]));
assign Wz38v6 = (~(Rxmiw6 & Yxmiw6));
assign Yxmiw6 = (~(G5j7z6[36] & Fymiw6));
assign Fymiw6 = (~(Kqmiw6 & L2miw6));
assign Pz38v6 = (!Mymiw6);
assign Mymiw6 = (M6j7z6[36] ? Azmiw6 : Tymiw6);
assign Azmiw6 = (~(Hzmiw6 & Rxmiw6));
assign Rxmiw6 = (~(Ozmiw6 & A5iov6));
assign Ozmiw6 = (Uuhov6 & Vzmiw6);
assign Hzmiw6 = (~(Osmiw6 & W52nv6));
assign Tymiw6 = (C0niw6 & J0niw6);
assign J0niw6 = (~(Jtmiw6 & W52nv6));
assign C0niw6 = (~(Qkj7z6[36] | Q0niw6));
assign Q0niw6 = (X0niw6 & Tib7z6[36]);
assign X0niw6 = (~(Jqj7z6[45] & G5j7z6[36]));
assign Iz38v6 = (~(E1niw6 & L1niw6));
assign L1niw6 = (~(G5j7z6[38] & S1niw6));
assign S1niw6 = (~(D3iov6 & F6miw6));
assign Bz38v6 = (!Z1niw6);
assign Z1niw6 = (M6j7z6[38] ? N2niw6 : G2niw6);
assign N2niw6 = (~(E1niw6 & U2niw6));
assign U2niw6 = (~(Osmiw6 & K62nv6));
assign E1niw6 = (~(B3niw6 & A5iov6));
assign B3niw6 = (Gnhov6 & I3niw6);
assign G2niw6 = (P3niw6 & W3niw6);
assign W3niw6 = (~(Jtmiw6 & K62nv6));
assign P3niw6 = (~(Qkj7z6[38] | D4niw6));
assign D4niw6 = (K4niw6 & Tib7z6[38]);
assign K4niw6 = (~(Jqj7z6[47] & G5j7z6[38]));
assign Uy38v6 = (~(R4niw6 & Y4niw6));
assign Y4niw6 = (~(F5niw6 & U4fov6));
assign R4niw6 = (M5niw6 & T5niw6);
assign M5niw6 = (Z3fov6 | A6niw6);
assign Ny38v6 = (!H6niw6);
assign H6niw6 = (M6j7z6[48] ? V6niw6 : O6niw6);
assign V6niw6 = (~(C7niw6 & T5niw6));
assign T5niw6 = (~(J7niw6 & Svliw6));
assign Svliw6 = (Q7niw6 & Rgjov6);
assign J7niw6 = (R4hov6 & A6niw6);
assign A6niw6 = (!G5j7z6[48]);
assign C7niw6 = (~(X7niw6 & Is5iw6));
assign O6niw6 = (E8niw6 & L8niw6);
assign L8niw6 = (~(S8niw6 & Is5iw6));
assign E8niw6 = (~(Qkj7z6[48] | Z8niw6));
assign Z8niw6 = (G9niw6 & Tib7z6[48]);
assign G9niw6 = (~(Jqj7z6[57] & G5j7z6[48]));
assign Gy38v6 = (~(N9niw6 & U9niw6));
assign U9niw6 = (~(Baniw6 & U4fov6));
assign N9niw6 = (Ianiw6 & Paniw6);
assign Ianiw6 = (Z3fov6 | Fs2nv6);
assign Fs2nv6 = (!G5j7z6[50]);
assign Zx38v6 = (!Waniw6);
assign Waniw6 = (M6j7z6[50] ? Kbniw6 : Dbniw6);
assign Kbniw6 = (~(Rbniw6 & Paniw6));
assign Paniw6 = (~(Ybniw6 & R4hov6));
assign Ybniw6 = (~(Rxgov6 | G5j7z6[50]));
assign Rbniw6 = (~(X7niw6 & Jp5iw6));
assign Dbniw6 = (Fcniw6 & Mcniw6);
assign Mcniw6 = (~(S8niw6 & Jp5iw6));
assign Fcniw6 = (~(Qkj7z6[50] | Tcniw6));
assign Tcniw6 = (Adniw6 & Tib7z6[50]);
assign Adniw6 = (~(Jqj7z6[59] & G5j7z6[50]));
assign Sx38v6 = (~(Hdniw6 & Odniw6));
assign Odniw6 = (~(G5j7z6[1] & Vdniw6));
assign Vdniw6 = (~(Vtliw6 & Ceniw6));
assign Lx38v6 = (!Jeniw6);
assign Jeniw6 = (M6j7z6[1] ? Xeniw6 : Qeniw6);
assign Xeniw6 = (~(Hdniw6 & Efniw6));
assign Efniw6 = (~(Gwliw6 & B52nv6));
assign Hdniw6 = (~(Lfniw6 & Sfniw6));
assign Lfniw6 = (~(Zvliw6 | G5j7z6[1]));
assign Qeniw6 = (Zfniw6 & Ggniw6);
assign Ggniw6 = (~(Bxliw6 & B52nv6));
assign Zfniw6 = (~(Qkj7z6[1] | Ngniw6));
assign Ngniw6 = (Ugniw6 & Tib7z6[1]);
assign Ugniw6 = (~(Jqj7z6[10] & G5j7z6[1]));
assign Ex38v6 = (~(Bhniw6 & Ihniw6));
assign Ihniw6 = (~(G5j7z6[3] & Phniw6));
assign Phniw6 = (~(Vtliw6 & Whniw6));
assign Xw38v6 = (!Diniw6);
assign Diniw6 = (M6j7z6[3] ? Riniw6 : Kiniw6);
assign Riniw6 = (~(Bhniw6 & Yiniw6));
assign Yiniw6 = (~(Gwliw6 & P52nv6));
assign Bhniw6 = (~(Fjniw6 & Mjniw6));
assign Fjniw6 = (~(Zvliw6 | G5j7z6[3]));
assign Zvliw6 = (!H0miw6);
assign Kiniw6 = (Tjniw6 & Akniw6);
assign Akniw6 = (~(Bxliw6 & P52nv6));
assign Tjniw6 = (~(Qkj7z6[3] | Hkniw6));
assign Hkniw6 = (Okniw6 & Tib7z6[3]);
assign Okniw6 = (~(Jqj7z6[12] & G5j7z6[3]));
assign Qw38v6 = (~(Vkniw6 & Clniw6));
assign Clniw6 = (~(G5j7z6[5] & Jlniw6));
assign Jlniw6 = (~(Vtliw6 & Qlniw6));
assign Jw38v6 = (!Xlniw6);
assign Xlniw6 = (M6j7z6[5] ? Lmniw6 : Emniw6);
assign Lmniw6 = (~(Vkniw6 & Smniw6));
assign Smniw6 = (~(Gwliw6 & D62nv6));
assign Vkniw6 = (~(Zmniw6 & H0miw6));
assign Zmniw6 = (Gnniw6 & Nnniw6);
assign Emniw6 = (Unniw6 & Boniw6);
assign Boniw6 = (~(Bxliw6 & D62nv6));
assign Unniw6 = (~(Qkj7z6[5] | Ioniw6));
assign Ioniw6 = (Poniw6 & Tib7z6[5]);
assign Poniw6 = (~(Jqj7z6[14] & G5j7z6[5]));
assign Cw38v6 = (~(Woniw6 & Dpniw6));
assign Dpniw6 = (~(G5j7z6[7] & Kpniw6));
assign Kpniw6 = (~(Vtliw6 & Rpniw6));
assign Vv38v6 = (!Ypniw6);
assign Ypniw6 = (M6j7z6[7] ? Mqniw6 : Fqniw6);
assign Mqniw6 = (~(Woniw6 & Tqniw6));
assign Tqniw6 = (~(Gwliw6 & R62nv6));
assign Gwliw6 = (~(Arniw6 | Twaiw6));
assign Woniw6 = (~(Hrniw6 & H0miw6));
assign Hrniw6 = (Orniw6 & Vrniw6);
assign Fqniw6 = (Csniw6 & Jsniw6);
assign Jsniw6 = (~(Bxliw6 & R62nv6));
assign Bxliw6 = (~(Qsniw6 | Twaiw6));
assign Csniw6 = (~(Qkj7z6[7] | Xsniw6));
assign Xsniw6 = (Etniw6 & Tib7z6[7]);
assign Etniw6 = (~(Jqj7z6[16] & G5j7z6[7]));
assign Ov38v6 = (~(Ltniw6 & Stniw6));
assign Stniw6 = (~(Ztniw6 & G5j7z6[17]));
assign Ztniw6 = (Guniw6 & U4fov6);
assign Guniw6 = (~(Cfmiw6 & Nuniw6));
assign Hv38v6 = (!Uuniw6);
assign Uuniw6 = (M6j7z6[17] ? Ivniw6 : Bvniw6);
assign Ivniw6 = (~(Ltniw6 & Pvniw6));
assign Pvniw6 = (~(Kcmiw6 & Gr5iw6));
assign Ltniw6 = (~(Wvniw6 & Sfniw6));
assign Wvniw6 = (Dcmiw6 & Ju2nv6);
assign Ju2nv6 = (!G5j7z6[17]);
assign Bvniw6 = (Dwniw6 & Kwniw6);
assign Kwniw6 = (~(Fdmiw6 & Gr5iw6));
assign Dwniw6 = (~(Qkj7z6[17] | Rwniw6));
assign Rwniw6 = (Ywniw6 & Tib7z6[17]);
assign Ywniw6 = (~(Jqj7z6[26] & G5j7z6[17]));
assign Av38v6 = (~(Fxniw6 & Mxniw6));
assign Mxniw6 = (~(Txniw6 & U4fov6));
assign Fxniw6 = (Ayniw6 & Hyniw6);
assign Ayniw6 = (Z3fov6 | Oyniw6);
assign Tu38v6 = (!Vyniw6);
assign Vyniw6 = (M6j7z6[19] ? Jzniw6 : Czniw6);
assign Jzniw6 = (~(Qzniw6 & Hyniw6));
assign Hyniw6 = (~(Xzniw6 & Mjniw6));
assign Xzniw6 = (Dcmiw6 & Oyniw6);
assign Oyniw6 = (!G5j7z6[19]);
assign Qzniw6 = (~(Kcmiw6 & Mn5iw6));
assign Czniw6 = (E0oiw6 & L0oiw6);
assign L0oiw6 = (~(Fdmiw6 & Mn5iw6));
assign E0oiw6 = (~(Qkj7z6[19] | S0oiw6));
assign S0oiw6 = (Z0oiw6 & Tib7z6[19]);
assign Z0oiw6 = (~(Jqj7z6[28] & G5j7z6[19]));
assign Mu38v6 = (~(G1oiw6 & N1oiw6));
assign N1oiw6 = (~(U1oiw6 & G5j7z6[21]));
assign U1oiw6 = (B2oiw6 & U4fov6);
assign B2oiw6 = (~(Cfmiw6 & I2oiw6));
assign Fu38v6 = (!P2oiw6);
assign P2oiw6 = (M6j7z6[21] ? D3oiw6 : W2oiw6);
assign D3oiw6 = (~(G1oiw6 & K3oiw6));
assign K3oiw6 = (~(Kcmiw6 & Ej5iw6));
assign G1oiw6 = (~(R3oiw6 & Dcmiw6));
assign R3oiw6 = (Gnniw6 & Y3oiw6);
assign W2oiw6 = (F4oiw6 & M4oiw6);
assign M4oiw6 = (~(Fdmiw6 & Ej5iw6));
assign F4oiw6 = (~(Qkj7z6[21] | T4oiw6));
assign T4oiw6 = (A5oiw6 & Tib7z6[21]);
assign A5oiw6 = (~(Jqj7z6[30] & G5j7z6[21]));
assign Yt38v6 = (~(H5oiw6 & O5oiw6));
assign O5oiw6 = (~(V5oiw6 & G5j7z6[23]));
assign V5oiw6 = (C6oiw6 & U4fov6);
assign C6oiw6 = (~(Cfmiw6 & J6oiw6));
assign Rt38v6 = (!Q6oiw6);
assign Q6oiw6 = (M6j7z6[23] ? E7oiw6 : X6oiw6);
assign E7oiw6 = (~(H5oiw6 & L7oiw6));
assign L7oiw6 = (~(Kcmiw6 & Cx4iw6));
assign Kcmiw6 = (~(Arniw6 | Ie5iw6));
assign H5oiw6 = (~(S7oiw6 & Dcmiw6));
assign S7oiw6 = (Orniw6 & Z7oiw6);
assign X6oiw6 = (G8oiw6 & N8oiw6);
assign N8oiw6 = (~(Fdmiw6 & Cx4iw6));
assign Fdmiw6 = (~(Qsniw6 | Ie5iw6));
assign G8oiw6 = (~(Qkj7z6[23] | U8oiw6));
assign U8oiw6 = (B9oiw6 & Tib7z6[23]);
assign B9oiw6 = (~(Jqj7z6[32] & G5j7z6[23]));
assign Kt38v6 = (~(I9oiw6 & P9oiw6));
assign P9oiw6 = (~(G5j7z6[33] & W9oiw6));
assign W9oiw6 = (~(D3iov6 & Ceniw6));
assign Ceniw6 = (~(U4fov6 & Daoiw6));
assign Dt38v6 = (!Kaoiw6);
assign Kaoiw6 = (M6j7z6[33] ? Yaoiw6 : Raoiw6);
assign Yaoiw6 = (~(I9oiw6 & Fboiw6));
assign Fboiw6 = (~(Osmiw6 & B52nv6));
assign I9oiw6 = (~(Mboiw6 & Sfniw6));
assign Mboiw6 = (A5iov6 & Tboiw6);
assign Raoiw6 = (Acoiw6 & Hcoiw6);
assign Hcoiw6 = (~(Jtmiw6 & B52nv6));
assign Acoiw6 = (~(Qkj7z6[33] | Ocoiw6));
assign Ocoiw6 = (Vcoiw6 & Tib7z6[33]);
assign Vcoiw6 = (~(Jqj7z6[42] & G5j7z6[33]));
assign Ws38v6 = (~(Cdoiw6 & Jdoiw6));
assign Jdoiw6 = (~(G5j7z6[35] & Qdoiw6));
assign Qdoiw6 = (~(D3iov6 & Whniw6));
assign Whniw6 = (~(Xdoiw6 & U4fov6));
assign Ps38v6 = (!Eeoiw6);
assign Eeoiw6 = (M6j7z6[35] ? Seoiw6 : Leoiw6);
assign Seoiw6 = (~(Cdoiw6 & Zeoiw6));
assign Zeoiw6 = (~(Osmiw6 & P52nv6));
assign Cdoiw6 = (~(Gfoiw6 & Mjniw6));
assign Gfoiw6 = (A5iov6 & Nfoiw6);
assign Leoiw6 = (Ufoiw6 & Bgoiw6);
assign Bgoiw6 = (~(Jtmiw6 & P52nv6));
assign Ufoiw6 = (~(Qkj7z6[35] | Igoiw6));
assign Igoiw6 = (Pgoiw6 & Tib7z6[35]);
assign Pgoiw6 = (~(Jqj7z6[44] & G5j7z6[35]));
assign Is38v6 = (~(Wgoiw6 & Dhoiw6));
assign Dhoiw6 = (~(G5j7z6[37] & Khoiw6));
assign Khoiw6 = (~(D3iov6 & Qlniw6));
assign Bs38v6 = (!Rhoiw6);
assign Rhoiw6 = (M6j7z6[37] ? Fioiw6 : Yhoiw6);
assign Fioiw6 = (~(Wgoiw6 & Mioiw6));
assign Mioiw6 = (~(Osmiw6 & D62nv6));
assign Wgoiw6 = (~(Tioiw6 & A5iov6));
assign Tioiw6 = (Gnniw6 & Ajoiw6);
assign Yhoiw6 = (Hjoiw6 & Ojoiw6);
assign Ojoiw6 = (~(Jtmiw6 & D62nv6));
assign Hjoiw6 = (~(Qkj7z6[37] | Vjoiw6));
assign Vjoiw6 = (Ckoiw6 & Tib7z6[37]);
assign Ckoiw6 = (~(Jqj7z6[46] & G5j7z6[37]));
assign Ur38v6 = (~(Jkoiw6 & Qkoiw6));
assign Qkoiw6 = (~(G5j7z6[39] & Xkoiw6));
assign Xkoiw6 = (~(D3iov6 & Rpniw6));
assign Nr38v6 = (!Eloiw6);
assign Eloiw6 = (M6j7z6[39] ? Sloiw6 : Lloiw6);
assign Sloiw6 = (~(Jkoiw6 & Zloiw6));
assign Zloiw6 = (~(Osmiw6 & R62nv6));
assign Osmiw6 = (Gmoiw6 & Bqi7z6[0]);
assign Gmoiw6 = (!Nmoiw6);
assign Jkoiw6 = (~(Umoiw6 & A5iov6));
assign Umoiw6 = (Orniw6 & Bnoiw6);
assign Lloiw6 = (Inoiw6 & Pnoiw6);
assign Pnoiw6 = (~(Jtmiw6 & R62nv6));
assign Jtmiw6 = (Wnoiw6 & Bqi7z6[0]);
assign Wnoiw6 = (!Dooiw6);
assign Inoiw6 = (~(Qkj7z6[39] | Kooiw6));
assign Kooiw6 = (Rooiw6 & Tib7z6[39]);
assign Rooiw6 = (~(Jqj7z6[48] & G5j7z6[39]));
assign Gr38v6 = (~(Yooiw6 & Fpoiw6));
assign Fpoiw6 = (Mpoiw6 | Fsliw6);
assign Yooiw6 = (Tpoiw6 & Aqoiw6);
assign Tpoiw6 = (Z3fov6 | Yr2nv6);
assign Zq38v6 = (!Hqoiw6);
assign Hqoiw6 = (M6j7z6[49] ? Vqoiw6 : Oqoiw6);
assign Vqoiw6 = (~(Croiw6 & Aqoiw6));
assign Aqoiw6 = (~(Jroiw6 & Sfniw6));
assign Sfniw6 = (~(Qroiw6 | P2j7z6[1]));
assign Jroiw6 = (R4hov6 & Yr2nv6);
assign Yr2nv6 = (!G5j7z6[49]);
assign Croiw6 = (~(X7niw6 & Gr5iw6));
assign Oqoiw6 = (Xroiw6 & Esoiw6);
assign Esoiw6 = (~(S8niw6 & Gr5iw6));
assign Xroiw6 = (~(Qkj7z6[49] | Lsoiw6));
assign Lsoiw6 = (Ssoiw6 & Tib7z6[49]);
assign Ssoiw6 = (~(Jqj7z6[58] & G5j7z6[49]));
assign Sq38v6 = (~(Zsoiw6 & Gtoiw6));
assign Gtoiw6 = (~(Ntoiw6 & U4fov6));
assign Zsoiw6 = (Utoiw6 & Buoiw6);
assign Utoiw6 = (Z3fov6 | Ms2nv6);
assign Lq38v6 = (!Iuoiw6);
assign Iuoiw6 = (M6j7z6[51] ? Wuoiw6 : Puoiw6);
assign Wuoiw6 = (~(Dvoiw6 & Buoiw6));
assign Buoiw6 = (~(Kvoiw6 & Mjniw6));
assign Kvoiw6 = (R4hov6 & Ms2nv6);
assign Ms2nv6 = (!G5j7z6[51]);
assign Dvoiw6 = (~(X7niw6 & Mn5iw6));
assign Puoiw6 = (Rvoiw6 & Yvoiw6);
assign Yvoiw6 = (~(S8niw6 & Mn5iw6));
assign Rvoiw6 = (~(Qkj7z6[51] | Fwoiw6));
assign Fwoiw6 = (Mwoiw6 & Tib7z6[51]);
assign Mwoiw6 = (~(Jqj7z6[60] & G5j7z6[51]));
assign Eq38v6 = (~(Twoiw6 & Axoiw6));
assign Axoiw6 = (~(Hxoiw6 & Oxoiw6));
assign Oxoiw6 = (~(A6oov6 | IFLUSH));
assign A6oov6 = (N8xnv6 & Znnov6);
assign Hxoiw6 = (D61ov6 & A3ddt6);
assign Twoiw6 = (~(Vxoiw6 & Cyoiw6));
assign Cyoiw6 = (M4xnv6 & Pj1ov6);
assign Vxoiw6 = (Jyoiw6 & Qyoiw6);
assign Jyoiw6 = (~(Xyoiw6 & Xloov6));
assign Xloov6 = (!J21ov6);
assign Xyoiw6 = (~(Wzcdt6 & D61ov6));
assign Xp38v6 = (~(Ezoiw6 & Lzoiw6));
assign Lzoiw6 = (~(Szoiw6 & Pj1ov6));
assign Ezoiw6 = (Zzoiw6 & G0piw6);
assign G0piw6 = (~(N0piw6 & U0piw6));
assign U0piw6 = (B1piw6 & Ldo7v6);
assign B1piw6 = (I1piw6 & V4jhw6);
assign I1piw6 = (~(P1piw6 & W1piw6));
assign W1piw6 = (~(Cgc7z6[0] & Qg2nv6));
assign N0piw6 = (D2piw6 & Cgc7z6[2]);
assign Zzoiw6 = (~(K2piw6 & R2piw6));
assign R2piw6 = (~(L7xnv6 | Y2piw6));
assign L7xnv6 = (N8xnv6 & Q0wnv6);
assign N8xnv6 = (Xg1ov6 & H11ov6);
assign Xg1ov6 = (F3piw6 & Kconv6);
assign F3piw6 = (~(Crcdt6 & M3piw6));
assign M3piw6 = (~(T3piw6 & Nlcdt6));
assign T3piw6 = (A4piw6 & H4piw6);
assign H4piw6 = (Fsc7z6[0] ^ Eh1ov6);
assign Eh1ov6 = (!Emoov6);
assign A4piw6 = (~(Fsc7z6[1] ^ Ghnov6));
assign K2piw6 = (Nbddt6 & O4piw6);
assign Qp38v6 = (V4piw6 & C5piw6);
assign C5piw6 = (J5piw6 & M4xnv6);
assign M4xnv6 = (!H11ov6);
assign J5piw6 = (~(IFLUSH | Sgcdt6));
assign V4piw6 = (Qyoiw6 & Q5piw6);
assign Q5piw6 = (~(L8oov6 & X5piw6));
assign X5piw6 = (~(J21ov6 & G2oov6));
assign J21ov6 = (E6piw6 & Cgc7z6[3]);
assign Qyoiw6 = (Ujnet6 | Tr9ov6);
assign Tr9ov6 = (X0oet6 & L6piw6);
assign L6piw6 = (~(S6piw6 & Z6piw6));
assign Z6piw6 = (~(G7piw6 & HRESPS[0]));
assign S6piw6 = (N7piw6 & U7piw6);
assign U7piw6 = (~(HRESPI[0] & B8piw6));
assign B8piw6 = (~(I8piw6 & P8piw6));
assign P8piw6 = (W8piw6 | D9piw6);
assign W8piw6 = (G7piw6 | K9piw6);
assign I8piw6 = (~(R9piw6 & Y9piw6));
assign Y9piw6 = (~(Fapiw6 & Hrb7z6[0]));
assign N7piw6 = (~(K9piw6 & Qhlov6));
assign Jp38v6 = (~(L3fov6 | Mapiw6));
assign L3fov6 = (Mjniw6 & Vzgov6);
assign Cp38v6 = (~(Tapiw6 & Abpiw6));
assign Abpiw6 = (~(S6cdt6 & Dcnov6));
assign Tapiw6 = (Vs9ov6 | V9i8v6);
assign V9i8v6 = (Xolhw6 & Trnov6);
assign Trnov6 = (~(Vs9ov6 | T7mov6));
assign Vo38v6 = (Dcnov6 ? Usbdt6 : Hbpiw6);
assign Oo38v6 = (~(Obpiw6 & Vbpiw6));
assign Vbpiw6 = (~(Ccpiw6 & Ple7z6[0]));
assign Obpiw6 = (Jcpiw6 & Qcpiw6);
assign Qcpiw6 = (~(Udkov6 & C5jhw6));
assign C5jhw6 = (~(Xcpiw6 & Edpiw6));
assign Edpiw6 = (~(Dfkov6 & Ldpiw6));
assign Ldpiw6 = (~(Sdpiw6 & Zdpiw6));
assign Zdpiw6 = (~(Z4hdt6 & Gepiw6));
assign Xcpiw6 = (~(Bsgdt6 & Nepiw6));
assign Jcpiw6 = (Uepiw6 | Xzhhw6);
assign Xzhhw6 = (Bfpiw6 & Ifpiw6);
assign Ifpiw6 = (Pfpiw6 & Wfpiw6);
assign Wfpiw6 = (~(Uqd7z6[22] & Dgpiw6));
assign Pfpiw6 = (Kgpiw6 & Rgpiw6);
assign Kgpiw6 = (~(Zec7z6[6] & Ygpiw6));
assign Bfpiw6 = (Fhpiw6 & Htfhw6);
assign Htfhw6 = (!Mhpiw6);
assign Fhpiw6 = (Thpiw6 & Aipiw6);
assign Aipiw6 = (~(Ovbdt6 & Hipiw6));
assign Thpiw6 = (~(Zec7z6[0] & Oipiw6));
assign Ho38v6 = (~(Vipiw6 & Cjpiw6));
assign Cjpiw6 = (~(Jjpiw6 & Dxghw6));
assign Dxghw6 = (~(Qjpiw6 & Xjpiw6));
assign Xjpiw6 = (Ekpiw6 & Lkpiw6);
assign Lkpiw6 = (Skpiw6 & Zkpiw6);
assign Zkpiw6 = (Glpiw6 | S9nhw6);
assign Skpiw6 = (Dsehw6 | B2phw6);
assign Ekpiw6 = (Nlpiw6 & Ulpiw6);
assign Ulpiw6 = (~(Zec7z6[7] & Oipiw6));
assign Nlpiw6 = (~(Hipiw6 & Oenhw6));
assign Qjpiw6 = (Bmpiw6 & Impiw6);
assign Impiw6 = (Pmpiw6 & Wmpiw6);
assign Wmpiw6 = (~(Q1s8v6 & J7ohw6));
assign Pmpiw6 = (Fcinv6 | E7phw6);
assign Bmpiw6 = (Dnpiw6 & Knpiw6);
assign Knpiw6 = (~(Zec7z6[5] & Zwlhw6));
assign Vipiw6 = (~(Ple7z6[7] & Ccpiw6));
assign Ao38v6 = (~(Rnpiw6 & Ynpiw6));
assign Ynpiw6 = (~(Jjpiw6 & C0hhw6));
assign C0hhw6 = (~(Fopiw6 & Mopiw6));
assign Mopiw6 = (Topiw6 & Appiw6);
assign Appiw6 = (Hppiw6 & Oppiw6);
assign Oppiw6 = (~(Ryr8v6 & J7ohw6));
assign Hppiw6 = (Vppiw6 & Cqpiw6);
assign Cqpiw6 = (~(Jqpiw6 & Zec7z6[10]));
assign Vppiw6 = (~(Uqd7z6[22] & Hipiw6));
assign Topiw6 = (Qqpiw6 & Xqpiw6);
assign Xqpiw6 = (~(Zec7z6[4] & Zwlhw6));
assign Qqpiw6 = (~(Zec7z6[6] & Oipiw6));
assign Fopiw6 = (Erpiw6 & Lrpiw6);
assign Lrpiw6 = (Srpiw6 & Zrpiw6);
assign Zrpiw6 = (Zpehw6 | E7phw6);
assign Srpiw6 = (Gspiw6 & Nspiw6);
assign Nspiw6 = (E9onv6 | B2phw6);
assign Gspiw6 = (Dsehw6 | S9nhw6);
assign Erpiw6 = (Qufhw6 & Uspiw6);
assign Uspiw6 = (~(Btpiw6 & Zec7z6[9]));
assign Rnpiw6 = (~(Ple7z6[6] & Ccpiw6));
assign Tn38v6 = (~(Itpiw6 & Ptpiw6));
assign Ptpiw6 = (Uepiw6 | Y4hhw6);
assign Y4hhw6 = (Wtpiw6 & Dupiw6);
assign Dupiw6 = (Kupiw6 & Rupiw6);
assign Rupiw6 = (Yupiw6 & Fvpiw6);
assign Fvpiw6 = (Mvpiw6 & Tvpiw6);
assign Tvpiw6 = (~(Awpiw6 & Hwpiw6));
assign Awpiw6 = (Owpiw6 & Vwpiw6);
assign Vwpiw6 = (Dsehw6 ^ E9onv6);
assign Mvpiw6 = (O0nhw6 | Rktov6);
assign Yupiw6 = (Cxpiw6 & Jxpiw6);
assign Jxpiw6 = (~(Jqpiw6 & Zec7z6[9]));
assign Cxpiw6 = (~(Uqd7z6[21] & Hipiw6));
assign Kupiw6 = (Qxpiw6 & Xxpiw6);
assign Xxpiw6 = (~(Zec7z6[5] & Oipiw6));
assign Qxpiw6 = (Eypiw6 & Lypiw6);
assign Lypiw6 = (~(Svr8v6 & J7ohw6));
assign Eypiw6 = (~(Zec7z6[3] & Zwlhw6));
assign Wtpiw6 = (Sypiw6 & Zypiw6);
assign Zypiw6 = (Gzpiw6 & Nzpiw6);
assign Nzpiw6 = (Qtnov6 | E7phw6);
assign Gzpiw6 = (Uzpiw6 & B0qiw6);
assign B0qiw6 = (Fjohw6 | B2phw6);
assign Uzpiw6 = (E9onv6 | S9nhw6);
assign Sypiw6 = (I0qiw6 & P0qiw6);
assign I0qiw6 = (W0qiw6 & D1qiw6);
assign D1qiw6 = (~(K1qiw6 & Zec7z6[10]));
assign W0qiw6 = (~(Btpiw6 & Zec7z6[7]));
assign Itpiw6 = (~(Ccpiw6 & Ple7z6[5]));
assign Mn38v6 = (~(R1qiw6 & Y1qiw6));
assign Y1qiw6 = (~(Ccpiw6 & Ple7z6[4]));
assign R1qiw6 = (F2qiw6 & M2qiw6);
assign M2qiw6 = (~(Udkov6 & J5jhw6));
assign J5jhw6 = (T2qiw6 | A3qiw6);
assign A3qiw6 = (Dfkov6 & H3qiw6);
assign H3qiw6 = (~(O3qiw6 & V3qiw6));
assign V3qiw6 = (~(Jwgdt6 & C4qiw6));
assign C4qiw6 = (J4qiw6 | Nygdt6);
assign T2qiw6 = (Mpe7z6[4] ? X4qiw6 : Q4qiw6);
assign X4qiw6 = (~(E5qiw6 | L5qiw6));
assign F2qiw6 = (~(Jjpiw6 & Wahhw6));
assign Wahhw6 = (~(S5qiw6 & Z5qiw6));
assign Z5qiw6 = (G6qiw6 & N6qiw6);
assign N6qiw6 = (U6qiw6 & B7qiw6);
assign B7qiw6 = (I7qiw6 & P7qiw6);
assign P7qiw6 = (~(Zec7z6[10] & W7qiw6));
assign I7qiw6 = (~(Jqpiw6 & Zec7z6[8]));
assign U6qiw6 = (D8qiw6 & K8qiw6);
assign K8qiw6 = (~(Uqd7z6[20] & Hipiw6));
assign D8qiw6 = (~(Zec7z6[30] & Dgpiw6));
assign G6qiw6 = (R8qiw6 & Y8qiw6);
assign Y8qiw6 = (T6onv6 | Dsehw6);
assign R8qiw6 = (F9qiw6 & M9qiw6);
assign M9qiw6 = (~(Tsr8v6 & J7ohw6));
assign F9qiw6 = (~(Zec7z6[2] & Zwlhw6));
assign S5qiw6 = (T9qiw6 & Aaqiw6);
assign Aaqiw6 = (Haqiw6 & Oaqiw6);
assign Oaqiw6 = (Vaqiw6 & Cbqiw6);
assign Cbqiw6 = (~(Zec7z6[4] & Oipiw6));
assign Vaqiw6 = (Jbqiw6 | B2phw6);
assign Haqiw6 = (Qbqiw6 & Xbqiw6);
assign Xbqiw6 = (Fjohw6 | S9nhw6);
assign Qbqiw6 = (U2ohw6 | E7phw6);
assign T9qiw6 = (Ecqiw6 & Lvfhw6);
assign Lvfhw6 = (!Lcqiw6);
assign Ecqiw6 = (Scqiw6 & Zcqiw6);
assign Zcqiw6 = (~(K1qiw6 & Zec7z6[9]));
assign Scqiw6 = (~(Btpiw6 & Zec7z6[6]));
assign Fn38v6 = (~(Gdqiw6 & Ndqiw6));
assign Ndqiw6 = (~(Ccpiw6 & Ple7z6[3]));
assign Gdqiw6 = (Udqiw6 & Beqiw6);
assign Beqiw6 = (~(Udkov6 & Q5jhw6));
assign Q5jhw6 = (~(Ieqiw6 & Peqiw6));
assign Peqiw6 = (~(Dfkov6 & Weqiw6));
assign Weqiw6 = (Nygdt6 ^ Dfqiw6);
assign Ieqiw6 = (Kfqiw6 & Wekov6);
assign Wekov6 = (!Q4qiw6);
assign Q4qiw6 = (Nepiw6 & L5qiw6);
assign L5qiw6 = (~(Mpe7z6[3] | Mpe7z6[2]));
assign Kfqiw6 = (~(Rfqiw6 & Mpe7z6[3]));
assign Rfqiw6 = (Mpe7z6[2] & Nepiw6);
assign Udqiw6 = (Uepiw6 | Vdhhw6);
assign Vdhhw6 = (Yfqiw6 & Fgqiw6);
assign Fgqiw6 = (Mgqiw6 & Tgqiw6);
assign Tgqiw6 = (Ahqiw6 & Hhqiw6);
assign Hhqiw6 = (Ohqiw6 & Vhqiw6);
assign Vhqiw6 = (~(J7ohw6 & Uonhw6));
assign Uonhw6 = (Nas8v6 & M6nhw6);
assign Ohqiw6 = (~(Zec7z6[9] & W7qiw6));
assign Ahqiw6 = (Ciqiw6 & Jiqiw6);
assign Jiqiw6 = (~(Jqpiw6 & Zec7z6[7]));
assign Ciqiw6 = (~(Uqd7z6[19] & Hipiw6));
assign Mgqiw6 = (Qiqiw6 & Xiqiw6);
assign Xiqiw6 = (T6onv6 | E9onv6);
assign Qiqiw6 = (Ejqiw6 & Ljqiw6);
assign Ljqiw6 = (~(Dgpiw6 & M6nhw6));
assign Ejqiw6 = (~(Zec7z6[1] & Zwlhw6));
assign Yfqiw6 = (Sjqiw6 & Zjqiw6);
assign Zjqiw6 = (Gkqiw6 & Nkqiw6);
assign Nkqiw6 = (Ukqiw6 & Blqiw6);
assign Blqiw6 = (~(Zec7z6[3] & Oipiw6));
assign Ukqiw6 = (Jgtov6 | B2phw6);
assign Gkqiw6 = (Ilqiw6 & Plqiw6);
assign Plqiw6 = (Jbqiw6 | S9nhw6);
assign Ilqiw6 = (T5ohw6 | E7phw6);
assign Sjqiw6 = (Wlqiw6 & Dmqiw6);
assign Wlqiw6 = (Kmqiw6 & Rmqiw6);
assign Rmqiw6 = (~(K1qiw6 & Zec7z6[8]));
assign Kmqiw6 = (~(Btpiw6 & Zec7z6[5]));
assign Ym38v6 = (~(Ymqiw6 & Fnqiw6));
assign Fnqiw6 = (~(Ccpiw6 & Ple7z6[2]));
assign Ymqiw6 = (Mnqiw6 & Tnqiw6);
assign Tnqiw6 = (~(Udkov6 & X5jhw6));
assign X5jhw6 = (~(Aoqiw6 & Hoqiw6));
assign Hoqiw6 = (~(Dfkov6 & Ooqiw6));
assign Ooqiw6 = (~(J4qiw6 & Voqiw6));
assign Voqiw6 = (~(R0hdt6 & Cpqiw6));
assign J4qiw6 = (!Dfqiw6);
assign Aoqiw6 = (E5qiw6 | Mpe7z6[2]);
assign Mnqiw6 = (~(Jjpiw6 & Kphhw6));
assign Kphhw6 = (~(Jpqiw6 & Qpqiw6));
assign Qpqiw6 = (Xpqiw6 & Eqqiw6);
assign Eqqiw6 = (Lqqiw6 & Sqqiw6);
assign Sqqiw6 = (Zqqiw6 & Grqiw6);
assign Grqiw6 = (~(Asnhw6 & J7ohw6));
assign Asnhw6 = (O7s8v6 & M6nhw6);
assign Zqqiw6 = (~(Jqpiw6 & Zec7z6[6]));
assign Jqpiw6 = (~(Nrqiw6 | Zec7z6[12]));
assign Lqqiw6 = (Urqiw6 & Bsqiw6);
assign Bsqiw6 = (~(Uqd7z6[18] & Hipiw6));
assign Urqiw6 = (~(Zec7z6[8] & Ygpiw6));
assign Xpqiw6 = (Isqiw6 & Psqiw6);
assign Psqiw6 = (~(Zec7z6[2] & Oipiw6));
assign Isqiw6 = (Wsqiw6 & Dtqiw6);
assign Dtqiw6 = (~(Dgpiw6 & Z9nhw6));
assign Wsqiw6 = (~(Zec7z6[0] & Zwlhw6));
assign Jpqiw6 = (Ktqiw6 & Rtqiw6);
assign Rtqiw6 = (Ytqiw6 & Fuqiw6);
assign Fuqiw6 = (S8ohw6 | E7phw6);
assign Ytqiw6 = (Muqiw6 & Tuqiw6);
assign Tuqiw6 = (Ctnov6 | B2phw6);
assign Muqiw6 = (Jgtov6 | S9nhw6);
assign Ktqiw6 = (Avqiw6 & Msfhw6);
assign Avqiw6 = (Hvqiw6 & Ovqiw6);
assign Ovqiw6 = (~(K1qiw6 & Zec7z6[7]));
assign Hvqiw6 = (~(Btpiw6 & Zec7z6[4]));
assign Rm38v6 = (~(Vvqiw6 & Cwqiw6));
assign Cwqiw6 = (~(Ccpiw6 & Ple7z6[1]));
assign Vvqiw6 = (Jwqiw6 & Qwqiw6);
assign Qwqiw6 = (~(Udkov6 & E6jhw6));
assign E6jhw6 = (~(Xwqiw6 & Exqiw6));
assign Exqiw6 = (~(Dfkov6 & Lxqiw6));
assign Lxqiw6 = (~(Cpqiw6 & Sxqiw6));
assign Sxqiw6 = (~(V2hdt6 & Sdpiw6));
assign Xwqiw6 = (L6jhw6 | E5qiw6);
assign E5qiw6 = (!Nepiw6);
assign Nepiw6 = (~(Dfkov6 | Mpe7z6[5]));
assign L6jhw6 = (!Xpgdt6);
assign Jwqiw6 = (~(Jjpiw6 & Ywhhw6));
assign Ywhhw6 = (~(Zxqiw6 & Gyqiw6));
assign Gyqiw6 = (Nyqiw6 & Uyqiw6);
assign Uyqiw6 = (Bzqiw6 & Izqiw6);
assign Izqiw6 = (~(Dgpiw6 & Oenhw6));
assign Dgpiw6 = (~(Pzqiw6 & Uqehw6));
assign Pzqiw6 = (Wzqiw6 & D0riw6);
assign Wzqiw6 = (O0nhw6 | K0riw6);
assign Bzqiw6 = (R0riw6 & Y0riw6);
assign Y0riw6 = (~(Uqd7z6[17] & Hipiw6));
assign Hipiw6 = (F1riw6 | Okohw6);
assign Okohw6 = (~(Prsov6 & Paohw6));
assign Paohw6 = (~(Mynhw6 & Xeinv6));
assign F1riw6 = (~(M1riw6 & T1riw6));
assign M1riw6 = (Yxnhw6 | Mqohw6);
assign Mqohw6 = (Kfa7z6 & M6nhw6);
assign Yxnhw6 = (~(A2riw6 & H2riw6));
assign R0riw6 = (~(Zec7z6[7] & Ygpiw6));
assign Ygpiw6 = (W7qiw6 | O2riw6);
assign O2riw6 = (!V2riw6);
assign W7qiw6 = (~(C3riw6 & J3riw6));
assign J3riw6 = (~(Rdfhw6 & Zec7z6[12]));
assign Nyqiw6 = (Q3riw6 & X3riw6);
assign X3riw6 = (~(Zunhw6 & J7ohw6));
assign J7ohw6 = (E4riw6 & Nvnhw6);
assign Nvnhw6 = (~(L4riw6 | H2riw6));
assign E4riw6 = (Zec7z6[10] & Zec7z6[30]);
assign Zunhw6 = (P4s8v6 & M6nhw6);
assign P4s8v6 = (C7t8v6 & Z9nhw6);
assign C7t8v6 = (~(Ctnov6 | Sfa7z6));
assign Q3riw6 = (~(Zec7z6[1] & Oipiw6));
assign Zxqiw6 = (S4riw6 & Z4riw6);
assign Z4riw6 = (G5riw6 & N5riw6);
assign N5riw6 = (~(K1qiw6 & Zec7z6[6]));
assign G5riw6 = (U5riw6 & B6riw6);
assign B6riw6 = (Ctnov6 | S9nhw6);
assign U5riw6 = (Baohw6 | E7phw6);
assign S4riw6 = (I6riw6 & P6riw6);
assign P6riw6 = (~(Btpiw6 & Zec7z6[3]));
assign Jjpiw6 = (!Uepiw6);
assign Uepiw6 = (Udkov6 | Ccpiw6);
assign Ccpiw6 = (~(W6riw6 | Udkov6));
assign Udkov6 = (D7riw6 & Bdf7z6[2]);
assign D7riw6 = (Bdf7z6[3] & Y4aov6);
assign Km38v6 = (K7riw6 | R7riw6);
assign K7riw6 = (Y7riw6 & Djgdt6);
assign Y7riw6 = (F8riw6 & M8riw6);
assign F8riw6 = (~(Ehgdt6 & Zbmnv6));
assign Zbmnv6 = (!T8riw6);
assign Dm38v6 = (~(A9riw6 & H9riw6));
assign H9riw6 = (~(O9riw6 & T8riw6));
assign O9riw6 = (Ehgdt6 & M8riw6);
assign A9riw6 = (~(V9riw6 & Cariw6));
assign Cariw6 = (~(Jariw6 & Qariw6));
assign Jariw6 = (~(W6riw6 & Xariw6));
assign Wl38v6 = (~(Ebriw6 & Lbriw6));
assign Lbriw6 = (Sbriw6 | Zbriw6);
assign Ebriw6 = (~(Dte7z6[0] & M8riw6));
assign Pl38v6 = (~(Gcriw6 & Ncriw6));
assign Ncriw6 = (~(Ucriw6 & Bdriw6));
assign Bdriw6 = (~(Idriw6 & Pdriw6));
assign Idriw6 = (Wdriw6 & Deriw6);
assign Gcriw6 = (~(Dte7z6[20] & M8riw6));
assign Il38v6 = (~(Keriw6 & Reriw6));
assign Reriw6 = (~(Ucriw6 & Yeriw6));
assign Yeriw6 = (~(Ffriw6 & Mfriw6));
assign Mfriw6 = (Tfriw6 & Agriw6);
assign Agriw6 = (~(Hgriw6 & Ogriw6));
assign Ogriw6 = (~(Vgriw6 & Chriw6));
assign Chriw6 = (Jhriw6 | H2riw6);
assign Vgriw6 = (Daphw6 & Dssov6);
assign Tfriw6 = (Qhriw6 & Xhriw6);
assign Ffriw6 = (Eiriw6 & Liriw6);
assign Eiriw6 = (Siriw6 & Wdriw6);
assign Keriw6 = (~(Dte7z6[19] & M8riw6));
assign Bl38v6 = (~(Ziriw6 & Gjriw6));
assign Gjriw6 = (~(Ucriw6 & Njriw6));
assign Njriw6 = (~(Ujriw6 & Bkriw6));
assign Bkriw6 = (Ikriw6 & Pkriw6);
assign Pkriw6 = (Qhriw6 & Wkriw6);
assign Qhriw6 = (~(Hgriw6 & Dlriw6));
assign Ikriw6 = (Klriw6 & Rlriw6);
assign Klriw6 = (~(Ylriw6 & Fmriw6));
assign Ylriw6 = (Hgriw6 & H2riw6);
assign Hgriw6 = (~(Qtnov6 | Mmriw6));
assign Ujriw6 = (Tmriw6 & Anriw6);
assign Tmriw6 = (V2riw6 & Aulhw6);
assign Ziriw6 = (~(Dte7z6[18] & M8riw6));
assign Uk38v6 = (Hnriw6 | Teliw6);
assign Hnriw6 = (N3onv6 ? Onriw6 : X0cdt6);
assign Onriw6 = (~(Vnriw6 & Coriw6));
assign Coriw6 = (Joriw6 & Qoriw6);
assign Qoriw6 = (~(Xoriw6 & Cyihw6));
assign Xoriw6 = (~(Epriw6 & Lpriw6));
assign Lpriw6 = (~(Spriw6 & S0ihw6));
assign Epriw6 = (~(Iwvnv6 & Dyfhw6));
assign Iwvnv6 = (Mqhhw6 & B8cdt6);
assign Joriw6 = (~(B8cdt6 & Zpriw6));
assign Zpriw6 = (~(Gqriw6 & Nqriw6));
assign Nqriw6 = (~(Uqriw6 & Brriw6));
assign Uqriw6 = (Oxihw6 & Irriw6);
assign Oxihw6 = (~(Prriw6 & Bylhw6));
assign Prriw6 = (Wrriw6 & Dsriw6);
assign Wrriw6 = (~(Ksriw6 & Zec7z6[5]));
assign Ksriw6 = (~(Rsriw6 | K0riw6));
assign Gqriw6 = (Ysriw6 & Ftriw6);
assign Ftriw6 = (~(Mtriw6 & Ttriw6));
assign Ttriw6 = (Auriw6 & Gifhw6);
assign Auriw6 = (Zhfhw6 & Shfhw6);
assign Mtriw6 = (~(Nifhw6 | Huriw6));
assign Huriw6 = (~(Ouriw6 | P6lhw6));
assign P6lhw6 = (Vuriw6 & Cvriw6);
assign Cvriw6 = (!Cyihw6);
assign Vuriw6 = (N3onv6 & Mzfhw6);
assign Mzfhw6 = (!Jvriw6);
assign Ysriw6 = (~(Qvriw6 & Xvriw6));
assign Xvriw6 = (Cyihw6 & F4ihw6);
assign Cyihw6 = (~(Ewriw6 & Lwriw6));
assign Lwriw6 = (Swriw6 & Yvihw6);
assign Swriw6 = (~(Zwriw6 | Gxriw6));
assign Ewriw6 = (Nxriw6 & Uxriw6);
assign Uxriw6 = (~(Zec7z6[4] & Byriw6));
assign Byriw6 = (~(Iyriw6 & Mefhw6));
assign Nxriw6 = (Pyriw6 & Wyriw6);
assign Wyriw6 = (~(Ydfhw6 & Dzriw6));
assign Dzriw6 = (Xgmhw6 | Kzriw6);
assign Pyriw6 = (~(Zec7z6[11] & Rzriw6));
assign Qvriw6 = (Wwvnv6 & Yzriw6);
assign Vnriw6 = (F0siw6 & M0siw6);
assign M0siw6 = (~(Spriw6 & Eilhw6));
assign Eilhw6 = (~(T0siw6 & A1siw6));
assign A1siw6 = (H1siw6 & O1siw6);
assign O1siw6 = (V1siw6 & C2siw6);
assign C2siw6 = (~(J2siw6 & Q2siw6));
assign Q2siw6 = (X2siw6 & E3siw6);
assign E3siw6 = (~(L3siw6 & Uqd7z6[20]));
assign L3siw6 = (Uqd7z6[18] & S3siw6);
assign X2siw6 = (~(Uqd7z6[19] & Z3siw6));
assign Z3siw6 = (~(G4siw6 & N4siw6));
assign N4siw6 = (~(Uqd7z6[17] & Ovbdt6));
assign G4siw6 = (Jbqiw6 & E9onv6);
assign J2siw6 = (U4siw6 & Kktov6);
assign V1siw6 = (B5siw6 & Xhriw6);
assign H1siw6 = (I5siw6 & P5siw6);
assign P5siw6 = (W5siw6 | D6siw6);
assign I5siw6 = (K6siw6 & R6siw6);
assign R6siw6 = (~(Y6siw6 & F7siw6));
assign F7siw6 = (M7siw6 & Rktov6);
assign Y6siw6 = (Tmsov6 & Ansov6);
assign K6siw6 = (~(T7siw6 & Gxlhw6));
assign Gxlhw6 = (~(A8siw6 & H8siw6));
assign H8siw6 = (O8siw6 & V8siw6);
assign V8siw6 = (C9siw6 & Daphw6);
assign Daphw6 = (!J9siw6);
assign C9siw6 = (Kaphw6 & Q9siw6);
assign O8siw6 = (O0nhw6 & Xosov6);
assign A8siw6 = (X9siw6 & Easiw6);
assign Easiw6 = (Lasiw6 & Sasiw6);
assign Lasiw6 = (Jhriw6 & Zasiw6);
assign Jhriw6 = (!Fmriw6);
assign X9siw6 = (Gbsiw6 & Nbsiw6);
assign T7siw6 = (~(Zec7z6[25] & Ubsiw6));
assign T0siw6 = (Bcsiw6 & Icsiw6);
assign Icsiw6 = (Pcsiw6 & Wcsiw6);
assign Pcsiw6 = (Ddsiw6 & S9nhw6);
assign Bcsiw6 = (Kdsiw6 & Rdsiw6);
assign Kdsiw6 = (Siriw6 & Ydsiw6);
assign Spriw6 = (Fesiw6 & Mesiw6);
assign Mesiw6 = (Tesiw6 & S4lhw6);
assign Tesiw6 = (L4lhw6 & Xehov6);
assign Fesiw6 = (~(I6lhw6 | Gaonv6));
assign Gaonv6 = (!B8cdt6);
assign F0siw6 = (~(X0cdt6 & V0onv6));
assign V0onv6 = (Afsiw6 & Hfsiw6);
assign Hfsiw6 = (Pxfov6 & Ofsiw6);
assign Afsiw6 = (Ecc7z6[3] & Pbadt6);
assign Nk38v6 = (Vfsiw6 ? Oyfdt6 : Ofsiw6);
assign Ofsiw6 = (Cgsiw6 | S0jnv6);
assign Gk38v6 = (~(Jgsiw6 & Qgsiw6));
assign Qgsiw6 = (~(Xgsiw6 & Ohe7z6[7]));
assign Jgsiw6 = (~(Vfsiw6 & Mfe7z6[7]));
assign Zj38v6 = (~(Ehsiw6 & Lhsiw6));
assign Lhsiw6 = (~(Xgsiw6 & Ohe7z6[6]));
assign Ehsiw6 = (~(Vfsiw6 & Mfe7z6[6]));
assign Sj38v6 = (~(Shsiw6 & Zhsiw6));
assign Zhsiw6 = (~(Xgsiw6 & Ohe7z6[5]));
assign Shsiw6 = (~(Vfsiw6 & Mfe7z6[5]));
assign Lj38v6 = (~(Gisiw6 & Nisiw6));
assign Nisiw6 = (~(Xgsiw6 & N0gdt6));
assign Gisiw6 = (~(Vfsiw6 & Mfe7z6[4]));
assign Ej38v6 = (~(Uisiw6 & Bjsiw6));
assign Bjsiw6 = (~(Xgsiw6 & Ohe7z6[4]));
assign Xgsiw6 = (~(Vfsiw6 | Sa2nv6));
assign Uisiw6 = (~(Vfsiw6 & Mfe7z6[3]));
assign Vfsiw6 = (Upfov6 & Ijsiw6);
assign Ijsiw6 = (~(N3onv6 & Oyfdt6));
assign Upfov6 = (Pjsiw6 & Wjsiw6);
assign Wjsiw6 = (Dksiw6 & P5mov6);
assign P5mov6 = (~(N3onv6 & Kksiw6));
assign Kksiw6 = (~(W4onv6 & G4mov6));
assign Dksiw6 = (Rksiw6 & Yksiw6);
assign Yksiw6 = (~(Flsiw6 & Mlsiw6));
assign Flsiw6 = (~(Wqfov6 | Tlsiw6));
assign Tlsiw6 = (!Ohe7z6[4]);
assign Rksiw6 = (!N4mov6);
assign N4mov6 = (Amsiw6 & Mlsiw6);
assign Mlsiw6 = (Hmsiw6 & Fsfov6);
assign Fsfov6 = (Omsiw6 & Vmsiw6);
assign Omsiw6 = (Cnsiw6 & Jnsiw6);
assign Cnsiw6 = (~(Qg2nv6 & Qnsiw6));
assign Qnsiw6 = (~(Xnsiw6 & Eosiw6));
assign Eosiw6 = (Losiw6 & Sosiw6);
assign Xnsiw6 = (Gd77z6 & Zosiw6);
assign Hmsiw6 = (~(Gpsiw6 | Npsiw6));
assign Npsiw6 = (Upsiw6 & Bqsiw6);
assign Bqsiw6 = (~(Iqsiw6 & N3onv6));
assign Iqsiw6 = (W4onv6 & Qg2nv6);
assign Upsiw6 = (~(Teliw6 & Pqsiw6));
assign Pqsiw6 = (Wqsiw6 | Drsiw6);
assign Amsiw6 = (Krsiw6 & Wqfov6);
assign Pjsiw6 = (Rrsiw6 & M0mov6);
assign M0mov6 = (Yrsiw6 & Fssiw6);
assign Fssiw6 = (~(Mssiw6 | Zo1ov6));
assign Mssiw6 = (Tssiw6 & Atsiw6);
assign Atsiw6 = (~(Htsiw6 & Otsiw6));
assign Tssiw6 = (~(Elphw6 & Vtsiw6));
assign Vtsiw6 = (~(Gmphw6 & Cusiw6));
assign Cusiw6 = (~(Mq9iw6 & Jusiw6));
assign Jusiw6 = (~(Qusiw6 & Ijmov6));
assign Yrsiw6 = (Xusiw6 & Evsiw6);
assign Evsiw6 = (~(Lvsiw6 & Gmphw6));
assign Gmphw6 = (Gr2et6 & Otsiw6);
assign Lvsiw6 = (Svsiw6 & Yioov6);
assign Svsiw6 = (~(Zvsiw6 & Xlinv6));
assign Xlinv6 = (Rhphw6 | Bwvnv6);
assign Zvsiw6 = (Gwsiw6 | Dwb7z6[5]);
assign Xusiw6 = (~(Xtvnv6 & Nwsiw6));
assign Nwsiw6 = (~(Uwsiw6 & Bxsiw6));
assign Bxsiw6 = (~(Ixsiw6 & Pxsiw6));
assign Pxsiw6 = (Bfo7v6 & Qtvnv6);
assign Ixsiw6 = (Wxsiw6 & Gr2et6);
assign Uwsiw6 = (~(Dysiw6 & C0ydt6));
assign C0ydt6 = (~(Qg2nv6 & Kysiw6));
assign Kysiw6 = (~(Hbo7v6 & Xsinv6));
assign Xtvnv6 = (~(Rysiw6 | Htsiw6));
assign Htsiw6 = (Yysiw6 & Fzsiw6);
assign Fzsiw6 = (~(L2nov6 | Mzmov6));
assign Yysiw6 = (~(Gwmov6 | Y5nov6));
assign Rrsiw6 = (Mzsiw6 & Po9iw6);
assign Po9iw6 = (~(F02nv6 & Qu1ov6));
assign Mzsiw6 = (~(Tzsiw6 & A0tiw6));
assign A0tiw6 = (~(F02nv6 | Yrfov6));
assign Tzsiw6 = (~(Krsiw6 | H0tiw6));
assign Krsiw6 = (Wqsiw6 | Rihov6);
assign Xi38v6 = (~(O0tiw6 & V0tiw6));
assign V0tiw6 = (~(Dte7z6[17] & M8riw6));
assign Qi38v6 = (C1tiw6 | J1tiw6);
assign J1tiw6 = (Dte7z6[16] & M8riw6);
assign Ji38v6 = (Q1tiw6 | X1tiw6);
assign X1tiw6 = (Dte7z6[15] & M8riw6);
assign Ci38v6 = (~(E2tiw6 & L2tiw6));
assign L2tiw6 = (~(Dte7z6[14] & M8riw6));
assign Vh38v6 = (~(S2tiw6 & Z2tiw6));
assign Z2tiw6 = (~(Dte7z6[13] & M8riw6));
assign Oh38v6 = (~(G3tiw6 & N3tiw6));
assign N3tiw6 = (~(D3bov6 & S7f7z6[1]));
assign G3tiw6 = (U3tiw6 & B4tiw6);
assign Hh38v6 = (~(P2bov6 & I4tiw6));
assign I4tiw6 = (~(D3bov6 & S7f7z6[2]));
assign Ah38v6 = (~(P4tiw6 & W4tiw6));
assign W4tiw6 = (D5tiw6 & B4tiw6);
assign B4tiw6 = (~(K5tiw6 & R5tiw6));
assign K5tiw6 = (~(Y5tiw6 | I4a7z6));
assign D5tiw6 = (F6tiw6 | Q4a7z6);
assign P4tiw6 = (P2bov6 & M6tiw6);
assign M6tiw6 = (~(D3bov6 & S7f7z6[3]));
assign Tg38v6 = (~(T6tiw6 & A7tiw6));
assign A7tiw6 = (~(D3bov6 & S7f7z6[4]));
assign T6tiw6 = (H7tiw6 & U3tiw6);
assign U3tiw6 = (~(O7tiw6 & V7tiw6));
assign V7tiw6 = (~(Rsi8v6 | I4a7z6));
assign O7tiw6 = (Abo7v6 & Y5tiw6);
assign H7tiw6 = (F6tiw6 | Y5tiw6);
assign Mg38v6 = (~(C8tiw6 & P2bov6));
assign P2bov6 = (Abo7v6 ? Q8tiw6 : J8tiw6);
assign Q8tiw6 = (~(X8tiw6 & Y5tiw6));
assign Y5tiw6 = (!Q4a7z6);
assign Q4a7z6 = (S9tiw6 ? L9tiw6 : E9tiw6);
assign L9tiw6 = (~(Z9tiw6 & Gatiw6));
assign Gatiw6 = (Natiw6 & Uatiw6);
assign Uatiw6 = (Bbtiw6 & Qariw6);
assign Bbtiw6 = (Ibtiw6 | Pbtiw6);
assign Natiw6 = (Wbtiw6 & Dctiw6);
assign Dctiw6 = (~(E9tiw6 & Kctiw6));
assign Kctiw6 = (~(Rctiw6 & Yctiw6));
assign Rctiw6 = (Fdtiw6 & Mdtiw6);
assign Fdtiw6 = (~(Tdtiw6 & Aetiw6));
assign Wbtiw6 = (~(Hetiw6 & Oetiw6));
assign Oetiw6 = (~(Vetiw6 & Cftiw6));
assign Cftiw6 = (Jftiw6 & Qftiw6);
assign Jftiw6 = (Xftiw6 | Egtiw6);
assign Vetiw6 = (Lgtiw6 & Sgtiw6);
assign Sgtiw6 = (Zgtiw6 | Ghtiw6);
assign Z9tiw6 = (Nhtiw6 & Uhtiw6);
assign Uhtiw6 = (Bitiw6 & Iitiw6);
assign Iitiw6 = (~(Ijnnv6 & Kfkov6));
assign Kfkov6 = (~(O3qiw6 ^ Fugdt6));
assign O3qiw6 = (~(Pitiw6 & Dfqiw6));
assign Dfqiw6 = (~(Cpqiw6 | R0hdt6));
assign Cpqiw6 = (Sdpiw6 | V2hdt6);
assign Sdpiw6 = (Gepiw6 | Z4hdt6);
assign Pitiw6 = (~(Nygdt6 | Jwgdt6));
assign Nhtiw6 = (Dfkov6 & Witiw6);
assign X8tiw6 = (Djtiw6 & I4a7z6);
assign J8tiw6 = (I4a7z6 | Kjtiw6);
assign Kjtiw6 = (~(Rsi8v6 | Rjtiw6));
assign Rsi8v6 = (!Djtiw6);
assign C8tiw6 = (Yjtiw6 & F6tiw6);
assign F6tiw6 = (~(R5tiw6 & I4a7z6));
assign I4a7z6 = (S9tiw6 ? Mktiw6 : Fktiw6);
assign Mktiw6 = (~(Tktiw6 & Altiw6));
assign Altiw6 = (Hltiw6 & Oltiw6);
assign Oltiw6 = (Vltiw6 & Cmtiw6);
assign Vltiw6 = (~(Jmtiw6 & Qmtiw6));
assign Qmtiw6 = (Xmtiw6 & Xftiw6);
assign Xmtiw6 = (Entiw6 & Lntiw6);
assign Jmtiw6 = (Hetiw6 & Qftiw6);
assign Hltiw6 = (Sntiw6 & Zntiw6);
assign Zntiw6 = (~(Gotiw6 & Notiw6));
assign Gotiw6 = (Ibtiw6 & R4aov6);
assign Ibtiw6 = (~(Uotiw6 & Egtiw6));
assign Sntiw6 = (~(Fktiw6 & Bptiw6));
assign Bptiw6 = (~(Iptiw6 & Pptiw6));
assign Pptiw6 = (~(Wptiw6 & Dqtiw6));
assign Wptiw6 = (Zgtiw6 & Aetiw6);
assign Tktiw6 = (Kqtiw6 & Witiw6);
assign Witiw6 = (Rqtiw6 & Yqtiw6);
assign Rqtiw6 = (~(Frtiw6 & Mrtiw6));
assign Mrtiw6 = (!Trtiw6);
assign Kqtiw6 = (Astiw6 & Hstiw6);
assign Hstiw6 = (~(Mpe7z6[5] & Y3bov6));
assign Fktiw6 = (E9tiw6 | Ouriw6);
assign Ouriw6 = (Rjtiw6 & Ostiw6);
assign Ostiw6 = (S2tiw6 ^ E2tiw6);
assign R5tiw6 = (Djtiw6 & Vstiw6);
assign Djtiw6 = (S9tiw6 ? Jttiw6 : Cttiw6);
assign Jttiw6 = (Qttiw6 & Xttiw6);
assign Xttiw6 = (Eutiw6 & Lutiw6);
assign Lutiw6 = (Cttiw6 | Iptiw6);
assign Iptiw6 = (Yctiw6 & E4lhw6);
assign Yctiw6 = (Sutiw6 & Zutiw6);
assign Zutiw6 = (~(Gvtiw6 | Nvtiw6));
assign Sutiw6 = (Uvtiw6 & Ol8iw6);
assign Eutiw6 = (Bwtiw6 & Z6jhw6);
assign Bwtiw6 = (~(Iwtiw6 & Zgtiw6));
assign Iwtiw6 = (~(Qariw6 & Pwtiw6));
assign Pwtiw6 = (Mdtiw6 | Cttiw6);
assign Qttiw6 = (Dfkov6 & Astiw6);
assign Astiw6 = (Wwtiw6 & Dxtiw6);
assign Wwtiw6 = (Kxtiw6 & Rxtiw6);
assign Rxtiw6 = (!Yxtiw6);
assign Cttiw6 = (~(E9tiw6 | Fytiw6));
assign Fytiw6 = (Q1tiw6 & Mytiw6);
assign E9tiw6 = (Tytiw6 & Rjtiw6);
assign Yjtiw6 = (~(D3bov6 & S7f7z6[0]));
assign D3bov6 = (Aztiw6 & Hztiw6);
assign Hztiw6 = (~(Oztiw6 | Rjtiw6));
assign Rjtiw6 = (Vztiw6 & C1tiw6);
assign Vztiw6 = (~(O0tiw6 | Q1tiw6));
assign Aztiw6 = (~(Ol8iw6 | Mytiw6));
assign Mytiw6 = (C0uiw6 & C1tiw6);
assign C0uiw6 = (J0uiw6 & E2tiw6);
assign J0uiw6 = (!O0tiw6);
assign O0tiw6 = (~(N3onv6 & Q0uiw6));
assign Q0uiw6 = (~(X0uiw6 & E1uiw6));
assign E1uiw6 = (L1uiw6 & S1uiw6);
assign L1uiw6 = (Z1uiw6 & G2uiw6);
assign X0uiw6 = (N2uiw6 & U2uiw6);
assign N2uiw6 = (Rdsiw6 & B3uiw6);
assign B3uiw6 = (~(K5onv6 & I3uiw6));
assign I3uiw6 = (~(P3uiw6 & Q9siw6));
assign Rdsiw6 = (W3uiw6 & D4uiw6);
assign D4uiw6 = (K4uiw6 & R4uiw6);
assign W3uiw6 = (Y4uiw6 & F5uiw6);
assign Fg38v6 = (~(M5uiw6 & T5uiw6));
assign T5uiw6 = (~(Y3bov6 & Yxf7z6[2]));
assign M5uiw6 = (A6uiw6 & H6uiw6);
assign H6uiw6 = (~(Rj2ov6 & Jamdt6));
assign A6uiw6 = (~(Yj2ov6 & Yxf7z6[6]));
assign Yf38v6 = (~(O6uiw6 & V6uiw6));
assign V6uiw6 = (~(Y3bov6 & Yxf7z6[6]));
assign O6uiw6 = (C7uiw6 & J7uiw6);
assign J7uiw6 = (~(Rj2ov6 & X1mdt6));
assign C7uiw6 = (~(Yj2ov6 & Yxf7z6[10]));
assign Rf38v6 = (~(Q7uiw6 & X7uiw6));
assign X7uiw6 = (~(Y3bov6 & Yxf7z6[10]));
assign Q7uiw6 = (E8uiw6 & L8uiw6);
assign L8uiw6 = (~(Rj2ov6 & Ltldt6));
assign E8uiw6 = (~(Yj2ov6 & Yxf7z6[14]));
assign Kf38v6 = (~(S8uiw6 & Z8uiw6));
assign Z8uiw6 = (~(Y3bov6 & Yxf7z6[14]));
assign S8uiw6 = (G9uiw6 & N9uiw6);
assign N9uiw6 = (~(Rj2ov6 & Zkldt6));
assign G9uiw6 = (~(Yj2ov6 & Yxf7z6[18]));
assign Df38v6 = (~(U9uiw6 & Bauiw6));
assign Bauiw6 = (~(Y3bov6 & Yxf7z6[18]));
assign U9uiw6 = (Iauiw6 & Pauiw6);
assign Pauiw6 = (~(Rj2ov6 & Ncldt6));
assign Iauiw6 = (~(Yj2ov6 & Yxf7z6[22]));
assign We38v6 = (~(Wauiw6 & Dbuiw6));
assign Dbuiw6 = (~(Y3bov6 & Yxf7z6[22]));
assign Wauiw6 = (Kbuiw6 & Rbuiw6);
assign Rbuiw6 = (~(Rj2ov6 & B4ldt6));
assign Kbuiw6 = (~(Yj2ov6 & Yxf7z6[26]));
assign Pe38v6 = (~(Ybuiw6 & Fcuiw6));
assign Fcuiw6 = (~(Y3bov6 & Yxf7z6[26]));
assign Ybuiw6 = (Mcuiw6 & Tcuiw6);
assign Tcuiw6 = (~(Rj2ov6 & Pvkdt6));
assign Mcuiw6 = (~(Yj2ov6 & Yxf7z6[30]));
assign Ie38v6 = (~(Aduiw6 & Hduiw6));
assign Hduiw6 = (~(Yj2ov6 & Yxf7z6[34]));
assign Aduiw6 = (~(Y3bov6 & Yxf7z6[30]));
assign Be38v6 = (~(Oduiw6 & Vduiw6));
assign Vduiw6 = (Wi2ov6 | Tmg7z6[32]);
assign Oduiw6 = (Ceuiw6 & Jeuiw6);
assign Jeuiw6 = (~(Rj2ov6 & Sgmdt6));
assign Ceuiw6 = (~(Yj2ov6 & Yxf7z6[3]));
assign Ud38v6 = (~(Qeuiw6 & Xeuiw6));
assign Xeuiw6 = (~(Y3bov6 & Yxf7z6[3]));
assign Qeuiw6 = (Efuiw6 & Lfuiw6);
assign Lfuiw6 = (~(Rj2ov6 & G8mdt6));
assign Efuiw6 = (~(Yj2ov6 & Yxf7z6[7]));
assign Nd38v6 = (~(Sfuiw6 & Zfuiw6));
assign Zfuiw6 = (~(Y3bov6 & Yxf7z6[7]));
assign Sfuiw6 = (Gguiw6 & Nguiw6);
assign Nguiw6 = (~(Rj2ov6 & Uzldt6));
assign Gguiw6 = (~(Yj2ov6 & Yxf7z6[11]));
assign Gd38v6 = (~(Uguiw6 & Bhuiw6));
assign Bhuiw6 = (~(Y3bov6 & Yxf7z6[11]));
assign Uguiw6 = (Ihuiw6 & Phuiw6);
assign Phuiw6 = (~(Rj2ov6 & Irldt6));
assign Ihuiw6 = (~(Yj2ov6 & Yxf7z6[15]));
assign Zc38v6 = (~(Whuiw6 & Diuiw6));
assign Diuiw6 = (~(Y3bov6 & Yxf7z6[15]));
assign Whuiw6 = (Kiuiw6 & Riuiw6);
assign Riuiw6 = (~(Rj2ov6 & Wildt6));
assign Kiuiw6 = (~(Yj2ov6 & Yxf7z6[19]));
assign Sc38v6 = (~(Yiuiw6 & Fjuiw6));
assign Fjuiw6 = (~(Y3bov6 & Yxf7z6[19]));
assign Yiuiw6 = (Mjuiw6 & Tjuiw6);
assign Tjuiw6 = (~(Rj2ov6 & Kaldt6));
assign Mjuiw6 = (~(Yj2ov6 & Yxf7z6[23]));
assign Lc38v6 = (~(Akuiw6 & Hkuiw6));
assign Hkuiw6 = (~(Y3bov6 & Yxf7z6[23]));
assign Akuiw6 = (Okuiw6 & Vkuiw6);
assign Vkuiw6 = (~(Rj2ov6 & Y1ldt6));
assign Okuiw6 = (~(Yj2ov6 & Yxf7z6[27]));
assign Ec38v6 = (~(Cluiw6 & Jluiw6));
assign Jluiw6 = (Rgpiw6 | Sbriw6);
assign Rgpiw6 = (~(Qluiw6 & Xluiw6));
assign Xluiw6 = (Uqd7z6[21] & Owpiw6);
assign Qluiw6 = (Hwpiw6 & Uqd7z6[20]);
assign Cluiw6 = (~(Dte7z6[12] & M8riw6));
assign Xb38v6 = (~(Emuiw6 & Lmuiw6));
assign Lmuiw6 = (Sbriw6 | Smuiw6);
assign Emuiw6 = (~(Dte7z6[11] & M8riw6));
assign Qb38v6 = (~(Zmuiw6 & Gnuiw6));
assign Gnuiw6 = (~(Ucriw6 & Nnuiw6));
assign Nnuiw6 = (~(Unuiw6 & Bouiw6));
assign Unuiw6 = (C3riw6 & A7onv6);
assign Zmuiw6 = (~(Dte7z6[10] & M8riw6));
assign Jb38v6 = (~(Iouiw6 & Pouiw6));
assign Pouiw6 = (~(Dte7z6[9] & M8riw6));
assign Iouiw6 = (~(Ucriw6 & Wouiw6));
assign Wouiw6 = (~(Dpuiw6 & Kpuiw6));
assign Kpuiw6 = (Rpuiw6 & Ypuiw6);
assign Ypuiw6 = (L4riw6 & Fquiw6);
assign Rpuiw6 = (Mquiw6 & M6onv6);
assign Dpuiw6 = (Tquiw6 & Aruiw6);
assign Tquiw6 = (L9onv6 & Bouiw6);
assign Cb38v6 = (~(Hruiw6 & Oruiw6));
assign Oruiw6 = (~(Ucriw6 & Vruiw6));
assign Vruiw6 = (~(Csuiw6 & Jsuiw6));
assign Jsuiw6 = (Qsuiw6 & Xsuiw6);
assign Xsuiw6 = (~(Etuiw6 & Zec7z6[5]));
assign Qsuiw6 = (Ltuiw6 & Stuiw6);
assign Csuiw6 = (Ztuiw6 & Guuiw6);
assign Ztuiw6 = (Nuuiw6 & Uuuiw6);
assign Uuuiw6 = (~(Bvuiw6 & Nbfhw6));
assign Nuuiw6 = (~(Uqd7z6[21] & Owpiw6));
assign Hruiw6 = (~(Dte7z6[7] & M8riw6));
assign Va38v6 = (~(Ivuiw6 & Pvuiw6));
assign Pvuiw6 = (~(Ucriw6 & Wvuiw6));
assign Wvuiw6 = (~(Dwuiw6 & Kwuiw6));
assign Kwuiw6 = (Rwuiw6 & Ywuiw6);
assign Ywuiw6 = (~(Fxuiw6 & V0nhw6));
assign Fxuiw6 = (Nbfhw6 & Mxuiw6);
assign Rwuiw6 = (Txuiw6 & Ayuiw6);
assign Txuiw6 = (~(Hyuiw6 & Oyuiw6));
assign Dwuiw6 = (Vyuiw6 & Guuiw6);
assign Guuiw6 = (Czuiw6 & Jzuiw6);
assign Jzuiw6 = (~(Bvuiw6 & Qzuiw6));
assign Czuiw6 = (Xzuiw6 & T6onv6);
assign Vyuiw6 = (E0viw6 & L0viw6);
assign L0viw6 = (~(Bvuiw6 & E3fhw6));
assign E0viw6 = (~(Uqd7z6[20] & Owpiw6));
assign Ivuiw6 = (~(Dte7z6[6] & M8riw6));
assign Oa38v6 = (~(S0viw6 & Z0viw6));
assign Z0viw6 = (~(G1viw6 & Fmriw6));
assign Fmriw6 = (~(L4riw6 | N1viw6));
assign G1viw6 = (~(Sbriw6 | H2riw6));
assign S0viw6 = (~(Dte7z6[5] & M8riw6));
assign Ha38v6 = (~(U1viw6 & B2viw6));
assign B2viw6 = (~(Ucriw6 & J9siw6));
assign U1viw6 = (~(Dte7z6[4] & M8riw6));
assign Aa38v6 = (~(I2viw6 & P2viw6));
assign P2viw6 = (~(Dte7z6[3] & M8riw6));
assign T938v6 = (~(W2viw6 & D3viw6));
assign D3viw6 = (Sbriw6 | K3viw6);
assign Sbriw6 = (!Ucriw6);
assign W2viw6 = (~(Dte7z6[2] & M8riw6));
assign M938v6 = (~(R3viw6 & Y3viw6));
assign Y3viw6 = (~(Ucriw6 & F4viw6));
assign F4viw6 = (~(M4viw6 & T4viw6));
assign T4viw6 = (A5viw6 & H5viw6);
assign H5viw6 = (O5viw6 & V5viw6);
assign V5viw6 = (Xhriw6 & C6viw6);
assign O5viw6 = (~(J6viw6 | Q6viw6));
assign A5viw6 = (X6viw6 & E7viw6);
assign E7viw6 = (L7viw6 & X9fhw6);
assign X6viw6 = (S7viw6 & Z7viw6);
assign M4viw6 = (G8viw6 & N8viw6);
assign N8viw6 = (U8viw6 & B9viw6);
assign B9viw6 = (I9viw6 & P9viw6);
assign I9viw6 = (~(W9viw6 & Daviw6));
assign W9viw6 = (Kaviw6 & Qtnov6);
assign U8viw6 = (Raviw6 & Yaviw6);
assign Yaviw6 = (W5siw6 | Gginv6);
assign Raviw6 = (~(Zafhw6 & V1fhw6));
assign G8viw6 = (Fbviw6 & Mbviw6);
assign Mbviw6 = (Tbviw6 & Acviw6);
assign Acviw6 = (Hcviw6 | Xeinv6);
assign Fbviw6 = (Zpsov6 & Ocviw6);
assign Zpsov6 = (Vcviw6 & Cdviw6);
assign Cdviw6 = (W5siw6 | Jdviw6);
assign Ucriw6 = (~(M8riw6 | Vs9ov6));
assign R3viw6 = (~(Dte7z6[1] & M8riw6));
assign F938v6 = (~(Qdviw6 & Xdviw6));
assign Xdviw6 = (~(Xwe7z6[1] & M8riw6));
assign Qdviw6 = (Eeviw6 & Leviw6);
assign Leviw6 = (~(Seviw6 & Gifhw6));
assign Gifhw6 = (~(Zeviw6 & Gfviw6));
assign Gfviw6 = (Nfviw6 | Bat8v6);
assign Zeviw6 = (Ufviw6 & Bgviw6);
assign Bgviw6 = (~(Uqd7z6[17] & Igviw6));
assign Ufviw6 = (~(Zec7z6[25] & Pgviw6));
assign Eeviw6 = (~(R7riw6 & Oac7z6[1]));
assign Y838v6 = (~(Wgviw6 & Dhviw6));
assign Dhviw6 = (~(Xwe7z6[2] & M8riw6));
assign Wgviw6 = (Khviw6 & Rhviw6);
assign Rhviw6 = (~(Seviw6 & Zhfhw6));
assign Zhfhw6 = (~(Yhviw6 & Fiviw6));
assign Fiviw6 = (~(Zec7z6[26] & Pgviw6));
assign Yhviw6 = (Miviw6 & Tiviw6);
assign Tiviw6 = (~(Uqd7z6[18] & Igviw6));
assign Miviw6 = (Adohw6 | Nfviw6);
assign Khviw6 = (~(R7riw6 & Oac7z6[2]));
assign R838v6 = (~(Ajviw6 & Hjviw6));
assign Hjviw6 = (~(Xwe7z6[3] & M8riw6));
assign Ajviw6 = (Ojviw6 & Vjviw6);
assign Vjviw6 = (~(Seviw6 & Shfhw6));
assign Shfhw6 = (~(Ckviw6 & Jkviw6));
assign Jkviw6 = (~(Zec7z6[27] & Pgviw6));
assign Ckviw6 = (Qkviw6 & Xkviw6);
assign Xkviw6 = (~(Uqd7z6[19] & Igviw6));
assign Qkviw6 = (Elviw6 | Nfviw6);
assign Ojviw6 = (~(R7riw6 & Oac7z6[3]));
assign K838v6 = (~(Llviw6 & Slviw6));
assign Slviw6 = (~(Xwe7z6[0] & M8riw6));
assign Llviw6 = (Zlviw6 & Gmviw6);
assign Gmviw6 = (~(Seviw6 & Nifhw6));
assign Nifhw6 = (~(Nmviw6 & Umviw6));
assign Umviw6 = (Nfviw6 | Kfa7z6);
assign Nfviw6 = (Bnviw6 & Inviw6);
assign Nmviw6 = (Pnviw6 & Wnviw6);
assign Wnviw6 = (~(Ovbdt6 & Igviw6));
assign Pnviw6 = (~(Zec7z6[24] & Pgviw6));
assign Seviw6 = (~(M8riw6 | Xariw6));
assign Zlviw6 = (~(R7riw6 & Oac7z6[0]));
assign R7riw6 = (W6riw6 & Xariw6);
assign W6riw6 = (!M8riw6);
assign M8riw6 = (~(Hmtov6 & Doviw6));
assign Doviw6 = (~(Koviw6 & Roviw6));
assign Roviw6 = (Tytiw6 & Yoviw6);
assign Yoviw6 = (~(Q1tiw6 | C1tiw6));
assign C1tiw6 = (N3onv6 & Fpviw6);
assign Fpviw6 = (~(Mpviw6 & Tpviw6));
assign Tpviw6 = (Aqviw6 & Hqviw6);
assign Hqviw6 = (~(M0fhw6 | Oqviw6));
assign Aqviw6 = (Vqviw6 & R4uiw6);
assign R4uiw6 = (Nqehw6 | Ubsiw6);
assign Vqviw6 = (~(Crviw6 & Jrviw6));
assign Jrviw6 = (!Kssov6);
assign Mpviw6 = (Qrviw6 & Xrviw6);
assign Qrviw6 = (F5uiw6 & Esviw6);
assign F5uiw6 = (Lsviw6 & Ssviw6);
assign Q1tiw6 = (N3onv6 & Zsviw6);
assign Zsviw6 = (~(Gtviw6 & Ntviw6));
assign Ntviw6 = (Utviw6 & Buviw6);
assign Utviw6 = (C3riw6 & Iuviw6);
assign Iuviw6 = (~(Puviw6 & K5onv6));
assign Puviw6 = (~(P3uiw6 & Sasiw6));
assign Sasiw6 = (Wuviw6 & Dvviw6);
assign Dvviw6 = (~(Bvuiw6 | Kvviw6));
assign Wuviw6 = (Rvviw6 & Yvviw6);
assign P3uiw6 = (Fwviw6 & Mwviw6);
assign Mwviw6 = (Twviw6 & Kaphw6);
assign Kaphw6 = (!Prehw6);
assign Prehw6 = (~(T6onv6 | Axviw6));
assign Axviw6 = (~(Nbfhw6 | Hxviw6));
assign Twviw6 = (~(Oxviw6 & Tmsov6));
assign Oxviw6 = (~(M0fhw6 | K0riw6));
assign M0fhw6 = (Vxviw6 & Tmsov6);
assign Tmsov6 = (!Hffhw6);
assign Vxviw6 = (Kssov6 & Rktov6);
assign Fwviw6 = (Vffhw6 & Cyviw6);
assign Cyviw6 = (~(U4siw6 & Ansov6));
assign Vffhw6 = (Jyviw6 & Qyviw6);
assign Qyviw6 = (Zasiw6 & L7viw6);
assign Jyviw6 = (Xyviw6 & S7viw6);
assign Xyviw6 = (~(Ezviw6 & Lzviw6));
assign Ezviw6 = (A2riw6 & K0riw6);
assign Gtviw6 = (Szviw6 & Y4uiw6);
assign Y4uiw6 = (Zzviw6 & G0wiw6);
assign G0wiw6 = (N0wiw6 & X9fhw6);
assign N0wiw6 = (~(V8fhw6 | Oqviw6));
assign Zzviw6 = (U0wiw6 & Aruiw6);
assign Aruiw6 = (B1wiw6 & Q9fhw6);
assign B1wiw6 = (I1wiw6 & Amtov6);
assign U0wiw6 = (~(P1wiw6 | Mtehw6));
assign Szviw6 = (W1wiw6 & D2wiw6);
assign Tytiw6 = (E2tiw6 & S2tiw6);
assign S2tiw6 = (~(N3onv6 & K2wiw6));
assign K2wiw6 = (~(R2wiw6 & Y2wiw6));
assign Y2wiw6 = (F3wiw6 & M3wiw6);
assign M3wiw6 = (T3wiw6 & Epsov6);
assign T3wiw6 = (A4wiw6 & H4wiw6);
assign F3wiw6 = (Lsviw6 & O4wiw6);
assign O4wiw6 = (~(Crviw6 & V4wiw6));
assign Crviw6 = (C5wiw6 & J5wiw6);
assign J5wiw6 = (~(Q5wiw6 | Ansov6));
assign C5wiw6 = (U4siw6 & Z1uiw6);
assign Lsviw6 = (X5wiw6 & E6wiw6);
assign X5wiw6 = (~(L6wiw6 & S6wiw6));
assign R2wiw6 = (Z6wiw6 & G7wiw6);
assign G7wiw6 = (N7wiw6 & Esviw6);
assign Esviw6 = (U7wiw6 & B8wiw6);
assign B8wiw6 = (~(P1wiw6 | Zbsov6));
assign P1wiw6 = (I8wiw6 & Uqd7z6[20]);
assign I8wiw6 = (X8onv6 & P8wiw6);
assign U7wiw6 = (D2wiw6 & W8wiw6);
assign W8wiw6 = (~(D9wiw6 & K5onv6));
assign D2wiw6 = (K9wiw6 & Ycnov6);
assign Ycnov6 = (~(Jhsov6 & Zec7z6[1]));
assign K9wiw6 = (~(R9wiw6 & Hftov6));
assign N7wiw6 = (Y9wiw6 & Fawiw6);
assign Fawiw6 = (~(Mawiw6 & Tawiw6));
assign Mawiw6 = (Abwiw6 | Hbwiw6);
assign Hbwiw6 = (Obwiw6 & Hxviw6);
assign Y9wiw6 = (Uqehw6 | Mmriw6);
assign Uqehw6 = (Rvviw6 & Xosov6);
assign Rvviw6 = (~(V0nhw6 & Nbfhw6));
assign Z6wiw6 = (Ocviw6 & U2uiw6);
assign U2uiw6 = (Vbwiw6 & Ccwiw6);
assign Ccwiw6 = (~(K5onv6 & Jcwiw6));
assign Jcwiw6 = (~(Qcwiw6 & Yvviw6));
assign Yvviw6 = (Xcwiw6 | Dsehw6);
assign Vbwiw6 = (~(U4siw6 & Kssov6));
assign Ocviw6 = (Edwiw6 & Ldwiw6);
assign Edwiw6 = (~(Sdwiw6 & E3fhw6));
assign Sdwiw6 = (Zdwiw6 & Tawiw6);
assign E2tiw6 = (~(N3onv6 & Gewiw6));
assign Gewiw6 = (~(Newiw6 & Uewiw6));
assign Uewiw6 = (Bfwiw6 & Ifwiw6);
assign Ifwiw6 = (Pfwiw6 & P9viw6);
assign P9viw6 = (~(Wfwiw6 & Rktov6));
assign Pfwiw6 = (Z7viw6 & H4wiw6);
assign Z7viw6 = (Dgwiw6 | K0riw6);
assign Bfwiw6 = (Kgwiw6 & Rgwiw6);
assign Rgwiw6 = (~(R9wiw6 & S3siw6));
assign S3siw6 = (!Hftov6);
assign Kgwiw6 = (E6wiw6 & V4wiw6);
assign V4wiw6 = (~(Ygwiw6 & Fhwiw6));
assign Fhwiw6 = (Ijtov6 & Kktov6);
assign E6wiw6 = (Q1ghw6 | Mhwiw6);
assign Newiw6 = (Thwiw6 & Aiwiw6);
assign Aiwiw6 = (Hiwiw6 & Oiwiw6);
assign Oiwiw6 = (~(Tawiw6 & Viwiw6));
assign Hiwiw6 = (Ssviw6 & Z1uiw6);
assign Z1uiw6 = (~(Cjwiw6 & Jjwiw6));
assign Jjwiw6 = (Ovbdt6 & Fjohw6);
assign Cjwiw6 = (U4siw6 & Qjwiw6);
assign Ssviw6 = (~(Xjwiw6 & L6wiw6));
assign Thwiw6 = (W1wiw6 & Ekwiw6);
assign W1wiw6 = (Lkwiw6 & Skwiw6);
assign Skwiw6 = (Zkwiw6 & S1uiw6);
assign S1uiw6 = (Mmriw6 | Nbsiw6);
assign Nbsiw6 = (Glwiw6 & Wrehw6);
assign Wrehw6 = (Nlwiw6 | E9onv6);
assign Glwiw6 = (Xcwiw6 | Uqd7z6[21]);
assign Xcwiw6 = (Nlwiw6 | Uqd7z6[20]);
assign Nlwiw6 = (~(Ulwiw6 & Bmwiw6));
assign Ulwiw6 = (Zec7z6[4] & Zpehw6);
assign Zkwiw6 = (~(Imwiw6 & K5onv6));
assign Imwiw6 = (~(Pmwiw6 & Wmwiw6));
assign Wmwiw6 = (Xosov6 & Q9siw6);
assign Q9siw6 = (!D9wiw6);
assign D9wiw6 = (Dnwiw6 & Knwiw6);
assign Knwiw6 = (Rnwiw6 & Zec7z6[4]);
assign Rnwiw6 = (E9onv6 & Dsehw6);
assign Dnwiw6 = (Bmwiw6 & Zec7z6[5]);
assign Xosov6 = (!Etuiw6);
assign Etuiw6 = (Ynwiw6 & V0nhw6);
assign Ynwiw6 = (Fowiw6 & Fcinv6);
assign Fowiw6 = (~(Hwpiw6 & Zec7z6[5]));
assign Pmwiw6 = (Qcwiw6 & O0nhw6);
assign O0nhw6 = (~(Mowiw6 & V0nhw6));
assign Mowiw6 = (Qzuiw6 & Xeinv6);
assign Qcwiw6 = (Zasiw6 | Xeinv6);
assign Zasiw6 = (~(Towiw6 & Mynhw6));
assign Towiw6 = (Nbfhw6 & Qtnov6);
assign Lkwiw6 = (Xrviw6 & K4uiw6);
assign Xrviw6 = (~(Apwiw6 | Q5wiw6));
assign Q5wiw6 = (Zhtov6 & R9wiw6);
assign R9wiw6 = (Ygwiw6 & Hpwiw6);
assign Hpwiw6 = (Gitov6 & Kktov6);
assign Ygwiw6 = (U4siw6 & Uqd7z6[20]);
assign U4siw6 = (~(Onlhw6 | Mmriw6));
assign Mmriw6 = (!K5onv6);
assign K5onv6 = (~(Opwiw6 & Zec7z6[25]));
assign Opwiw6 = (Ubsiw6 & Vpwiw6);
assign Vpwiw6 = (~(Tawiw6 & Cqwiw6));
assign Cqwiw6 = (~(Jqwiw6 & Qqwiw6));
assign Qqwiw6 = (~(Hxviw6 & Xqwiw6));
assign Jqwiw6 = (~(Abwiw6 | Erwiw6));
assign Tawiw6 = (!Wrsov6);
assign Zhtov6 = (Uqd7z6[17] & Ovbdt6);
assign Apwiw6 = (Jhsov6 & Zec7z6[0]);
assign Jhsov6 = (Lrwiw6 & Srwiw6);
assign Srwiw6 = (Zrwiw6 & Zec7z6[5]);
assign Lrwiw6 = (Ttehw6 & Cvehw6);
assign Koviw6 = (Gswiw6 & Xhlhw6);
assign Gswiw6 = (Nswiw6 & I2viw6);
assign I2viw6 = (~(N3onv6 & Uswiw6));
assign Uswiw6 = (~(Btwiw6 & Itwiw6));
assign Itwiw6 = (Ptwiw6 & L7viw6);
assign L7viw6 = (~(Wtwiw6 & K0riw6));
assign Wtwiw6 = (!Dgwiw6);
assign Dgwiw6 = (~(Duwiw6 & Qzuiw6));
assign Duwiw6 = (Owpiw6 & Zdwiw6);
assign Ptwiw6 = (X9fhw6 & Xhriw6);
assign Btwiw6 = (K3viw6 & S7viw6);
assign S7viw6 = (~(Wfwiw6 & K0riw6));
assign Wfwiw6 = (Kuwiw6 & A2riw6);
assign Kuwiw6 = (Qzuiw6 & Zdwiw6);
assign K3viw6 = (Ruwiw6 & Yuwiw6);
assign Yuwiw6 = (Fvwiw6 & Mvwiw6);
assign Mvwiw6 = (Tvwiw6 & S9nhw6);
assign Tvwiw6 = (B5siw6 & Wkriw6);
assign Fvwiw6 = (V2riw6 & Ddsiw6);
assign Ruwiw6 = (Awwiw6 & Hwwiw6);
assign Hwwiw6 = (Wdriw6 & Wcsiw6);
assign Awwiw6 = (Liriw6 & Gbsiw6);
assign Gbsiw6 = (~(Dlriw6 | Owwiw6));
assign Owwiw6 = (Vwwiw6 & Kaviw6);
assign Kaviw6 = (!Prsov6);
assign Vwwiw6 = (Cxwiw6 & Qtnov6);
assign Cxwiw6 = (Daviw6 | Abwiw6);
assign Abwiw6 = (Zdwiw6 & Hxviw6);
assign Daviw6 = (E3fhw6 & Zec7z6[7]);
assign Dlriw6 = (~(Jxwiw6 & Qxwiw6));
assign Qxwiw6 = (Xxwiw6 & Zbriw6);
assign Zbriw6 = (W9phw6 & Eywiw6);
assign Eywiw6 = (~(Lywiw6 & A2riw6));
assign Lywiw6 = (Sywiw6 & Nbfhw6);
assign W9phw6 = (~(Zywiw6 & Sywiw6));
assign Zywiw6 = (Owpiw6 & Nbfhw6);
assign Xxwiw6 = (~(Gzwiw6 | Mbphw6));
assign Mbphw6 = (Nzwiw6 & Hxviw6);
assign Gzwiw6 = (Uzwiw6 & A2riw6);
assign Uzwiw6 = (B0xiw6 & Hxviw6);
assign Jxwiw6 = (Pdriw6 & Tbviw6);
assign Tbviw6 = (Tbphw6 & I0xiw6);
assign I0xiw6 = (~(A2riw6 & Erwiw6));
assign Tbphw6 = (P0xiw6 & Deriw6);
assign Deriw6 = (~(Nzwiw6 & Qzuiw6));
assign P0xiw6 = (~(Erwiw6 & Owpiw6));
assign Pdriw6 = (W0xiw6 & D1xiw6);
assign D1xiw6 = (~(K1xiw6 & A2riw6));
assign K1xiw6 = (Nbfhw6 & B0xiw6);
assign W0xiw6 = (~(Fbphw6 | J6viw6));
assign J6viw6 = (R1xiw6 & A2riw6);
assign A2riw6 = (!L4riw6);
assign R1xiw6 = (Qzuiw6 & B0xiw6);
assign Fbphw6 = (Nzwiw6 & Nbfhw6);
assign Nzwiw6 = (~(D0riw6 | Y1xiw6));
assign Nswiw6 = (~(J9siw6 & N3onv6));
assign J9siw6 = (~(D0riw6 | N1viw6));
assign N1viw6 = (F2xiw6 & M2xiw6);
assign F2xiw6 = (!Viwiw6);
assign Viwiw6 = (~(T2xiw6 & A3xiw6));
assign A3xiw6 = (~(H3xiw6 & Zdwiw6));
assign H3xiw6 = (Nbfhw6 & Rktov6);
assign T2xiw6 = (~(Obwiw6 & Hxviw6));
assign Hmtov6 = (!Dcnov6);
assign D838v6 = (Sidiw6 ? U6i7z6[0] : O3xiw6);
assign O3xiw6 = (Vxihw6 & V3xiw6);
assign V3xiw6 = (~(C4xiw6 & J4xiw6));
assign J4xiw6 = (~(Q4xiw6 & Ecc7z6[11]));
assign Q4xiw6 = (Mwphw6 & Cwlnv6);
assign C4xiw6 = (~(X4xiw6 & E5xiw6));
assign E5xiw6 = (~(L5xiw6 & S5xiw6));
assign S5xiw6 = (~(Z5xiw6 & G6xiw6));
assign Z5xiw6 = (~(N6xiw6 | Ecc7z6[10]));
assign W738v6 = (~(U6xiw6 & B7xiw6));
assign B7xiw6 = (I7xiw6 & P7xiw6);
assign P7xiw6 = (~(Td2ov6 & W7xiw6));
assign I7xiw6 = (D8xiw6 & K8xiw6);
assign K8xiw6 = (C12ov6 | Utjnv6);
assign Utjnv6 = (R8xiw6 & Y8xiw6);
assign Y8xiw6 = (F9xiw6 & M9xiw6);
assign M9xiw6 = (T9xiw6 & Aaxiw6);
assign Aaxiw6 = (Haxiw6 & Oaxiw6);
assign Oaxiw6 = (~(vis_psp_o[26] & N32ov6));
assign Haxiw6 = (~(U32ov6 & Pic7z6[26]));
assign T9xiw6 = (Vaxiw6 & Cbxiw6);
assign Cbxiw6 = (~(vis_msp_o[26] & P42ov6));
assign Vaxiw6 = (~(vis_r12_o[26] & W42ov6));
assign F9xiw6 = (Jbxiw6 & Qbxiw6);
assign Qbxiw6 = (Xbxiw6 & Ecxiw6);
assign Ecxiw6 = (~(vis_r11_o[26] & F62ov6));
assign Xbxiw6 = (~(vis_r10_o[26] & M62ov6));
assign Jbxiw6 = (Lcxiw6 & Scxiw6);
assign Scxiw6 = (~(vis_r9_o[26] & H72ov6));
assign Lcxiw6 = (~(vis_r8_o[26] & O72ov6));
assign R8xiw6 = (Zcxiw6 & Gdxiw6);
assign Gdxiw6 = (Ndxiw6 & Udxiw6);
assign Udxiw6 = (Bexiw6 & Iexiw6);
assign Iexiw6 = (~(vis_r7_o[26] & L92ov6));
assign Bexiw6 = (~(vis_r6_o[26] & S92ov6));
assign Ndxiw6 = (Pexiw6 & Wexiw6);
assign Wexiw6 = (~(vis_r5_o[26] & Na2ov6));
assign Pexiw6 = (~(vis_r4_o[26] & Ua2ov6));
assign Zcxiw6 = (Dfxiw6 & Kfxiw6);
assign Kfxiw6 = (Rfxiw6 & Yfxiw6);
assign Yfxiw6 = (~(vis_r3_o[26] & Dc2ov6));
assign Rfxiw6 = (~(vis_r2_o[26] & Kc2ov6));
assign Dfxiw6 = (Fgxiw6 & Mgxiw6);
assign Mgxiw6 = (~(vis_r1_o[26] & Fd2ov6));
assign Fgxiw6 = (~(vis_r0_o[26] & Md2ov6));
assign D8xiw6 = (~(H02ov6 & Qw97z6));
assign U6xiw6 = (Tgxiw6 & Ahxiw6);
assign Ahxiw6 = (~(Ve2ov6 & vis_pc_o[26]));
assign Tgxiw6 = (~(Fhc7z6[26] & Cf2ov6));
assign P738v6 = (~(Hhxiw6 & Ohxiw6));
assign Ohxiw6 = (Vhxiw6 & Cixiw6);
assign Cixiw6 = (~(H02ov6 & Yw97z6));
assign Vhxiw6 = (Jixiw6 & Qixiw6);
assign Qixiw6 = (C12ov6 | W8knv6);
assign W8knv6 = (Xixiw6 & Ejxiw6);
assign Ejxiw6 = (Ljxiw6 & Sjxiw6);
assign Sjxiw6 = (Zjxiw6 & Gkxiw6);
assign Gkxiw6 = (Nkxiw6 & Ukxiw6);
assign Ukxiw6 = (~(vis_psp_o[18] & N32ov6));
assign Nkxiw6 = (~(U32ov6 & Pic7z6[18]));
assign Zjxiw6 = (Blxiw6 & Ilxiw6);
assign Ilxiw6 = (~(vis_msp_o[18] & P42ov6));
assign Blxiw6 = (~(vis_r12_o[18] & W42ov6));
assign Ljxiw6 = (Plxiw6 & Wlxiw6);
assign Wlxiw6 = (Dmxiw6 & Kmxiw6);
assign Kmxiw6 = (~(vis_r11_o[18] & F62ov6));
assign Dmxiw6 = (~(vis_r10_o[18] & M62ov6));
assign Plxiw6 = (Rmxiw6 & Ymxiw6);
assign Ymxiw6 = (~(vis_r9_o[18] & H72ov6));
assign Rmxiw6 = (~(vis_r8_o[18] & O72ov6));
assign Xixiw6 = (Fnxiw6 & Mnxiw6);
assign Mnxiw6 = (Tnxiw6 & Aoxiw6);
assign Aoxiw6 = (Hoxiw6 & Ooxiw6);
assign Ooxiw6 = (~(vis_r7_o[18] & L92ov6));
assign Hoxiw6 = (~(vis_r6_o[18] & S92ov6));
assign Tnxiw6 = (Voxiw6 & Cpxiw6);
assign Cpxiw6 = (~(vis_r5_o[18] & Na2ov6));
assign Voxiw6 = (~(vis_r4_o[18] & Ua2ov6));
assign Fnxiw6 = (Jpxiw6 & Qpxiw6);
assign Qpxiw6 = (Xpxiw6 & Eqxiw6);
assign Eqxiw6 = (~(vis_r3_o[18] & Dc2ov6));
assign Xpxiw6 = (~(vis_r2_o[18] & Kc2ov6));
assign Jpxiw6 = (Lqxiw6 & Sqxiw6);
assign Sqxiw6 = (~(vis_r1_o[18] & Fd2ov6));
assign Lqxiw6 = (~(vis_r0_o[18] & Md2ov6));
assign Jixiw6 = (~(Td2ov6 & Zqxiw6));
assign Hhxiw6 = (Grxiw6 & Nrxiw6);
assign Nrxiw6 = (~(Ve2ov6 & vis_pc_o[18]));
assign Grxiw6 = (~(Fhc7z6[18] & Cf2ov6));
assign I738v6 = (~(Urxiw6 & Bsxiw6));
assign Bsxiw6 = (Isxiw6 & Psxiw6);
assign Psxiw6 = (~(H02ov6 & Gx97z6));
assign Isxiw6 = (Wsxiw6 & Dtxiw6);
assign Dtxiw6 = (~(Ktxiw6 & Imknv6));
assign Imknv6 = (~(Rtxiw6 & Ytxiw6));
assign Ytxiw6 = (Fuxiw6 & Muxiw6);
assign Muxiw6 = (Tuxiw6 & Avxiw6);
assign Avxiw6 = (Hvxiw6 & Ovxiw6);
assign Ovxiw6 = (~(vis_psp_o[10] & N32ov6));
assign Hvxiw6 = (~(U32ov6 & Pic7z6[10]));
assign Tuxiw6 = (Vvxiw6 & Cwxiw6);
assign Cwxiw6 = (~(vis_msp_o[10] & P42ov6));
assign Vvxiw6 = (~(vis_r12_o[10] & W42ov6));
assign Fuxiw6 = (Jwxiw6 & Qwxiw6);
assign Qwxiw6 = (Xwxiw6 & Exxiw6);
assign Exxiw6 = (~(vis_r11_o[10] & F62ov6));
assign Xwxiw6 = (~(vis_r10_o[10] & M62ov6));
assign Jwxiw6 = (Lxxiw6 & Sxxiw6);
assign Sxxiw6 = (~(vis_r9_o[10] & H72ov6));
assign Lxxiw6 = (~(vis_r8_o[10] & O72ov6));
assign Rtxiw6 = (Zxxiw6 & Gyxiw6);
assign Gyxiw6 = (Nyxiw6 & Uyxiw6);
assign Uyxiw6 = (Bzxiw6 & Izxiw6);
assign Izxiw6 = (~(vis_r7_o[10] & L92ov6));
assign Bzxiw6 = (~(vis_r6_o[10] & S92ov6));
assign Nyxiw6 = (Pzxiw6 & Wzxiw6);
assign Wzxiw6 = (~(vis_r5_o[10] & Na2ov6));
assign Pzxiw6 = (~(vis_r4_o[10] & Ua2ov6));
assign Zxxiw6 = (D0yiw6 & K0yiw6);
assign K0yiw6 = (R0yiw6 & Y0yiw6);
assign Y0yiw6 = (~(vis_r3_o[10] & Dc2ov6));
assign R0yiw6 = (~(vis_r2_o[10] & Kc2ov6));
assign D0yiw6 = (F1yiw6 & M1yiw6);
assign M1yiw6 = (~(vis_r1_o[10] & Fd2ov6));
assign F1yiw6 = (~(vis_r0_o[10] & Md2ov6));
assign Wsxiw6 = (~(Td2ov6 & T1yiw6));
assign Urxiw6 = (A2yiw6 & H2yiw6);
assign H2yiw6 = (~(Ve2ov6 & vis_pc_o[10]));
assign A2yiw6 = (~(Fhc7z6[10] & Cf2ov6));
assign B738v6 = (~(O2yiw6 & V2yiw6));
assign V2yiw6 = (~(Eji7z6[2] & C3yiw6));
assign O2yiw6 = (J3yiw6 & Q3yiw6);
assign Q3yiw6 = (~(Bhi7z6[2] & X3yiw6));
assign J3yiw6 = (~(E4yiw6 & vis_pc_o[2]));
assign U638v6 = (~(L4yiw6 & S4yiw6));
assign S4yiw6 = (Z4yiw6 & G5yiw6);
assign G5yiw6 = (Eu9ov6 | N5yiw6);
assign Z4yiw6 = (U5yiw6 & B6yiw6);
assign B6yiw6 = (~(Gv9ov6 & Bskov6));
assign U5yiw6 = (~(Uv9ov6 & As97z6));
assign L4yiw6 = (I6yiw6 & P6yiw6);
assign P6yiw6 = (~(Pw9ov6 & Kxb7z6[2]));
assign I6yiw6 = (W6yiw6 & D7yiw6);
assign D7yiw6 = (~(Kx9ov6 & vis_pc_o[2]));
assign W6yiw6 = (~(Gli7z6[2] & Rx9ov6));
assign N638v6 = (K7yiw6 ? vis_psp_o[2] : Bskov6);
assign G638v6 = (K7yiw6 ? vis_psp_o[31] : Ae2ov6);
assign Z538v6 = (K7yiw6 ? vis_psp_o[30] : Fi4ov6);
assign S538v6 = (K7yiw6 ? vis_psp_o[29] : Slbov6);
assign L538v6 = (K7yiw6 ? vis_psp_o[28] : C7aov6);
assign E538v6 = (K7yiw6 ? vis_psp_o[27] : S2gov6);
assign X438v6 = (K7yiw6 ? vis_psp_o[26] : W7xiw6);
assign Q438v6 = (K7yiw6 ? vis_psp_o[25] : R7yiw6);
assign J438v6 = (K7yiw6 ? vis_psp_o[24] : Y7yiw6);
assign C438v6 = (K7yiw6 ? vis_psp_o[23] : F8yiw6);
assign V338v6 = (K7yiw6 ? vis_psp_o[22] : M8yiw6);
assign O338v6 = (K7yiw6 ? vis_psp_o[21] : T8yiw6);
assign H338v6 = (K7yiw6 ? vis_psp_o[20] : A9yiw6);
assign A338v6 = (K7yiw6 ? vis_psp_o[19] : H9yiw6);
assign T238v6 = (K7yiw6 ? vis_psp_o[18] : Zqxiw6);
assign M238v6 = (K7yiw6 ? vis_psp_o[17] : O9yiw6);
assign F238v6 = (K7yiw6 ? vis_psp_o[16] : V9yiw6);
assign Y138v6 = (K7yiw6 ? vis_psp_o[15] : Qccov6);
assign R138v6 = (K7yiw6 ? vis_psp_o[14] : Cayiw6);
assign K138v6 = (K7yiw6 ? vis_psp_o[13] : Jayiw6);
assign D138v6 = (K7yiw6 ? vis_psp_o[12] : Qayiw6);
assign W038v6 = (K7yiw6 ? vis_psp_o[11] : Xayiw6);
assign P038v6 = (K7yiw6 ? vis_psp_o[10] : T1yiw6);
assign K7yiw6 = (!Ebyiw6);
assign I038v6 = (Ebyiw6 ? Lbyiw6 : vis_psp_o[9]);
assign B038v6 = (Ebyiw6 ? W7kov6 : vis_psp_o[8]);
assign Uz28v6 = (Ebyiw6 ? Sbyiw6 : vis_psp_o[7]);
assign Nz28v6 = (Ebyiw6 ? Zbyiw6 : vis_psp_o[6]);
assign Gz28v6 = (Ebyiw6 ? Gcyiw6 : vis_psp_o[5]);
assign Zy28v6 = (Ebyiw6 ? W6lov6 : vis_psp_o[4]);
assign Sy28v6 = (Ebyiw6 ? Ncyiw6 : vis_psp_o[3]);
assign Ebyiw6 = (Ucyiw6 & Bdyiw6);
assign Ly28v6 = (Idyiw6 ? Pic7z6[0] : B2bov6);
assign Ey28v6 = (Idyiw6 ? Pic7z6[31] : Ae2ov6);
assign Xx28v6 = (Idyiw6 ? Pic7z6[30] : Fi4ov6);
assign Qx28v6 = (Idyiw6 ? Pic7z6[29] : Slbov6);
assign Jx28v6 = (Idyiw6 ? Pic7z6[28] : C7aov6);
assign Cx28v6 = (Idyiw6 ? Pic7z6[27] : S2gov6);
assign Vw28v6 = (Idyiw6 ? Pic7z6[26] : W7xiw6);
assign Ow28v6 = (Idyiw6 ? Pic7z6[25] : R7yiw6);
assign Hw28v6 = (Idyiw6 ? Pic7z6[24] : Y7yiw6);
assign Aw28v6 = (Idyiw6 ? Pic7z6[23] : F8yiw6);
assign Tv28v6 = (Idyiw6 ? Pic7z6[22] : M8yiw6);
assign Mv28v6 = (Idyiw6 ? Pic7z6[21] : T8yiw6);
assign Fv28v6 = (Idyiw6 ? Pic7z6[20] : A9yiw6);
assign Yu28v6 = (Idyiw6 ? Pic7z6[19] : H9yiw6);
assign Ru28v6 = (Idyiw6 ? Pic7z6[18] : Zqxiw6);
assign Ku28v6 = (Idyiw6 ? Pic7z6[17] : O9yiw6);
assign Du28v6 = (Idyiw6 ? Pic7z6[16] : V9yiw6);
assign Wt28v6 = (Idyiw6 ? Pic7z6[15] : Qccov6);
assign Pt28v6 = (Idyiw6 ? Pic7z6[14] : Cayiw6);
assign It28v6 = (Idyiw6 ? Pic7z6[13] : Jayiw6);
assign Bt28v6 = (Idyiw6 ? Pic7z6[12] : Qayiw6);
assign Us28v6 = (Idyiw6 ? Pic7z6[11] : Xayiw6);
assign Ns28v6 = (Idyiw6 ? Pic7z6[10] : T1yiw6);
assign Gs28v6 = (Idyiw6 ? Pic7z6[9] : Lbyiw6);
assign Zr28v6 = (Idyiw6 ? Pic7z6[8] : W7kov6);
assign Idyiw6 = (!Pdyiw6);
assign Sr28v6 = (Pdyiw6 ? Sbyiw6 : Pic7z6[7]);
assign Lr28v6 = (Pdyiw6 ? Zbyiw6 : Pic7z6[6]);
assign Er28v6 = (Pdyiw6 ? Gcyiw6 : Pic7z6[5]);
assign Xq28v6 = (Pdyiw6 ? W6lov6 : Pic7z6[4]);
assign Qq28v6 = (Pdyiw6 ? Ncyiw6 : Pic7z6[3]);
assign Jq28v6 = (Pdyiw6 ? Bskov6 : Pic7z6[2]);
assign Cq28v6 = (Pdyiw6 ? Nv9ov6 : Pic7z6[1]);
assign Pdyiw6 = (Ucyiw6 & Wdyiw6);
assign Vp28v6 = (Deyiw6 ? vis_msp_o[2] : Bskov6);
assign Op28v6 = (Deyiw6 ? vis_msp_o[31] : Ae2ov6);
assign Hp28v6 = (Deyiw6 ? vis_msp_o[30] : Fi4ov6);
assign Ap28v6 = (Deyiw6 ? vis_msp_o[29] : Slbov6);
assign To28v6 = (Deyiw6 ? vis_msp_o[28] : C7aov6);
assign Mo28v6 = (Deyiw6 ? vis_msp_o[27] : S2gov6);
assign Fo28v6 = (Deyiw6 ? vis_msp_o[26] : W7xiw6);
assign Yn28v6 = (Deyiw6 ? vis_msp_o[25] : R7yiw6);
assign Rn28v6 = (Deyiw6 ? vis_msp_o[24] : Y7yiw6);
assign Kn28v6 = (Deyiw6 ? vis_msp_o[23] : F8yiw6);
assign Dn28v6 = (Deyiw6 ? vis_msp_o[22] : M8yiw6);
assign Wm28v6 = (Deyiw6 ? vis_msp_o[21] : T8yiw6);
assign Pm28v6 = (Deyiw6 ? vis_msp_o[20] : A9yiw6);
assign Im28v6 = (Deyiw6 ? vis_msp_o[19] : H9yiw6);
assign Bm28v6 = (Deyiw6 ? vis_msp_o[18] : Zqxiw6);
assign Ul28v6 = (Deyiw6 ? vis_msp_o[17] : O9yiw6);
assign Nl28v6 = (Deyiw6 ? vis_msp_o[16] : V9yiw6);
assign Gl28v6 = (Deyiw6 ? vis_msp_o[15] : Qccov6);
assign Zk28v6 = (Deyiw6 ? vis_msp_o[14] : Cayiw6);
assign Sk28v6 = (Deyiw6 ? vis_msp_o[13] : Jayiw6);
assign Lk28v6 = (Deyiw6 ? vis_msp_o[12] : Qayiw6);
assign Ek28v6 = (Deyiw6 ? vis_msp_o[11] : Xayiw6);
assign Xj28v6 = (Deyiw6 ? vis_msp_o[10] : T1yiw6);
assign Qj28v6 = (Deyiw6 ? vis_msp_o[9] : Lbyiw6);
assign Jj28v6 = (Deyiw6 ? vis_msp_o[8] : W7kov6);
assign Cj28v6 = (Deyiw6 ? vis_msp_o[7] : Sbyiw6);
assign Deyiw6 = (!Keyiw6);
assign Vi28v6 = (Keyiw6 ? Zbyiw6 : vis_msp_o[6]);
assign Oi28v6 = (Keyiw6 ? Gcyiw6 : vis_msp_o[5]);
assign Hi28v6 = (Keyiw6 ? W6lov6 : vis_msp_o[4]);
assign Ai28v6 = (Keyiw6 ? Ncyiw6 : vis_msp_o[3]);
assign Keyiw6 = (~(Reyiw6 | Yeyiw6));
assign Th28v6 = (Ffyiw6 ? vis_r12_o[0] : B2bov6);
assign Mh28v6 = (Ffyiw6 ? vis_r12_o[31] : Ae2ov6);
assign Fh28v6 = (Ffyiw6 ? vis_r12_o[30] : Fi4ov6);
assign Yg28v6 = (Ffyiw6 ? vis_r12_o[29] : Slbov6);
assign Rg28v6 = (Ffyiw6 ? vis_r12_o[28] : C7aov6);
assign Kg28v6 = (Ffyiw6 ? vis_r12_o[27] : S2gov6);
assign Dg28v6 = (Ffyiw6 ? vis_r12_o[26] : W7xiw6);
assign Wf28v6 = (Ffyiw6 ? vis_r12_o[25] : R7yiw6);
assign Pf28v6 = (Ffyiw6 ? vis_r12_o[24] : Y7yiw6);
assign If28v6 = (Ffyiw6 ? vis_r12_o[23] : F8yiw6);
assign Bf28v6 = (Ffyiw6 ? vis_r12_o[22] : M8yiw6);
assign Ue28v6 = (Ffyiw6 ? vis_r12_o[21] : T8yiw6);
assign Ne28v6 = (Ffyiw6 ? vis_r12_o[20] : A9yiw6);
assign Ge28v6 = (Ffyiw6 ? vis_r12_o[19] : H9yiw6);
assign Zd28v6 = (Ffyiw6 ? vis_r12_o[18] : Zqxiw6);
assign Sd28v6 = (Ffyiw6 ? vis_r12_o[17] : O9yiw6);
assign Ld28v6 = (Ffyiw6 ? vis_r12_o[16] : V9yiw6);
assign Ed28v6 = (Ffyiw6 ? vis_r12_o[15] : Qccov6);
assign Xc28v6 = (Ffyiw6 ? vis_r12_o[14] : Cayiw6);
assign Qc28v6 = (Ffyiw6 ? vis_r12_o[13] : Jayiw6);
assign Jc28v6 = (Ffyiw6 ? vis_r12_o[12] : Qayiw6);
assign Cc28v6 = (Ffyiw6 ? vis_r12_o[11] : Xayiw6);
assign Vb28v6 = (Ffyiw6 ? vis_r12_o[10] : T1yiw6);
assign Ob28v6 = (Ffyiw6 ? vis_r12_o[9] : Lbyiw6);
assign Hb28v6 = (Ffyiw6 ? vis_r12_o[8] : W7kov6);
assign Ab28v6 = (Ffyiw6 ? vis_r12_o[7] : Sbyiw6);
assign Ta28v6 = (Ffyiw6 ? vis_r12_o[6] : Zbyiw6);
assign Ma28v6 = (Ffyiw6 ? vis_r12_o[5] : Gcyiw6);
assign Ffyiw6 = (!Mfyiw6);
assign Fa28v6 = (Mfyiw6 ? W6lov6 : vis_r12_o[4]);
assign Y928v6 = (Mfyiw6 ? Ncyiw6 : vis_r12_o[3]);
assign R928v6 = (Mfyiw6 ? Bskov6 : vis_r12_o[2]);
assign K928v6 = (Mfyiw6 ? Nv9ov6 : vis_r12_o[1]);
assign Mfyiw6 = (~(Reyiw6 | Tfyiw6));
assign D928v6 = (Agyiw6 ? vis_r11_o[0] : B2bov6);
assign W828v6 = (Agyiw6 ? vis_r11_o[31] : Ae2ov6);
assign P828v6 = (Agyiw6 ? vis_r11_o[30] : Fi4ov6);
assign I828v6 = (Agyiw6 ? vis_r11_o[29] : Slbov6);
assign B828v6 = (Agyiw6 ? vis_r11_o[28] : C7aov6);
assign U728v6 = (Agyiw6 ? vis_r11_o[27] : S2gov6);
assign N728v6 = (Agyiw6 ? vis_r11_o[26] : W7xiw6);
assign G728v6 = (Agyiw6 ? vis_r11_o[25] : R7yiw6);
assign Z628v6 = (Agyiw6 ? vis_r11_o[24] : Y7yiw6);
assign S628v6 = (Agyiw6 ? vis_r11_o[23] : F8yiw6);
assign L628v6 = (Agyiw6 ? vis_r11_o[22] : M8yiw6);
assign E628v6 = (Agyiw6 ? vis_r11_o[21] : T8yiw6);
assign X528v6 = (Agyiw6 ? vis_r11_o[20] : A9yiw6);
assign Q528v6 = (Agyiw6 ? vis_r11_o[19] : H9yiw6);
assign J528v6 = (Agyiw6 ? vis_r11_o[18] : Zqxiw6);
assign C528v6 = (Agyiw6 ? vis_r11_o[17] : O9yiw6);
assign V428v6 = (Agyiw6 ? vis_r11_o[16] : V9yiw6);
assign O428v6 = (Agyiw6 ? vis_r11_o[15] : Qccov6);
assign H428v6 = (Agyiw6 ? vis_r11_o[14] : Cayiw6);
assign A428v6 = (Agyiw6 ? vis_r11_o[13] : Jayiw6);
assign T328v6 = (Agyiw6 ? vis_r11_o[12] : Qayiw6);
assign M328v6 = (Agyiw6 ? vis_r11_o[11] : Xayiw6);
assign F328v6 = (Agyiw6 ? vis_r11_o[10] : T1yiw6);
assign Y228v6 = (Agyiw6 ? vis_r11_o[9] : Lbyiw6);
assign R228v6 = (Agyiw6 ? vis_r11_o[8] : W7kov6);
assign Agyiw6 = (!Hgyiw6);
assign K228v6 = (Hgyiw6 ? Sbyiw6 : vis_r11_o[7]);
assign D228v6 = (Hgyiw6 ? Zbyiw6 : vis_r11_o[6]);
assign W128v6 = (Hgyiw6 ? Gcyiw6 : vis_r11_o[5]);
assign P128v6 = (Hgyiw6 ? W6lov6 : vis_r11_o[4]);
assign I128v6 = (Hgyiw6 ? Ncyiw6 : vis_r11_o[3]);
assign B128v6 = (Hgyiw6 ? Bskov6 : vis_r11_o[2]);
assign U028v6 = (Hgyiw6 ? Nv9ov6 : vis_r11_o[1]);
assign Hgyiw6 = (Ogyiw6 & Bdyiw6);
assign Bdyiw6 = (!Yeyiw6);
assign N028v6 = (Vgyiw6 ? vis_r10_o[0] : B2bov6);
assign G028v6 = (Vgyiw6 ? vis_r10_o[31] : Ae2ov6);
assign Zz18v6 = (Vgyiw6 ? vis_r10_o[30] : Fi4ov6);
assign Sz18v6 = (Vgyiw6 ? vis_r10_o[29] : Slbov6);
assign Lz18v6 = (Vgyiw6 ? vis_r10_o[28] : C7aov6);
assign Ez18v6 = (Vgyiw6 ? vis_r10_o[27] : S2gov6);
assign Xy18v6 = (Vgyiw6 ? vis_r10_o[26] : W7xiw6);
assign Qy18v6 = (Vgyiw6 ? vis_r10_o[25] : R7yiw6);
assign Jy18v6 = (Vgyiw6 ? vis_r10_o[24] : Y7yiw6);
assign Cy18v6 = (Vgyiw6 ? vis_r10_o[23] : F8yiw6);
assign Vx18v6 = (Vgyiw6 ? vis_r10_o[22] : M8yiw6);
assign Ox18v6 = (Vgyiw6 ? vis_r10_o[21] : T8yiw6);
assign Hx18v6 = (Vgyiw6 ? vis_r10_o[20] : A9yiw6);
assign Ax18v6 = (Vgyiw6 ? vis_r10_o[19] : H9yiw6);
assign Tw18v6 = (Vgyiw6 ? vis_r10_o[18] : Zqxiw6);
assign Mw18v6 = (Vgyiw6 ? vis_r10_o[17] : O9yiw6);
assign Fw18v6 = (Vgyiw6 ? vis_r10_o[16] : V9yiw6);
assign Yv18v6 = (Vgyiw6 ? vis_r10_o[15] : Qccov6);
assign Rv18v6 = (Vgyiw6 ? vis_r10_o[14] : Cayiw6);
assign Kv18v6 = (Vgyiw6 ? vis_r10_o[13] : Jayiw6);
assign Dv18v6 = (Vgyiw6 ? vis_r10_o[12] : Qayiw6);
assign Wu18v6 = (Vgyiw6 ? vis_r10_o[11] : Xayiw6);
assign Pu18v6 = (Vgyiw6 ? vis_r10_o[10] : T1yiw6);
assign Iu18v6 = (Vgyiw6 ? vis_r10_o[9] : Lbyiw6);
assign Bu18v6 = (Vgyiw6 ? vis_r10_o[8] : W7kov6);
assign Vgyiw6 = (!Chyiw6);
assign Ut18v6 = (Chyiw6 ? Sbyiw6 : vis_r10_o[7]);
assign Nt18v6 = (Chyiw6 ? Zbyiw6 : vis_r10_o[6]);
assign Gt18v6 = (Chyiw6 ? Gcyiw6 : vis_r10_o[5]);
assign Zs18v6 = (Chyiw6 ? W6lov6 : vis_r10_o[4]);
assign Ss18v6 = (Chyiw6 ? Ncyiw6 : vis_r10_o[3]);
assign Ls18v6 = (Chyiw6 ? Bskov6 : vis_r10_o[2]);
assign Es18v6 = (Chyiw6 ? Nv9ov6 : vis_r10_o[1]);
assign Chyiw6 = (Ogyiw6 & Wdyiw6);
assign Wdyiw6 = (!Tfyiw6);
assign Xr18v6 = (Jhyiw6 ? vis_r9_o[0] : B2bov6);
assign Qr18v6 = (Jhyiw6 ? vis_r9_o[31] : Ae2ov6);
assign Jr18v6 = (Jhyiw6 ? vis_r9_o[30] : Fi4ov6);
assign Cr18v6 = (Jhyiw6 ? vis_r9_o[29] : Slbov6);
assign Vq18v6 = (Jhyiw6 ? vis_r9_o[28] : C7aov6);
assign Oq18v6 = (Jhyiw6 ? vis_r9_o[27] : S2gov6);
assign Hq18v6 = (Jhyiw6 ? vis_r9_o[26] : W7xiw6);
assign Aq18v6 = (Jhyiw6 ? vis_r9_o[25] : R7yiw6);
assign Tp18v6 = (Jhyiw6 ? vis_r9_o[24] : Y7yiw6);
assign Mp18v6 = (Jhyiw6 ? vis_r9_o[23] : F8yiw6);
assign Fp18v6 = (Jhyiw6 ? vis_r9_o[22] : M8yiw6);
assign Yo18v6 = (Jhyiw6 ? vis_r9_o[21] : T8yiw6);
assign Ro18v6 = (Jhyiw6 ? vis_r9_o[20] : A9yiw6);
assign Ko18v6 = (Jhyiw6 ? vis_r9_o[19] : H9yiw6);
assign Do18v6 = (Jhyiw6 ? vis_r9_o[18] : Zqxiw6);
assign Wn18v6 = (Jhyiw6 ? vis_r9_o[17] : O9yiw6);
assign Pn18v6 = (Jhyiw6 ? vis_r9_o[16] : V9yiw6);
assign In18v6 = (Jhyiw6 ? vis_r9_o[15] : Qccov6);
assign Bn18v6 = (Jhyiw6 ? vis_r9_o[14] : Cayiw6);
assign Um18v6 = (Jhyiw6 ? vis_r9_o[13] : Jayiw6);
assign Nm18v6 = (Jhyiw6 ? vis_r9_o[12] : Qayiw6);
assign Gm18v6 = (Jhyiw6 ? vis_r9_o[11] : Xayiw6);
assign Zl18v6 = (Jhyiw6 ? vis_r9_o[10] : T1yiw6);
assign Sl18v6 = (Jhyiw6 ? vis_r9_o[9] : Lbyiw6);
assign Ll18v6 = (Jhyiw6 ? vis_r9_o[8] : W7kov6);
assign El18v6 = (Jhyiw6 ? vis_r9_o[7] : Sbyiw6);
assign Jhyiw6 = (!Qhyiw6);
assign Xk18v6 = (Qhyiw6 ? Zbyiw6 : vis_r9_o[6]);
assign Qk18v6 = (Qhyiw6 ? Gcyiw6 : vis_r9_o[5]);
assign Jk18v6 = (Qhyiw6 ? W6lov6 : vis_r9_o[4]);
assign Ck18v6 = (Qhyiw6 ? Ncyiw6 : vis_r9_o[3]);
assign Vj18v6 = (Qhyiw6 ? Bskov6 : vis_r9_o[2]);
assign Oj18v6 = (Qhyiw6 ? Nv9ov6 : vis_r9_o[1]);
assign Qhyiw6 = (~(Yeyiw6 | Xhyiw6));
assign Yeyiw6 = (~(Eiyiw6 & Liyiw6));
assign Eiyiw6 = (Siyiw6 & Ziyiw6);
assign Hj18v6 = (Gjyiw6 ? vis_r8_o[0] : B2bov6);
assign Aj18v6 = (Gjyiw6 ? vis_r8_o[31] : Ae2ov6);
assign Ti18v6 = (Gjyiw6 ? vis_r8_o[30] : Fi4ov6);
assign Mi18v6 = (Gjyiw6 ? vis_r8_o[29] : Slbov6);
assign Fi18v6 = (Gjyiw6 ? vis_r8_o[28] : C7aov6);
assign Yh18v6 = (Gjyiw6 ? vis_r8_o[27] : S2gov6);
assign Rh18v6 = (Gjyiw6 ? vis_r8_o[26] : W7xiw6);
assign Kh18v6 = (Gjyiw6 ? vis_r8_o[25] : R7yiw6);
assign Dh18v6 = (Gjyiw6 ? vis_r8_o[24] : Y7yiw6);
assign Wg18v6 = (Gjyiw6 ? vis_r8_o[23] : F8yiw6);
assign Pg18v6 = (Gjyiw6 ? vis_r8_o[22] : M8yiw6);
assign Ig18v6 = (Gjyiw6 ? vis_r8_o[21] : T8yiw6);
assign Bg18v6 = (Gjyiw6 ? vis_r8_o[20] : A9yiw6);
assign Uf18v6 = (Gjyiw6 ? vis_r8_o[19] : H9yiw6);
assign Nf18v6 = (Gjyiw6 ? vis_r8_o[18] : Zqxiw6);
assign Gf18v6 = (Gjyiw6 ? vis_r8_o[17] : O9yiw6);
assign Ze18v6 = (Gjyiw6 ? vis_r8_o[16] : V9yiw6);
assign Se18v6 = (Gjyiw6 ? vis_r8_o[15] : Qccov6);
assign Le18v6 = (Gjyiw6 ? vis_r8_o[14] : Cayiw6);
assign Ee18v6 = (Gjyiw6 ? vis_r8_o[13] : Jayiw6);
assign Xd18v6 = (Gjyiw6 ? vis_r8_o[12] : Qayiw6);
assign Qd18v6 = (Gjyiw6 ? vis_r8_o[11] : Xayiw6);
assign Jd18v6 = (Gjyiw6 ? vis_r8_o[10] : T1yiw6);
assign Cd18v6 = (Gjyiw6 ? vis_r8_o[9] : Lbyiw6);
assign Vc18v6 = (Gjyiw6 ? vis_r8_o[8] : W7kov6);
assign Oc18v6 = (Gjyiw6 ? vis_r8_o[7] : Sbyiw6);
assign Gjyiw6 = (!Njyiw6);
assign Hc18v6 = (Njyiw6 ? Zbyiw6 : vis_r8_o[6]);
assign Ac18v6 = (Njyiw6 ? Gcyiw6 : vis_r8_o[5]);
assign Tb18v6 = (Njyiw6 ? W6lov6 : vis_r8_o[4]);
assign Mb18v6 = (Njyiw6 ? Ncyiw6 : vis_r8_o[3]);
assign Fb18v6 = (Njyiw6 ? Bskov6 : vis_r8_o[2]);
assign Ya18v6 = (Njyiw6 ? Nv9ov6 : vis_r8_o[1]);
assign Njyiw6 = (~(Tfyiw6 | Xhyiw6));
assign Tfyiw6 = (~(Ujyiw6 & Liyiw6));
assign Ujyiw6 = (Ziyiw6 & Bkyiw6);
assign Ra18v6 = (Ikyiw6 ? vis_r7_o[0] : B2bov6);
assign Ka18v6 = (Ikyiw6 ? vis_r7_o[31] : Ae2ov6);
assign Da18v6 = (Ikyiw6 ? vis_r7_o[30] : Fi4ov6);
assign W918v6 = (Ikyiw6 ? vis_r7_o[29] : Slbov6);
assign P918v6 = (Ikyiw6 ? vis_r7_o[28] : C7aov6);
assign I918v6 = (Ikyiw6 ? vis_r7_o[27] : S2gov6);
assign B918v6 = (Ikyiw6 ? vis_r7_o[26] : W7xiw6);
assign U818v6 = (Ikyiw6 ? vis_r7_o[25] : R7yiw6);
assign N818v6 = (Ikyiw6 ? vis_r7_o[24] : Y7yiw6);
assign G818v6 = (Ikyiw6 ? vis_r7_o[23] : F8yiw6);
assign Z718v6 = (Ikyiw6 ? vis_r7_o[22] : M8yiw6);
assign S718v6 = (Ikyiw6 ? vis_r7_o[21] : T8yiw6);
assign L718v6 = (Ikyiw6 ? vis_r7_o[20] : A9yiw6);
assign E718v6 = (Ikyiw6 ? vis_r7_o[19] : H9yiw6);
assign X618v6 = (Ikyiw6 ? vis_r7_o[18] : Zqxiw6);
assign Q618v6 = (Ikyiw6 ? vis_r7_o[17] : O9yiw6);
assign J618v6 = (Ikyiw6 ? vis_r7_o[16] : V9yiw6);
assign C618v6 = (Ikyiw6 ? vis_r7_o[15] : Qccov6);
assign V518v6 = (Ikyiw6 ? vis_r7_o[14] : Cayiw6);
assign O518v6 = (Ikyiw6 ? vis_r7_o[13] : Jayiw6);
assign H518v6 = (Ikyiw6 ? vis_r7_o[12] : Qayiw6);
assign A518v6 = (Ikyiw6 ? vis_r7_o[11] : Xayiw6);
assign T418v6 = (Ikyiw6 ? vis_r7_o[10] : T1yiw6);
assign M418v6 = (Ikyiw6 ? vis_r7_o[9] : Lbyiw6);
assign F418v6 = (Ikyiw6 ? vis_r7_o[8] : W7kov6);
assign Ikyiw6 = (!Pkyiw6);
assign Y318v6 = (Pkyiw6 ? Sbyiw6 : vis_r7_o[7]);
assign R318v6 = (Pkyiw6 ? Zbyiw6 : vis_r7_o[6]);
assign K318v6 = (Pkyiw6 ? Gcyiw6 : vis_r7_o[5]);
assign D318v6 = (Pkyiw6 ? W6lov6 : vis_r7_o[4]);
assign W218v6 = (Pkyiw6 ? Ncyiw6 : vis_r7_o[3]);
assign P218v6 = (Pkyiw6 ? Bskov6 : vis_r7_o[2]);
assign I218v6 = (Pkyiw6 ? Nv9ov6 : vis_r7_o[1]);
assign Pkyiw6 = (Ucyiw6 & Wkyiw6);
assign B218v6 = (Dlyiw6 ? vis_r6_o[0] : B2bov6);
assign U118v6 = (Dlyiw6 ? vis_r6_o[31] : Ae2ov6);
assign N118v6 = (Dlyiw6 ? vis_r6_o[30] : Fi4ov6);
assign G118v6 = (Dlyiw6 ? vis_r6_o[29] : Slbov6);
assign Z018v6 = (Dlyiw6 ? vis_r6_o[28] : C7aov6);
assign S018v6 = (Dlyiw6 ? vis_r6_o[27] : S2gov6);
assign L018v6 = (Dlyiw6 ? vis_r6_o[26] : W7xiw6);
assign E018v6 = (Dlyiw6 ? vis_r6_o[25] : R7yiw6);
assign Xz08v6 = (Dlyiw6 ? vis_r6_o[24] : Y7yiw6);
assign Qz08v6 = (Dlyiw6 ? vis_r6_o[23] : F8yiw6);
assign Jz08v6 = (Dlyiw6 ? vis_r6_o[22] : M8yiw6);
assign Cz08v6 = (Dlyiw6 ? vis_r6_o[21] : T8yiw6);
assign Vy08v6 = (Dlyiw6 ? vis_r6_o[20] : A9yiw6);
assign Oy08v6 = (Dlyiw6 ? vis_r6_o[19] : H9yiw6);
assign Hy08v6 = (Dlyiw6 ? vis_r6_o[18] : Zqxiw6);
assign Ay08v6 = (Dlyiw6 ? vis_r6_o[17] : O9yiw6);
assign Tx08v6 = (Dlyiw6 ? vis_r6_o[16] : V9yiw6);
assign Mx08v6 = (Dlyiw6 ? vis_r6_o[15] : Qccov6);
assign Fx08v6 = (Dlyiw6 ? vis_r6_o[14] : Cayiw6);
assign Yw08v6 = (Dlyiw6 ? vis_r6_o[13] : Jayiw6);
assign Rw08v6 = (Dlyiw6 ? vis_r6_o[12] : Qayiw6);
assign Kw08v6 = (Dlyiw6 ? vis_r6_o[11] : Xayiw6);
assign Dw08v6 = (Dlyiw6 ? vis_r6_o[10] : T1yiw6);
assign Wv08v6 = (Dlyiw6 ? vis_r6_o[9] : Lbyiw6);
assign Pv08v6 = (Dlyiw6 ? vis_r6_o[8] : W7kov6);
assign Dlyiw6 = (!Klyiw6);
assign Iv08v6 = (Klyiw6 ? Sbyiw6 : vis_r6_o[7]);
assign Bv08v6 = (Klyiw6 ? Zbyiw6 : vis_r6_o[6]);
assign Uu08v6 = (Klyiw6 ? Gcyiw6 : vis_r6_o[5]);
assign Nu08v6 = (Klyiw6 ? W6lov6 : vis_r6_o[4]);
assign Gu08v6 = (Klyiw6 ? Ncyiw6 : vis_r6_o[3]);
assign Zt08v6 = (Klyiw6 ? Bskov6 : vis_r6_o[2]);
assign St08v6 = (Klyiw6 ? Nv9ov6 : vis_r6_o[1]);
assign Klyiw6 = (Ucyiw6 & Rlyiw6);
assign Ucyiw6 = (Ylyiw6 & Fmyiw6);
assign Lt08v6 = (Mmyiw6 ? vis_r5_o[0] : B2bov6);
assign Et08v6 = (Mmyiw6 ? vis_r5_o[31] : Ae2ov6);
assign Xs08v6 = (Mmyiw6 ? vis_r5_o[30] : Fi4ov6);
assign Qs08v6 = (Mmyiw6 ? vis_r5_o[29] : Slbov6);
assign Js08v6 = (Mmyiw6 ? vis_r5_o[28] : C7aov6);
assign Cs08v6 = (Mmyiw6 ? vis_r5_o[27] : S2gov6);
assign Vr08v6 = (Mmyiw6 ? vis_r5_o[26] : W7xiw6);
assign Or08v6 = (Mmyiw6 ? vis_r5_o[25] : R7yiw6);
assign Hr08v6 = (Mmyiw6 ? vis_r5_o[24] : Y7yiw6);
assign Ar08v6 = (Mmyiw6 ? vis_r5_o[23] : F8yiw6);
assign Tq08v6 = (Mmyiw6 ? vis_r5_o[22] : M8yiw6);
assign Mq08v6 = (Mmyiw6 ? vis_r5_o[21] : T8yiw6);
assign Fq08v6 = (Mmyiw6 ? vis_r5_o[20] : A9yiw6);
assign Yp08v6 = (Mmyiw6 ? vis_r5_o[19] : H9yiw6);
assign Rp08v6 = (Mmyiw6 ? vis_r5_o[18] : Zqxiw6);
assign Kp08v6 = (Mmyiw6 ? vis_r5_o[17] : O9yiw6);
assign Dp08v6 = (Mmyiw6 ? vis_r5_o[16] : V9yiw6);
assign Wo08v6 = (Mmyiw6 ? vis_r5_o[15] : Qccov6);
assign Po08v6 = (Mmyiw6 ? vis_r5_o[14] : Cayiw6);
assign Io08v6 = (Mmyiw6 ? vis_r5_o[13] : Jayiw6);
assign Bo08v6 = (Mmyiw6 ? vis_r5_o[12] : Qayiw6);
assign Un08v6 = (Mmyiw6 ? vis_r5_o[11] : Xayiw6);
assign Nn08v6 = (Mmyiw6 ? vis_r5_o[10] : T1yiw6);
assign Gn08v6 = (Mmyiw6 ? vis_r5_o[9] : Lbyiw6);
assign Zm08v6 = (Mmyiw6 ? vis_r5_o[8] : W7kov6);
assign Sm08v6 = (Mmyiw6 ? vis_r5_o[7] : Sbyiw6);
assign Lm08v6 = (Mmyiw6 ? vis_r5_o[6] : Zbyiw6);
assign Em08v6 = (Mmyiw6 ? vis_r5_o[5] : Gcyiw6);
assign Mmyiw6 = (!Tmyiw6);
assign Xl08v6 = (Tmyiw6 ? W6lov6 : vis_r5_o[4]);
assign Ql08v6 = (Tmyiw6 ? Ncyiw6 : vis_r5_o[3]);
assign Jl08v6 = (Tmyiw6 ? Bskov6 : vis_r5_o[2]);
assign Cl08v6 = (Tmyiw6 ? Nv9ov6 : vis_r5_o[1]);
assign Tmyiw6 = (~(Anyiw6 | Reyiw6));
assign Vk08v6 = (Hnyiw6 ? vis_r4_o[0] : B2bov6);
assign Ok08v6 = (Hnyiw6 ? vis_r4_o[31] : Ae2ov6);
assign Hk08v6 = (Hnyiw6 ? vis_r4_o[30] : Fi4ov6);
assign Ak08v6 = (Hnyiw6 ? vis_r4_o[29] : Slbov6);
assign Tj08v6 = (Hnyiw6 ? vis_r4_o[28] : C7aov6);
assign Mj08v6 = (Hnyiw6 ? vis_r4_o[27] : S2gov6);
assign Fj08v6 = (Hnyiw6 ? vis_r4_o[26] : W7xiw6);
assign Yi08v6 = (Hnyiw6 ? vis_r4_o[25] : R7yiw6);
assign Ri08v6 = (Hnyiw6 ? vis_r4_o[24] : Y7yiw6);
assign Ki08v6 = (Hnyiw6 ? vis_r4_o[23] : F8yiw6);
assign Di08v6 = (Hnyiw6 ? vis_r4_o[22] : M8yiw6);
assign Wh08v6 = (Hnyiw6 ? vis_r4_o[21] : T8yiw6);
assign Ph08v6 = (Hnyiw6 ? vis_r4_o[20] : A9yiw6);
assign Ih08v6 = (Hnyiw6 ? vis_r4_o[19] : H9yiw6);
assign Bh08v6 = (Hnyiw6 ? vis_r4_o[18] : Zqxiw6);
assign Ug08v6 = (Hnyiw6 ? vis_r4_o[17] : O9yiw6);
assign Ng08v6 = (Hnyiw6 ? vis_r4_o[16] : V9yiw6);
assign Gg08v6 = (Hnyiw6 ? vis_r4_o[15] : Qccov6);
assign Zf08v6 = (Hnyiw6 ? vis_r4_o[14] : Cayiw6);
assign Sf08v6 = (Hnyiw6 ? vis_r4_o[13] : Jayiw6);
assign Lf08v6 = (Hnyiw6 ? vis_r4_o[12] : Qayiw6);
assign Ef08v6 = (Hnyiw6 ? vis_r4_o[11] : Xayiw6);
assign Xe08v6 = (Hnyiw6 ? vis_r4_o[10] : T1yiw6);
assign Qe08v6 = (Hnyiw6 ? vis_r4_o[9] : Lbyiw6);
assign Je08v6 = (Hnyiw6 ? vis_r4_o[8] : W7kov6);
assign Hnyiw6 = (!Onyiw6);
assign Ce08v6 = (Onyiw6 ? Sbyiw6 : vis_r4_o[7]);
assign Vd08v6 = (Onyiw6 ? Zbyiw6 : vis_r4_o[6]);
assign Od08v6 = (Onyiw6 ? Gcyiw6 : vis_r4_o[5]);
assign Hd08v6 = (Onyiw6 ? W6lov6 : vis_r4_o[4]);
assign Ad08v6 = (Onyiw6 ? Ncyiw6 : vis_r4_o[3]);
assign Tc08v6 = (Onyiw6 ? Bskov6 : vis_r4_o[2]);
assign Mc08v6 = (Onyiw6 ? Nv9ov6 : vis_r4_o[1]);
assign Onyiw6 = (~(Reyiw6 | Vnyiw6));
assign Reyiw6 = (Ylyiw6 | Coyiw6);
assign Fc08v6 = (Joyiw6 ? vis_r3_o[0] : B2bov6);
assign Yb08v6 = (Joyiw6 ? vis_r3_o[31] : Ae2ov6);
assign Rb08v6 = (Joyiw6 ? vis_r3_o[30] : Fi4ov6);
assign Kb08v6 = (Joyiw6 ? vis_r3_o[29] : Slbov6);
assign Db08v6 = (Joyiw6 ? vis_r3_o[28] : C7aov6);
assign Wa08v6 = (Joyiw6 ? vis_r3_o[27] : S2gov6);
assign Pa08v6 = (Joyiw6 ? vis_r3_o[26] : W7xiw6);
assign Ia08v6 = (Joyiw6 ? vis_r3_o[25] : R7yiw6);
assign Ba08v6 = (Joyiw6 ? vis_r3_o[24] : Y7yiw6);
assign U908v6 = (Joyiw6 ? vis_r3_o[23] : F8yiw6);
assign N908v6 = (Joyiw6 ? vis_r3_o[22] : M8yiw6);
assign G908v6 = (Joyiw6 ? vis_r3_o[21] : T8yiw6);
assign Z808v6 = (Joyiw6 ? vis_r3_o[20] : A9yiw6);
assign S808v6 = (Joyiw6 ? vis_r3_o[19] : H9yiw6);
assign L808v6 = (Joyiw6 ? vis_r3_o[18] : Zqxiw6);
assign E808v6 = (Joyiw6 ? vis_r3_o[17] : O9yiw6);
assign X708v6 = (Joyiw6 ? vis_r3_o[16] : V9yiw6);
assign Q708v6 = (Joyiw6 ? vis_r3_o[15] : Qccov6);
assign J708v6 = (Joyiw6 ? vis_r3_o[14] : Cayiw6);
assign C708v6 = (Joyiw6 ? vis_r3_o[13] : Jayiw6);
assign V608v6 = (Joyiw6 ? vis_r3_o[12] : Qayiw6);
assign O608v6 = (Joyiw6 ? vis_r3_o[11] : Xayiw6);
assign H608v6 = (Joyiw6 ? vis_r3_o[10] : T1yiw6);
assign A608v6 = (Joyiw6 ? vis_r3_o[9] : Lbyiw6);
assign T508v6 = (Joyiw6 ? vis_r3_o[8] : W7kov6);
assign Joyiw6 = (!Qoyiw6);
assign M508v6 = (Qoyiw6 ? Sbyiw6 : vis_r3_o[7]);
assign F508v6 = (Qoyiw6 ? Zbyiw6 : vis_r3_o[6]);
assign Y408v6 = (Qoyiw6 ? Gcyiw6 : vis_r3_o[5]);
assign R408v6 = (Qoyiw6 ? W6lov6 : vis_r3_o[4]);
assign K408v6 = (Qoyiw6 ? Ncyiw6 : vis_r3_o[3]);
assign D408v6 = (Qoyiw6 ? Bskov6 : vis_r3_o[2]);
assign W308v6 = (Qoyiw6 ? Nv9ov6 : vis_r3_o[1]);
assign Qoyiw6 = (Ogyiw6 & Wkyiw6);
assign Wkyiw6 = (!Anyiw6);
assign P308v6 = (Xoyiw6 ? vis_r2_o[0] : B2bov6);
assign I308v6 = (Xoyiw6 ? vis_r2_o[31] : Ae2ov6);
assign B308v6 = (Xoyiw6 ? vis_r2_o[30] : Fi4ov6);
assign U208v6 = (Xoyiw6 ? vis_r2_o[29] : Slbov6);
assign N208v6 = (Xoyiw6 ? vis_r2_o[28] : C7aov6);
assign G208v6 = (Xoyiw6 ? vis_r2_o[27] : S2gov6);
assign Z108v6 = (Xoyiw6 ? vis_r2_o[26] : W7xiw6);
assign S108v6 = (Xoyiw6 ? vis_r2_o[25] : R7yiw6);
assign L108v6 = (Xoyiw6 ? vis_r2_o[24] : Y7yiw6);
assign E108v6 = (Xoyiw6 ? vis_r2_o[23] : F8yiw6);
assign X008v6 = (Xoyiw6 ? vis_r2_o[22] : M8yiw6);
assign Q008v6 = (Xoyiw6 ? vis_r2_o[21] : T8yiw6);
assign J008v6 = (Xoyiw6 ? vis_r2_o[20] : A9yiw6);
assign C008v6 = (Xoyiw6 ? vis_r2_o[19] : H9yiw6);
assign Vzz7v6 = (Xoyiw6 ? vis_r2_o[18] : Zqxiw6);
assign Ozz7v6 = (Xoyiw6 ? vis_r2_o[17] : O9yiw6);
assign Hzz7v6 = (Xoyiw6 ? vis_r2_o[16] : V9yiw6);
assign Azz7v6 = (Xoyiw6 ? vis_r2_o[15] : Qccov6);
assign Tyz7v6 = (Xoyiw6 ? vis_r2_o[14] : Cayiw6);
assign Myz7v6 = (Xoyiw6 ? vis_r2_o[13] : Jayiw6);
assign Fyz7v6 = (Xoyiw6 ? vis_r2_o[12] : Qayiw6);
assign Yxz7v6 = (Xoyiw6 ? vis_r2_o[11] : Xayiw6);
assign Rxz7v6 = (Xoyiw6 ? vis_r2_o[10] : T1yiw6);
assign Kxz7v6 = (Xoyiw6 ? vis_r2_o[9] : Lbyiw6);
assign Dxz7v6 = (Xoyiw6 ? vis_r2_o[8] : W7kov6);
assign Xoyiw6 = (!Epyiw6);
assign Wwz7v6 = (Epyiw6 ? Sbyiw6 : vis_r2_o[7]);
assign Pwz7v6 = (Epyiw6 ? Zbyiw6 : vis_r2_o[6]);
assign Iwz7v6 = (Epyiw6 ? Gcyiw6 : vis_r2_o[5]);
assign Bwz7v6 = (Epyiw6 ? W6lov6 : vis_r2_o[4]);
assign Uvz7v6 = (Epyiw6 ? Ncyiw6 : vis_r2_o[3]);
assign Nvz7v6 = (Epyiw6 ? Bskov6 : vis_r2_o[2]);
assign Gvz7v6 = (Epyiw6 ? Nv9ov6 : vis_r2_o[1]);
assign Epyiw6 = (Ogyiw6 & Rlyiw6);
assign Ogyiw6 = (Coyiw6 & Ylyiw6);
assign Zuz7v6 = (Lpyiw6 ? vis_r1_o[0] : B2bov6);
assign Suz7v6 = (Lpyiw6 ? vis_r1_o[31] : Ae2ov6);
assign Ae2ov6 = (Spyiw6 ? Wt97z6 : Gli7z6[31]);
assign Wt97z6 = (~(Zpyiw6 & Gqyiw6));
assign Gqyiw6 = (~(Nqyiw6 & Bvwnv6));
assign Bvwnv6 = (~(Uqyiw6 & Bryiw6));
assign Bryiw6 = (Iryiw6 & Pryiw6);
assign Pryiw6 = (~(Wryiw6 & Hjjnv6));
assign Iryiw6 = (Dsyiw6 & Ksyiw6);
assign Ksyiw6 = (~(Ju1ov6 & Rsyiw6));
assign Dsyiw6 = (~(Nqh7z6[31] & Ysyiw6));
assign Uqyiw6 = (Ftyiw6 & Mtyiw6);
assign Mtyiw6 = (~(Fth7z6[31] & Ttyiw6));
assign Zpyiw6 = (Auyiw6 & Huyiw6);
assign Huyiw6 = (~(Pdc7z6[31] & Ouyiw6));
assign Auyiw6 = (~(Vuyiw6 & Cvyiw6));
assign Cvyiw6 = (~(Jvyiw6 & Qvyiw6));
assign Qvyiw6 = (Xvyiw6 & Ewyiw6);
assign Ewyiw6 = (Lwyiw6 & Swyiw6);
assign Swyiw6 = (Zwyiw6 & Gxyiw6);
assign Gxyiw6 = (~(Nxyiw6 & Rje7z6[31]));
assign Nxyiw6 = (Uxyiw6 & Kxb7z6[31]);
assign Zwyiw6 = (~(Byyiw6 & Wx1ov6));
assign Byyiw6 = (Dy1ov6 & J1gov6);
assign Lwyiw6 = (Iyyiw6 & Pyyiw6);
assign Pyyiw6 = (~(Wyyiw6 & V5bov6));
assign Wyyiw6 = (~(Dzyiw6 & Kzyiw6));
assign Dzyiw6 = (Rzyiw6 & Yzyiw6);
assign Yzyiw6 = (~(F0ziw6 & M0ziw6));
assign Rzyiw6 = (Ninnv6 | Rje7z6[31]);
assign Iyyiw6 = (~(T0ziw6 & Rje7z6[31]));
assign Xvyiw6 = (A1ziw6 & H1ziw6);
assign H1ziw6 = (~(L0g7z6[15] & O1ziw6));
assign A1ziw6 = (V1ziw6 & C2ziw6);
assign C2ziw6 = (~(L0g7z6[31] & J2ziw6));
assign V1ziw6 = (~(Cqf7z6[15] & Q2ziw6));
assign Jvyiw6 = (X2ziw6 & E3ziw6);
assign E3ziw6 = (L3ziw6 & S3ziw6);
assign S3ziw6 = (~(Z3ziw6 & E3c7z6[0]));
assign L3ziw6 = (G4ziw6 & N4ziw6);
assign N4ziw6 = (~(U4ziw6 & V1c7z6[31]));
assign G4ziw6 = (~(B5ziw6 & O4gdt6));
assign X2ziw6 = (I5ziw6 & Ry1ov6);
assign Ry1ov6 = (P5ziw6 & W5ziw6);
assign W5ziw6 = (D6ziw6 & K6ziw6);
assign K6ziw6 = (~(R6ziw6 & Y6ziw6));
assign D6ziw6 = (~(F7ziw6 & M7ziw6));
assign P5ziw6 = (T7ziw6 & A8ziw6);
assign A8ziw6 = (~(J73ov6 & H8ziw6));
assign I5ziw6 = (Ky1ov6 & O8ziw6);
assign O8ziw6 = (~(Mtkdt6 & Oztiw6));
assign Ky1ov6 = (J9ziw6 ? C9ziw6 : V8ziw6);
assign J9ziw6 = (!N2aov6);
assign N2aov6 = (Q9ziw6 ^ Dte7z6[0]);
assign Q9ziw6 = (~(X9ziw6 & Eaziw6));
assign Eaziw6 = (~(Yxf7z6[15] & Laziw6));
assign X9ziw6 = (Saziw6 & Zaziw6);
assign Zaziw6 = (~(Gbziw6 & Yxf7z6[31]));
assign Saziw6 = (~(Kxb7z6[31] & Nbziw6));
assign C9ziw6 = (~(B3aov6 & Ubziw6));
assign V8ziw6 = (B3aov6 ? Icziw6 : Bcziw6);
assign B3aov6 = (Mennv6 ^ Pcziw6);
assign Pcziw6 = (Wcziw6 & Ddziw6);
assign Ddziw6 = (~(Kdziw6 & Rdziw6));
assign Wcziw6 = (~(Ydziw6 & Feziw6));
assign Feziw6 = (~(Meziw6 & Teziw6));
assign Teziw6 = (Afziw6 & Hfziw6);
assign Hfziw6 = (~(Onf7z6[31] & Ofziw6));
assign Afziw6 = (Vfziw6 & Cgziw6);
assign Cgziw6 = (~(Kxb7z6[31] & Jgziw6));
assign Jgziw6 = (~(Z6jhw6 & Qgziw6));
assign Vfziw6 = (~(Gvtiw6 & Xgziw6));
assign Xgziw6 = (~(Ehziw6 & Lhziw6));
assign Lhziw6 = (Shziw6 & Zhziw6);
assign Zhziw6 = (~(Yxf7z6[31] & Giziw6));
assign Shziw6 = (~(Yxf7z6[32] & Niziw6));
assign Ehziw6 = (Uiziw6 & Bjziw6);
assign Bjziw6 = (~(Yxf7z6[33] & Ijziw6));
assign Uiziw6 = (~(Yxf7z6[34] & Pjziw6));
assign Meziw6 = (Wjziw6 & Dkziw6);
assign Dkziw6 = (Ebmnv6 | Kkziw6);
assign Ebmnv6 = (!Alf7z6[31]);
assign Wjziw6 = (~(Alf7z6[15] & Rkziw6));
assign Luz7v6 = (Lpyiw6 ? vis_r1_o[30] : Fi4ov6);
assign Euz7v6 = (Lpyiw6 ? vis_r1_o[29] : Slbov6);
assign Xtz7v6 = (Lpyiw6 ? vis_r1_o[28] : C7aov6);
assign Qtz7v6 = (Lpyiw6 ? vis_r1_o[27] : S2gov6);
assign Jtz7v6 = (Lpyiw6 ? vis_r1_o[26] : W7xiw6);
assign Ctz7v6 = (Lpyiw6 ? vis_r1_o[25] : R7yiw6);
assign Vsz7v6 = (Lpyiw6 ? vis_r1_o[24] : Y7yiw6);
assign Osz7v6 = (Lpyiw6 ? vis_r1_o[23] : F8yiw6);
assign Hsz7v6 = (Lpyiw6 ? vis_r1_o[22] : M8yiw6);
assign Asz7v6 = (Lpyiw6 ? vis_r1_o[21] : T8yiw6);
assign Trz7v6 = (Lpyiw6 ? vis_r1_o[20] : A9yiw6);
assign Mrz7v6 = (Lpyiw6 ? vis_r1_o[19] : H9yiw6);
assign Frz7v6 = (Lpyiw6 ? vis_r1_o[18] : Zqxiw6);
assign Yqz7v6 = (Lpyiw6 ? vis_r1_o[17] : O9yiw6);
assign Rqz7v6 = (Lpyiw6 ? vis_r1_o[16] : V9yiw6);
assign Kqz7v6 = (Lpyiw6 ? vis_r1_o[15] : Qccov6);
assign Dqz7v6 = (Lpyiw6 ? vis_r1_o[14] : Cayiw6);
assign Wpz7v6 = (Lpyiw6 ? vis_r1_o[13] : Jayiw6);
assign Ppz7v6 = (Lpyiw6 ? vis_r1_o[12] : Qayiw6);
assign Ipz7v6 = (Lpyiw6 ? vis_r1_o[11] : Xayiw6);
assign Bpz7v6 = (Lpyiw6 ? vis_r1_o[10] : T1yiw6);
assign Uoz7v6 = (Lpyiw6 ? vis_r1_o[9] : Lbyiw6);
assign Noz7v6 = (Lpyiw6 ? vis_r1_o[8] : W7kov6);
assign Goz7v6 = (Lpyiw6 ? vis_r1_o[7] : Sbyiw6);
assign Lpyiw6 = (!Ykziw6);
assign Znz7v6 = (Ykziw6 ? Zbyiw6 : vis_r1_o[6]);
assign Snz7v6 = (Ykziw6 ? Gcyiw6 : vis_r1_o[5]);
assign Lnz7v6 = (Ykziw6 ? W6lov6 : vis_r1_o[4]);
assign Enz7v6 = (Ykziw6 ? Ncyiw6 : vis_r1_o[3]);
assign Xmz7v6 = (Ykziw6 ? Bskov6 : vis_r1_o[2]);
assign Qmz7v6 = (Ykziw6 ? Nv9ov6 : vis_r1_o[1]);
assign Ykziw6 = (~(Anyiw6 | Xhyiw6));
assign Anyiw6 = (~(Flziw6 & Liyiw6));
assign Flziw6 = (Mlziw6 & Siyiw6);
assign Jmz7v6 = (Tbbov6 ? vis_r0_o[0] : B2bov6);
assign B2bov6 = (~(Spyiw6 & Tlziw6));
assign Tlziw6 = (~(Gghov6 & Amziw6));
assign Gghov6 = (~(Hmziw6 & Omziw6));
assign Omziw6 = (~(Pdc7z6[0] & Ouyiw6));
assign Hmziw6 = (Vmziw6 & Cnziw6);
assign Cnziw6 = (~(Vuyiw6 & Jnziw6));
assign Jnziw6 = (~(Qnziw6 & Xnziw6));
assign Xnziw6 = (Eoziw6 & Loziw6);
assign Loziw6 = (Soziw6 & Zoziw6);
assign Zoziw6 = (Gpziw6 & Npziw6);
assign Npziw6 = (~(Upziw6 & C1gov6));
assign Upziw6 = (Bqziw6 & Tkbdt6);
assign Gpziw6 = (Iqziw6 & Pqziw6);
assign Pqziw6 = (~(Wqziw6 & Drziw6));
assign Drziw6 = (Krziw6 & Rrziw6);
assign Rrziw6 = (~(Yrziw6 & Fsziw6));
assign Fsziw6 = (~(Dte7z6[14] & Inadt6));
assign Yrziw6 = (~(Dte7z6[13] & Nmadt6));
assign Krziw6 = (N99iw6 & Msziw6);
assign Wqziw6 = (Dte7z6[15] & Dte7z6[16]);
assign Iqziw6 = (~(Tsziw6 & Uxyiw6));
assign Tsziw6 = (Kxb7z6[0] & Atziw6);
assign Soziw6 = (Htziw6 & Otziw6);
assign Otziw6 = (~(Vtziw6 & Cuziw6));
assign Vtziw6 = (~(Juziw6 & Quziw6));
assign Juziw6 = (Xuziw6 & Evziw6);
assign Xuziw6 = (Atziw6 | Ninnv6);
assign Atziw6 = (Lvziw6 | Rje7z6[0]);
assign Htziw6 = (~(Svziw6 & Rknnv6));
assign Rknnv6 = (~(Zvziw6 & Gwziw6));
assign Gwziw6 = (Nwziw6 & Uwziw6);
assign Uwziw6 = (~(Bxziw6 & Ixziw6));
assign Ixziw6 = (~(Pxziw6 & Wxziw6));
assign Wxziw6 = (~(Dyziw6 & Kyziw6));
assign Kyziw6 = (~(Ryziw6 & Yyziw6));
assign Ryziw6 = (Tzziw6 ? Mzziw6 : Fzziw6);
assign Mzziw6 = (~(A00jw6 & H00jw6));
assign A00jw6 = (O00jw6 | V00jw6);
assign V00jw6 = (~(C10jw6 | J10jw6));
assign J10jw6 = (!Q10jw6);
assign Fzziw6 = (H00jw6 | X10jw6);
assign X10jw6 = (O00jw6 & E20jw6);
assign E20jw6 = (~(Q10jw6 & C10jw6));
assign Pxziw6 = (~(L20jw6 & S20jw6));
assign Nwziw6 = (Z20jw6 & G30jw6);
assign G30jw6 = (~(N30jw6 & U30jw6));
assign N30jw6 = (B40jw6 & I40jw6);
assign Z20jw6 = (~(P40jw6 & W40jw6));
assign W40jw6 = (~(D50jw6 & K50jw6));
assign K50jw6 = (~(R50jw6 & Y50jw6));
assign Y50jw6 = (~(F60jw6 & M60jw6));
assign F60jw6 = (Tzziw6 ? A70jw6 : T60jw6);
assign A70jw6 = (~(H70jw6 & O70jw6));
assign H70jw6 = (V70jw6 | C80jw6);
assign C80jw6 = (~(J80jw6 | Q80jw6));
assign Q80jw6 = (!X80jw6);
assign T60jw6 = (O70jw6 | E90jw6);
assign E90jw6 = (V70jw6 & L90jw6);
assign L90jw6 = (~(X80jw6 & J80jw6));
assign D50jw6 = (S90jw6 | Z90jw6);
assign Zvziw6 = (Ga0jw6 & Na0jw6);
assign Na0jw6 = (~(Ua0jw6 & Bb0jw6));
assign Bb0jw6 = (~(Ib0jw6 & Pb0jw6));
assign Pb0jw6 = (~(Wb0jw6 & Dc0jw6));
assign Dc0jw6 = (~(Kc0jw6 & Rc0jw6));
assign Kc0jw6 = (Tzziw6 ? Fd0jw6 : Yc0jw6);
assign Fd0jw6 = (~(Md0jw6 & Td0jw6));
assign Md0jw6 = (Ae0jw6 | He0jw6);
assign He0jw6 = (~(Oe0jw6 | Ve0jw6));
assign Ve0jw6 = (!Cf0jw6);
assign Yc0jw6 = (Td0jw6 | Jf0jw6);
assign Jf0jw6 = (Ae0jw6 & Qf0jw6);
assign Qf0jw6 = (~(Cf0jw6 & Oe0jw6));
assign Ib0jw6 = (Xf0jw6 | Eg0jw6);
assign Ga0jw6 = (~(Lg0jw6 & Sg0jw6));
assign Lg0jw6 = (~(Zg0jw6 & Gh0jw6));
assign Zg0jw6 = (Tzziw6 ? Uh0jw6 : Nh0jw6);
assign Uh0jw6 = (~(Bi0jw6 & Ii0jw6));
assign Bi0jw6 = (Pi0jw6 | Wi0jw6);
assign Wi0jw6 = (Dj0jw6 & Kj0jw6);
assign Nh0jw6 = (Ii0jw6 | Rj0jw6);
assign Rj0jw6 = (Pi0jw6 & Yj0jw6);
assign Yj0jw6 = (Fk0jw6 | Kj0jw6);
assign Eoziw6 = (Mk0jw6 & Tk0jw6);
assign Tk0jw6 = (Al0jw6 & Hl0jw6);
assign Hl0jw6 = (~(Ol0jw6 & Bo3ov6));
assign Al0jw6 = (~(J73ov6 & Pa3ov6));
assign Mk0jw6 = (Vl0jw6 & Cm0jw6);
assign Cm0jw6 = (~(Tj3ov6 & C73ov6));
assign Vl0jw6 = (~(Jm0jw6 & Qm0jw6));
assign Qnziw6 = (Xm0jw6 & En0jw6);
assign En0jw6 = (Ln0jw6 & Sn0jw6);
assign Sn0jw6 = (Zn0jw6 & Go0jw6);
assign Go0jw6 = (~(L0g7z6[0] & J2ziw6));
assign Zn0jw6 = (No0jw6 & Uo0jw6);
assign Uo0jw6 = (~(T0ziw6 & Rje7z6[0]));
assign No0jw6 = (Ryfov6 | Bp0jw6);
assign Ln0jw6 = (Ip0jw6 & Pp0jw6);
assign Pp0jw6 = (~(L0g7z6[16] & Q2ziw6));
assign Ip0jw6 = (~(O1ziw6 & Onf7z6[0]));
assign Xm0jw6 = (Wp0jw6 & Dq0jw6);
assign Dq0jw6 = (Kq0jw6 & Rq0jw6);
assign Rq0jw6 = (~(U4ziw6 & E3c7z6[0]));
assign Kq0jw6 = (~(Z3ziw6 & Fhc7z6[31]));
assign Wp0jw6 = (Dq2ov6 & Yq0jw6);
assign Yq0jw6 = (~(Bnmdt6 & Oztiw6));
assign Dq2ov6 = (Fr0jw6 & Mr0jw6);
assign Mr0jw6 = (~(Tr0jw6 & As0jw6));
assign Tr0jw6 = (~(Hs0jw6 | Icziw6));
assign Hs0jw6 = (!Zannv6);
assign Fr0jw6 = (~(Os0jw6 & Ubziw6));
assign Os0jw6 = (As0jw6 ^ Zannv6);
assign Zannv6 = (~(Vs0jw6 ^ Mennv6));
assign Vs0jw6 = (~(Ct0jw6 & Jt0jw6));
assign Jt0jw6 = (Qt0jw6 & Xt0jw6);
assign Xt0jw6 = (Eu0jw6 & Lu0jw6);
assign Lu0jw6 = (~(Yxf7z6[2] & Su0jw6));
assign Eu0jw6 = (Zu0jw6 & Gv0jw6);
assign Gv0jw6 = (~(Yxf7z6[0] & Nv0jw6));
assign Zu0jw6 = (~(Yxf7z6[1] & Uv0jw6));
assign Qt0jw6 = (Bw0jw6 & Iw0jw6);
assign Iw0jw6 = (~(Yxf7z6[3] & Pw0jw6));
assign Bw0jw6 = (Ww0jw6 | Dx0jw6);
assign Ct0jw6 = (Kx0jw6 & Rx0jw6);
assign Rx0jw6 = (Yx0jw6 & Fy0jw6);
assign Fy0jw6 = (~(Onf7z6[0] & My0jw6));
assign Yx0jw6 = (Ty0jw6 & Az0jw6);
assign Az0jw6 = (~(Hz0jw6 & Kxb7z6[0]));
assign Ty0jw6 = (~(Oz0jw6 & E3c7z6[0]));
assign Kx0jw6 = (Vz0jw6 & C01jw6);
assign C01jw6 = (~(Onf7z6[16] & J01jw6));
assign Vz0jw6 = (~(Alf7z6[0] & Q01jw6));
assign As0jw6 = (!Lannv6);
assign Lannv6 = (X01jw6 ^ Tennv6);
assign X01jw6 = (~(E11jw6 & L11jw6));
assign L11jw6 = (~(Kxb7z6[0] & S11jw6));
assign E11jw6 = (~(Yxf7z6[0] & Gbziw6));
assign Vmziw6 = (Z11jw6 | G21jw6);
assign Cmz7v6 = (Tbbov6 ? vis_r0_o[30] : Fi4ov6);
assign Vlz7v6 = (Tbbov6 ? vis_r0_o[29] : Slbov6);
assign Slbov6 = (Spyiw6 ? Cv97z6 : Gli7z6[29]);
assign Cv97z6 = (~(N21jw6 & U21jw6));
assign U21jw6 = (~(Nqyiw6 & Pgxnv6));
assign N21jw6 = (B31jw6 & I31jw6);
assign I31jw6 = (~(Pdc7z6[29] & Ouyiw6));
assign B31jw6 = (~(Vuyiw6 & P31jw6));
assign P31jw6 = (~(W31jw6 & D41jw6));
assign D41jw6 = (K41jw6 & R41jw6);
assign R41jw6 = (Y41jw6 & F51jw6);
assign F51jw6 = (M51jw6 & T51jw6);
assign T51jw6 = (~(A61jw6 & Uxyiw6));
assign A61jw6 = (Kxb7z6[29] & H61jw6);
assign M51jw6 = (~(Lt3ov6 & O61jw6));
assign O61jw6 = (~(V61jw6 & Quziw6));
assign V61jw6 = (C71jw6 & J71jw6);
assign J71jw6 = (H61jw6 | Ninnv6);
assign H61jw6 = (Q71jw6 | Rje7z6[29]);
assign C71jw6 = (~(Ofnnv6 & Q71jw6));
assign Y41jw6 = (X71jw6 & E81jw6);
assign E81jw6 = (~(F7ziw6 & Rb3ov6));
assign X71jw6 = (~(J73ov6 & Nn3ov6));
assign K41jw6 = (L81jw6 & S81jw6);
assign S81jw6 = (Z81jw6 & G91jw6);
assign G91jw6 = (~(R6ziw6 & Kb3ov6));
assign Z81jw6 = (~(T0ziw6 & Rje7z6[29]));
assign L81jw6 = (N91jw6 & U91jw6);
assign U91jw6 = (Ryfov6 | Ba1jw6);
assign Ba1jw6 = (!Q71jw6);
assign N91jw6 = (~(L0g7z6[29] & J2ziw6));
assign W31jw6 = (Ia1jw6 & Pa1jw6);
assign Pa1jw6 = (Wa1jw6 & Db1jw6);
assign Db1jw6 = (Kb1jw6 & Rb1jw6);
assign Rb1jw6 = (~(Cqf7z6[13] & Q2ziw6));
assign Kb1jw6 = (~(L0g7z6[13] & O1ziw6));
assign Wa1jw6 = (Yb1jw6 & Fc1jw6);
assign Fc1jw6 = (~(U4ziw6 & V1c7z6[29]));
assign Yb1jw6 = (~(B5ziw6 & S7gdt6));
assign Ia1jw6 = (Mc1jw6 & Tc1jw6);
assign Tc1jw6 = (Ad1jw6 & Hd1jw6);
assign Hd1jw6 = (~(Z3ziw6 & E3c7z6[2]));
assign Ad1jw6 = (~(Sxkdt6 & Oztiw6));
assign Mc1jw6 = (Yq2ov6 & T7ziw6);
assign Yq2ov6 = (Od1jw6 & Vd1jw6);
assign Vd1jw6 = (~(Ce1jw6 & Dzmnv6));
assign Ce1jw6 = (~(Kzmnv6 | Icziw6));
assign Od1jw6 = (~(Je1jw6 & Ubziw6));
assign Je1jw6 = (~(Dzmnv6 ^ Kzmnv6));
assign Kzmnv6 = (Qe1jw6 ^ Mennv6);
assign Qe1jw6 = (~(Xe1jw6 & Ef1jw6));
assign Ef1jw6 = (Lf1jw6 & Sf1jw6);
assign Sf1jw6 = (Zf1jw6 & Gg1jw6);
assign Gg1jw6 = (~(Su0jw6 & Yxf7z6[31]));
assign Zf1jw6 = (Ng1jw6 & Ug1jw6);
assign Ug1jw6 = (~(Yxf7z6[29] & Nv0jw6));
assign Ng1jw6 = (~(Yxf7z6[30] & Uv0jw6));
assign Lf1jw6 = (Bh1jw6 & Ih1jw6);
assign Ih1jw6 = (~(Pw0jw6 & Yxf7z6[32]));
assign Bh1jw6 = (~(Ph1jw6 & Rdziw6));
assign Xe1jw6 = (Wh1jw6 & Di1jw6);
assign Di1jw6 = (Ki1jw6 & Ri1jw6);
assign Ri1jw6 = (~(Onf7z6[29] & My0jw6));
assign Ki1jw6 = (Yi1jw6 & Fj1jw6);
assign Fj1jw6 = (~(Hz0jw6 & Kxb7z6[29]));
assign Yi1jw6 = (~(Oz0jw6 & Fhc7z6[29]));
assign Wh1jw6 = (Mj1jw6 & Tj1jw6);
assign Tj1jw6 = (~(Alf7z6[13] & J01jw6));
assign Mj1jw6 = (~(Alf7z6[29] & Q01jw6));
assign Dzmnv6 = (~(Ak1jw6 ^ Tennv6));
assign Ak1jw6 = (~(Hk1jw6 & Ok1jw6));
assign Ok1jw6 = (~(Yxf7z6[13] & Laziw6));
assign Hk1jw6 = (Vk1jw6 & Cl1jw6);
assign Cl1jw6 = (~(Yxf7z6[29] & Gbziw6));
assign Vk1jw6 = (~(Kxb7z6[29] & Nbziw6));
assign Olz7v6 = (Tbbov6 ? vis_r0_o[28] : C7aov6);
assign Hlz7v6 = (Tbbov6 ? vis_r0_o[27] : S2gov6);
assign Alz7v6 = (Tbbov6 ? vis_r0_o[26] : W7xiw6);
assign Tkz7v6 = (Tbbov6 ? vis_r0_o[25] : R7yiw6);
assign Mkz7v6 = (Tbbov6 ? vis_r0_o[24] : Y7yiw6);
assign Fkz7v6 = (Tbbov6 ? vis_r0_o[23] : F8yiw6);
assign Yjz7v6 = (Tbbov6 ? vis_r0_o[22] : M8yiw6);
assign Rjz7v6 = (Tbbov6 ? vis_r0_o[21] : T8yiw6);
assign Kjz7v6 = (Tbbov6 ? vis_r0_o[20] : A9yiw6);
assign Djz7v6 = (Tbbov6 ? vis_r0_o[19] : H9yiw6);
assign Wiz7v6 = (Tbbov6 ? vis_r0_o[18] : Zqxiw6);
assign Piz7v6 = (Tbbov6 ? vis_r0_o[17] : O9yiw6);
assign Iiz7v6 = (Tbbov6 ? vis_r0_o[16] : V9yiw6);
assign Biz7v6 = (Tbbov6 ? vis_r0_o[15] : Qccov6);
assign Uhz7v6 = (Tbbov6 ? vis_r0_o[14] : Cayiw6);
assign Nhz7v6 = (Tbbov6 ? vis_r0_o[13] : Jayiw6);
assign Ghz7v6 = (Tbbov6 ? vis_r0_o[12] : Qayiw6);
assign Zgz7v6 = (Tbbov6 ? vis_r0_o[11] : Xayiw6);
assign Sgz7v6 = (Tbbov6 ? vis_r0_o[10] : T1yiw6);
assign Lgz7v6 = (Tbbov6 ? vis_r0_o[9] : Lbyiw6);
assign Egz7v6 = (Tbbov6 ? vis_r0_o[8] : W7kov6);
assign Xfz7v6 = (Tbbov6 ? vis_r0_o[7] : Sbyiw6);
assign Qfz7v6 = (Tbbov6 ? vis_r0_o[6] : Zbyiw6);
assign Jfz7v6 = (Tbbov6 ? vis_r0_o[5] : Gcyiw6);
assign Tbbov6 = (!Jl1jw6);
assign Cfz7v6 = (Jl1jw6 ? W6lov6 : vis_r0_o[4]);
assign Vez7v6 = (Jl1jw6 ? Ncyiw6 : vis_r0_o[3]);
assign Oez7v6 = (Jl1jw6 ? Bskov6 : vis_r0_o[2]);
assign Bskov6 = (Spyiw6 ? As97z6 : Gli7z6[2]);
assign As97z6 = (~(Ql1jw6 & Xl1jw6));
assign Xl1jw6 = (~(Nqyiw6 & Qo0ov6));
assign Ql1jw6 = (Em1jw6 & Lm1jw6);
assign Lm1jw6 = (~(Pdc7z6[2] & Ouyiw6));
assign Em1jw6 = (~(Vuyiw6 & Sm1jw6));
assign Sm1jw6 = (~(Zm1jw6 & Gn1jw6));
assign Gn1jw6 = (Nn1jw6 & Un1jw6);
assign Un1jw6 = (Bo1jw6 & Io1jw6);
assign Io1jw6 = (Po1jw6 & Wo1jw6);
assign Wo1jw6 = (~(Dp1jw6 & Kp1jw6));
assign Dp1jw6 = (~(Quziw6 & Rp1jw6));
assign Rp1jw6 = (~(Yp1jw6 & Fq1jw6));
assign Yp1jw6 = (~(Ninnv6 | Rje7z6[2]));
assign Po1jw6 = (~(Rje7z6[2] & Mq1jw6));
assign Mq1jw6 = (T0ziw6 | Tq1jw6);
assign Tq1jw6 = (Uxyiw6 & Kxb7z6[2]);
assign Bo1jw6 = (Ar1jw6 & Hr1jw6);
assign Hr1jw6 = (~(Or1jw6 & Vr1jw6));
assign Or1jw6 = (~(Cs1jw6 & Js1jw6));
assign Js1jw6 = (~(Uxyiw6 & Kxb7z6[2]));
assign Cs1jw6 = (Qs1jw6 & Ryfov6);
assign Qs1jw6 = (~(Ofnnv6 & Kp1jw6));
assign Ar1jw6 = (~(Svziw6 & Dknnv6));
assign Dknnv6 = (~(Xs1jw6 & Et1jw6));
assign Et1jw6 = (Lt1jw6 & St1jw6);
assign St1jw6 = (~(Zt1jw6 & Gu1jw6));
assign Zt1jw6 = (Nu1jw6 & I40jw6);
assign Lt1jw6 = (~(P40jw6 & Uu1jw6));
assign Xs1jw6 = (Bv1jw6 & Iv1jw6);
assign Iv1jw6 = (~(Bxziw6 & Pv1jw6));
assign Bv1jw6 = (~(Ua0jw6 & Wv1jw6));
assign Nn1jw6 = (Dw1jw6 & Kw1jw6);
assign Kw1jw6 = (Rw1jw6 & Yw1jw6);
assign Yw1jw6 = (~(Hk3ov6 & C73ov6));
assign Rw1jw6 = (~(Ol0jw6 & Un3ov6));
assign Dw1jw6 = (Fx1jw6 & Mx1jw6);
assign Mx1jw6 = (~(Jm0jw6 & Tx1jw6));
assign Fx1jw6 = (~(J73ov6 & Db3ov6));
assign Zm1jw6 = (Ay1jw6 & Hy1jw6);
assign Hy1jw6 = (Oy1jw6 & Vy1jw6);
assign Vy1jw6 = (Cz1jw6 & Jz1jw6);
assign Jz1jw6 = (~(L0g7z6[2] & J2ziw6));
assign Cz1jw6 = (~(L0g7z6[18] & Q2ziw6));
assign Oy1jw6 = (Qz1jw6 & Xz1jw6);
assign Xz1jw6 = (~(O1ziw6 & Onf7z6[2]));
assign Qz1jw6 = (~(U4ziw6 & E3c7z6[2]));
assign Ay1jw6 = (E02jw6 & Rq2ov6);
assign Rq2ov6 = (L02jw6 & S02jw6);
assign S02jw6 = (~(Z02jw6 & Pymnv6));
assign Z02jw6 = (~(Wymnv6 | Icziw6));
assign L02jw6 = (~(G12jw6 & Ubziw6));
assign G12jw6 = (~(Pymnv6 ^ Wymnv6));
assign Wymnv6 = (N12jw6 ^ Mennv6);
assign N12jw6 = (~(U12jw6 & B22jw6));
assign B22jw6 = (I22jw6 & P22jw6);
assign P22jw6 = (W22jw6 & D32jw6);
assign D32jw6 = (~(Yxf7z6[4] & Su0jw6));
assign W22jw6 = (K32jw6 & R32jw6);
assign R32jw6 = (~(Yxf7z6[2] & Nv0jw6));
assign K32jw6 = (~(Yxf7z6[3] & Uv0jw6));
assign I22jw6 = (Y32jw6 & F42jw6);
assign F42jw6 = (~(Yxf7z6[5] & Pw0jw6));
assign Y32jw6 = (M42jw6 | Dx0jw6);
assign U12jw6 = (T42jw6 & A52jw6);
assign A52jw6 = (H52jw6 & O52jw6);
assign O52jw6 = (~(Onf7z6[2] & My0jw6));
assign H52jw6 = (V52jw6 & C62jw6);
assign C62jw6 = (~(Hz0jw6 & Kxb7z6[2]));
assign V52jw6 = (~(Oz0jw6 & E3c7z6[2]));
assign T42jw6 = (J62jw6 & Q62jw6);
assign Q62jw6 = (~(Onf7z6[18] & J01jw6));
assign J62jw6 = (~(Alf7z6[2] & Q01jw6));
assign Pymnv6 = (~(X62jw6 ^ Tennv6));
assign X62jw6 = (~(E72jw6 & L72jw6));
assign L72jw6 = (~(Yxf7z6[2] & Gbziw6));
assign E72jw6 = (~(Kxb7z6[2] & Nbziw6));
assign E02jw6 = (S72jw6 & Z72jw6);
assign Z72jw6 = (~(Z3ziw6 & Fhc7z6[29]));
assign S72jw6 = (~(Vimdt6 & Oztiw6));
assign Hez7v6 = (Jl1jw6 ? Nv9ov6 : vis_r0_o[1]);
assign Jl1jw6 = (~(Vnyiw6 | Xhyiw6));
assign Xhyiw6 = (Fmyiw6 | Ylyiw6);
assign Vnyiw6 = (!Rlyiw6);
assign Rlyiw6 = (G82jw6 & Liyiw6);
assign G82jw6 = (Mlziw6 & Bkyiw6);
assign Nv9ov6 = (Spyiw6 ? N82jw6 : Gli7z6[1]);
assign N82jw6 = (Amziw6 & Mu97z6);
assign Mu97z6 = (~(U82jw6 & B92jw6));
assign B92jw6 = (Z11jw6 | Kdmhw6);
assign U82jw6 = (I92jw6 & P92jw6);
assign P92jw6 = (~(Pdc7z6[1] & Ouyiw6));
assign I92jw6 = (~(Vuyiw6 & W92jw6));
assign W92jw6 = (~(Da2jw6 & Ka2jw6));
assign Ka2jw6 = (Ra2jw6 & Ya2jw6);
assign Ya2jw6 = (Fb2jw6 & Mb2jw6);
assign Mb2jw6 = (Tb2jw6 & Ac2jw6);
assign Ac2jw6 = (~(Hc2jw6 & Jm0jw6));
assign Hc2jw6 = (Nob7z6[1] & Rslov6);
assign Tb2jw6 = (Oc2jw6 & Vc2jw6);
assign Vc2jw6 = (~(Cd2jw6 & Uxyiw6));
assign Cd2jw6 = (Kxb7z6[1] & Jd2jw6);
assign Oc2jw6 = (~(Qd2jw6 & C1gov6));
assign Qd2jw6 = (Bqziw6 & Jjbdt6);
assign Fb2jw6 = (Xd2jw6 & Ee2jw6);
assign Ee2jw6 = (~(Le2jw6 & Se2jw6));
assign Le2jw6 = (~(Ze2jw6 & Quziw6));
assign Ze2jw6 = (Gf2jw6 & Nf2jw6);
assign Nf2jw6 = (Jd2jw6 | Ninnv6);
assign Jd2jw6 = (Uf2jw6 | Rje7z6[1]);
assign Gf2jw6 = (~(Ofnnv6 & Uf2jw6));
assign Xd2jw6 = (~(Ol0jw6 & Io3ov6));
assign Ra2jw6 = (Bg2jw6 & Ig2jw6);
assign Ig2jw6 = (Pg2jw6 & Wg2jw6);
assign Wg2jw6 = (Lf3ov6 | U93ov6);
assign Pg2jw6 = (~(Ak3ov6 & C73ov6));
assign Bg2jw6 = (Dh2jw6 & Kh2jw6);
assign Kh2jw6 = (~(T0ziw6 & Rje7z6[1]));
assign Dh2jw6 = (Ryfov6 | Rh2jw6);
assign Da2jw6 = (Yh2jw6 & Fi2jw6);
assign Fi2jw6 = (Mi2jw6 & Ti2jw6);
assign Ti2jw6 = (Aj2jw6 & Hj2jw6);
assign Hj2jw6 = (~(L0g7z6[1] & J2ziw6));
assign Aj2jw6 = (~(L0g7z6[17] & Q2ziw6));
assign Mi2jw6 = (Oj2jw6 & Vj2jw6);
assign Vj2jw6 = (~(O1ziw6 & Onf7z6[1]));
assign Oj2jw6 = (~(U4ziw6 & E3c7z6[1]));
assign Yh2jw6 = (Ck2jw6 & Jk2jw6);
assign Jk2jw6 = (Qk2jw6 & Xk2jw6);
assign Xk2jw6 = (~(Z3ziw6 & Fhc7z6[30]));
assign Qk2jw6 = (~(Svziw6 & Kknnv6));
assign Ck2jw6 = (As2ov6 & El2jw6);
assign El2jw6 = (~(Ykmdt6 & Oztiw6));
assign As2ov6 = (Ll2jw6 & Sl2jw6);
assign Sl2jw6 = (~(Zl2jw6 & N4nnv6));
assign Zl2jw6 = (~(U4nnv6 | Icziw6));
assign Ll2jw6 = (~(Gm2jw6 & Ubziw6));
assign Gm2jw6 = (~(N4nnv6 ^ U4nnv6));
assign U4nnv6 = (Nm2jw6 ^ Mennv6);
assign Nm2jw6 = (~(Um2jw6 & Bn2jw6));
assign Bn2jw6 = (In2jw6 & Pn2jw6);
assign Pn2jw6 = (Wn2jw6 & Do2jw6);
assign Do2jw6 = (~(Yxf7z6[3] & Su0jw6));
assign Wn2jw6 = (Ko2jw6 & Ro2jw6);
assign Ro2jw6 = (~(Yxf7z6[1] & Nv0jw6));
assign Ko2jw6 = (~(Yxf7z6[2] & Uv0jw6));
assign In2jw6 = (Yo2jw6 & Fp2jw6);
assign Fp2jw6 = (~(Yxf7z6[4] & Pw0jw6));
assign Yo2jw6 = (Mp2jw6 | Dx0jw6);
assign Um2jw6 = (Tp2jw6 & Aq2jw6);
assign Aq2jw6 = (Hq2jw6 & Oq2jw6);
assign Oq2jw6 = (~(Onf7z6[1] & My0jw6));
assign Hq2jw6 = (Vq2jw6 & Cr2jw6);
assign Cr2jw6 = (~(Hz0jw6 & Kxb7z6[1]));
assign Vq2jw6 = (~(Oz0jw6 & E3c7z6[1]));
assign Tp2jw6 = (Jr2jw6 & Qr2jw6);
assign Qr2jw6 = (~(Onf7z6[17] & J01jw6));
assign Jr2jw6 = (~(Alf7z6[1] & Q01jw6));
assign N4nnv6 = (~(Xr2jw6 ^ Tennv6));
assign Xr2jw6 = (~(Es2jw6 & Ls2jw6));
assign Ls2jw6 = (~(Kxb7z6[1] & S11jw6));
assign S11jw6 = (~(Ss2jw6 & Zs2jw6));
assign Ss2jw6 = (Dx0jw6 | Usbdt6);
assign Es2jw6 = (~(Yxf7z6[1] & Gbziw6));
assign Amziw6 = (!Gt2jw6);
assign Aez7v6 = (Ut2jw6 ? A4a7z6 : Nt2jw6);
assign Nt2jw6 = (Pkbet6 | C3yiw6);
assign Tdz7v6 = (~(Bu2jw6 & Iu2jw6));
assign Iu2jw6 = (~(Eji7z6[1] & C3yiw6));
assign Bu2jw6 = (Pu2jw6 & Wu2jw6);
assign Wu2jw6 = (~(Bhi7z6[1] & X3yiw6));
assign Pu2jw6 = (~(E4yiw6 & vis_pc_o[1]));
assign Mdz7v6 = (~(Dv2jw6 & Kv2jw6));
assign Kv2jw6 = (~(Eji7z6[3] & C3yiw6));
assign Dv2jw6 = (Rv2jw6 & Yv2jw6);
assign Yv2jw6 = (~(Bhi7z6[3] & X3yiw6));
assign Rv2jw6 = (~(E4yiw6 & vis_pc_o[3]));
assign Fdz7v6 = (~(Fw2jw6 & Mw2jw6));
assign Mw2jw6 = (~(Eji7z6[4] & C3yiw6));
assign Fw2jw6 = (Tw2jw6 & Ax2jw6);
assign Ax2jw6 = (~(Bhi7z6[4] & X3yiw6));
assign Tw2jw6 = (~(E4yiw6 & vis_pc_o[4]));
assign Ycz7v6 = (~(Hx2jw6 & Ox2jw6));
assign Ox2jw6 = (Vx2jw6 & Cy2jw6);
assign Cy2jw6 = (Eu9ov6 | Jy2jw6);
assign Vx2jw6 = (Qy2jw6 & Xy2jw6);
assign Xy2jw6 = (~(Gv9ov6 & W6lov6));
assign W6lov6 = (Spyiw6 ? Iw97z6 : Gli7z6[4]);
assign Qy2jw6 = (~(Uv9ov6 & Iw97z6));
assign Iw97z6 = (~(Ez2jw6 & Lz2jw6));
assign Lz2jw6 = (~(Nqyiw6 & Og0ov6));
assign Ez2jw6 = (Sz2jw6 & Zz2jw6);
assign Zz2jw6 = (~(Pdc7z6[4] & Ouyiw6));
assign Sz2jw6 = (~(Vuyiw6 & G03jw6));
assign G03jw6 = (~(N03jw6 & U03jw6));
assign U03jw6 = (B13jw6 & I13jw6);
assign I13jw6 = (P13jw6 & W13jw6);
assign W13jw6 = (D23jw6 & K23jw6);
assign K23jw6 = (~(R23jw6 & Uxyiw6));
assign R23jw6 = (Kxb7z6[4] & Y23jw6);
assign D23jw6 = (~(F33jw6 & Jm0jw6));
assign F33jw6 = (Nob7z6[4] & Rslov6);
assign P13jw6 = (M33jw6 & T33jw6);
assign T33jw6 = (~(Et3ov6 & A43jw6));
assign A43jw6 = (~(H43jw6 & Quziw6));
assign H43jw6 = (O43jw6 & V43jw6);
assign V43jw6 = (Y23jw6 | Ninnv6);
assign Y23jw6 = (C53jw6 | Rje7z6[4]);
assign O43jw6 = (~(Ofnnv6 & C53jw6));
assign M33jw6 = (~(Svziw6 & Pjnnv6));
assign Pjnnv6 = (Bxziw6 | P40jw6);
assign B13jw6 = (J53jw6 & Q53jw6);
assign Q53jw6 = (X53jw6 & E63jw6);
assign E63jw6 = (~(Ol0jw6 & Em3ov6));
assign X53jw6 = (~(Ki3ov6 & C73ov6));
assign J53jw6 = (L63jw6 & S63jw6);
assign S63jw6 = (~(J73ov6 & Xe3ov6));
assign L63jw6 = (~(T0ziw6 & Rje7z6[4]));
assign N03jw6 = (Z63jw6 & G73jw6);
assign G73jw6 = (N73jw6 & U73jw6);
assign U73jw6 = (B83jw6 & I83jw6);
assign I83jw6 = (Ryfov6 | P83jw6);
assign B83jw6 = (~(L0g7z6[4] & J2ziw6));
assign N73jw6 = (W83jw6 & D93jw6);
assign D93jw6 = (~(L0g7z6[20] & Q2ziw6));
assign W83jw6 = (~(O1ziw6 & Onf7z6[4]));
assign Z63jw6 = (K93jw6 & R93jw6);
assign R93jw6 = (Y93jw6 & Fa3jw6);
assign Fa3jw6 = (~(U4ziw6 & E3c7z6[4]));
assign Y93jw6 = (~(Z3ziw6 & Fhc7z6[27]));
assign K93jw6 = (Tr2ov6 & Ma3jw6);
assign Ma3jw6 = (~(Pemdt6 & Oztiw6));
assign Tr2ov6 = (Ta3jw6 & Ab3jw6);
assign Ab3jw6 = (~(Hb3jw6 & Zwmnv6));
assign Hb3jw6 = (~(Gxmnv6 | Icziw6));
assign Ta3jw6 = (~(Ob3jw6 & Ubziw6));
assign Ob3jw6 = (~(Zwmnv6 ^ Gxmnv6));
assign Gxmnv6 = (Vb3jw6 ^ Mennv6);
assign Vb3jw6 = (~(Cc3jw6 & Jc3jw6));
assign Jc3jw6 = (Qc3jw6 & Xc3jw6);
assign Xc3jw6 = (Ed3jw6 & Ld3jw6);
assign Ld3jw6 = (~(Yxf7z6[6] & Su0jw6));
assign Ed3jw6 = (Sd3jw6 & Zd3jw6);
assign Zd3jw6 = (~(Yxf7z6[4] & Nv0jw6));
assign Sd3jw6 = (~(Yxf7z6[5] & Uv0jw6));
assign Qc3jw6 = (Ge3jw6 & Ne3jw6);
assign Ne3jw6 = (~(Yxf7z6[7] & Pw0jw6));
assign Ge3jw6 = (~(Ue3jw6 & Rdziw6));
assign Cc3jw6 = (Bf3jw6 & If3jw6);
assign If3jw6 = (Pf3jw6 & Wf3jw6);
assign Wf3jw6 = (~(Onf7z6[4] & My0jw6));
assign Pf3jw6 = (Dg3jw6 & Kg3jw6);
assign Kg3jw6 = (~(Hz0jw6 & Kxb7z6[4]));
assign Dg3jw6 = (~(Oz0jw6 & E3c7z6[4]));
assign Bf3jw6 = (Rg3jw6 & Yg3jw6);
assign Yg3jw6 = (~(Onf7z6[20] & J01jw6));
assign Rg3jw6 = (~(Alf7z6[4] & Q01jw6));
assign Zwmnv6 = (~(Fh3jw6 ^ Tennv6));
assign Fh3jw6 = (~(Mh3jw6 & Th3jw6));
assign Th3jw6 = (~(Yxf7z6[4] & Gbziw6));
assign Mh3jw6 = (~(Kxb7z6[4] & Nbziw6));
assign Hx2jw6 = (Ai3jw6 & Hi3jw6);
assign Hi3jw6 = (~(Pw9ov6 & Kxb7z6[4]));
assign Ai3jw6 = (Oi3jw6 & Vi3jw6);
assign Vi3jw6 = (~(Kx9ov6 & vis_pc_o[4]));
assign Oi3jw6 = (~(Gli7z6[4] & Rx9ov6));
assign Rcz7v6 = (~(Cj3jw6 & Jj3jw6));
assign Jj3jw6 = (~(Eji7z6[5] & C3yiw6));
assign Cj3jw6 = (Qj3jw6 & Xj3jw6);
assign Xj3jw6 = (~(Bhi7z6[5] & X3yiw6));
assign Qj3jw6 = (~(E4yiw6 & vis_pc_o[5]));
assign Kcz7v6 = (~(Ek3jw6 & Lk3jw6));
assign Lk3jw6 = (~(Eji7z6[6] & C3yiw6));
assign Ek3jw6 = (Sk3jw6 & Zk3jw6);
assign Zk3jw6 = (~(Bhi7z6[6] & X3yiw6));
assign Sk3jw6 = (~(E4yiw6 & vis_pc_o[6]));
assign Dcz7v6 = (~(Gl3jw6 & Nl3jw6));
assign Nl3jw6 = (~(Eji7z6[7] & C3yiw6));
assign Gl3jw6 = (Ul3jw6 & Bm3jw6);
assign Bm3jw6 = (~(Bhi7z6[7] & X3yiw6));
assign Ul3jw6 = (~(E4yiw6 & vis_pc_o[7]));
assign Wbz7v6 = (~(Im3jw6 & Pm3jw6));
assign Pm3jw6 = (~(Eji7z6[8] & C3yiw6));
assign Im3jw6 = (Wm3jw6 & Dn3jw6);
assign Dn3jw6 = (~(Bhi7z6[8] & X3yiw6));
assign Wm3jw6 = (~(E4yiw6 & vis_pc_o[8]));
assign Pbz7v6 = (~(Kn3jw6 & Rn3jw6));
assign Rn3jw6 = (Yn3jw6 & Fo3jw6);
assign Fo3jw6 = (Eu9ov6 | Mo3jw6);
assign Yn3jw6 = (To3jw6 & Ap3jw6);
assign Ap3jw6 = (~(Gv9ov6 & W7kov6));
assign W7kov6 = (Spyiw6 ? Aw97z6 : Gli7z6[8]);
assign To3jw6 = (~(Uv9ov6 & Aw97z6));
assign Aw97z6 = (~(Hp3jw6 & Op3jw6));
assign Op3jw6 = (~(Nqyiw6 & K00ov6));
assign Hp3jw6 = (Vp3jw6 & Cq3jw6);
assign Cq3jw6 = (~(Pdc7z6[8] & Ouyiw6));
assign Vp3jw6 = (~(Vuyiw6 & Jq3jw6));
assign Jq3jw6 = (~(Qq3jw6 & Xq3jw6));
assign Xq3jw6 = (Er3jw6 & Lr3jw6);
assign Lr3jw6 = (Sr3jw6 & Zr3jw6);
assign Zr3jw6 = (Gs3jw6 & Ns3jw6);
assign Gs3jw6 = (~(Us3jw6 & Uxyiw6));
assign Us3jw6 = (Kxb7z6[8] & Bt3jw6);
assign Sr3jw6 = (It3jw6 & Pt3jw6);
assign Pt3jw6 = (~(Wt3jw6 & Jm0jw6));
assign Wt3jw6 = (Nob7z6[8] & Rslov6);
assign It3jw6 = (~(Du3jw6 & Ku3jw6));
assign Du3jw6 = (~(Ru3jw6 & Quziw6));
assign Ru3jw6 = (Yu3jw6 & Fv3jw6);
assign Fv3jw6 = (Bt3jw6 | Ninnv6);
assign Bt3jw6 = (Mv3jw6 | Rje7z6[8]);
assign Yu3jw6 = (~(Ofnnv6 & Mv3jw6));
assign Er3jw6 = (Tv3jw6 & Aw3jw6);
assign Aw3jw6 = (Hw3jw6 & Ow3jw6);
assign Ow3jw6 = (~(Bo3ov6 & C73ov6));
assign Hw3jw6 = (~(Tj3ov6 & Ug3ov6));
assign Tv3jw6 = (Vw3jw6 & Cx3jw6);
assign Cx3jw6 = (Lf3ov6 | Ba3ov6);
assign Vw3jw6 = (~(T0ziw6 & Rje7z6[8]));
assign Qq3jw6 = (Jx3jw6 & Qx3jw6);
assign Qx3jw6 = (Xx3jw6 & Ey3jw6);
assign Ey3jw6 = (Ly3jw6 & Sy3jw6);
assign Sy3jw6 = (Ryfov6 | Zy3jw6);
assign Ly3jw6 = (~(L0g7z6[8] & J2ziw6));
assign Xx3jw6 = (Gz3jw6 & Nz3jw6);
assign Nz3jw6 = (~(L0g7z6[24] & Q2ziw6));
assign Gz3jw6 = (~(O1ziw6 & Onf7z6[8]));
assign Jx3jw6 = (Uz3jw6 & B04jw6);
assign B04jw6 = (I04jw6 & P04jw6);
assign P04jw6 = (~(U4ziw6 & Fhc7z6[8]));
assign I04jw6 = (~(Z3ziw6 & Fhc7z6[23]));
assign Uz3jw6 = (Os2ov6 & W04jw6);
assign W04jw6 = (~(D6mdt6 & Oztiw6));
assign Os2ov6 = (D14jw6 & K14jw6);
assign K14jw6 = (~(R14jw6 & Vumnv6));
assign R14jw6 = (~(Cvmnv6 | Icziw6));
assign D14jw6 = (~(Y14jw6 & Ubziw6));
assign Y14jw6 = (~(Vumnv6 ^ Cvmnv6));
assign Cvmnv6 = (F24jw6 ^ Mennv6);
assign F24jw6 = (~(M24jw6 & T24jw6));
assign T24jw6 = (A34jw6 & H34jw6);
assign H34jw6 = (O34jw6 & V34jw6);
assign V34jw6 = (~(Yxf7z6[10] & Su0jw6));
assign O34jw6 = (C44jw6 & J44jw6);
assign J44jw6 = (~(Yxf7z6[8] & Nv0jw6));
assign C44jw6 = (~(Yxf7z6[9] & Uv0jw6));
assign A34jw6 = (Q44jw6 & X44jw6);
assign X44jw6 = (~(Yxf7z6[11] & Pw0jw6));
assign Q44jw6 = (E54jw6 | Dx0jw6);
assign M24jw6 = (L54jw6 & S54jw6);
assign S54jw6 = (Z54jw6 & G64jw6);
assign G64jw6 = (~(Onf7z6[8] & My0jw6));
assign Z54jw6 = (N64jw6 & U64jw6);
assign U64jw6 = (~(Hz0jw6 & Kxb7z6[8]));
assign N64jw6 = (~(Oz0jw6 & Fhc7z6[8]));
assign L54jw6 = (B74jw6 & I74jw6);
assign I74jw6 = (~(Onf7z6[24] & J01jw6));
assign B74jw6 = (~(Alf7z6[8] & Q01jw6));
assign Vumnv6 = (~(P74jw6 ^ Tennv6));
assign P74jw6 = (~(W74jw6 & D84jw6));
assign D84jw6 = (~(Yxf7z6[8] & Gbziw6));
assign W74jw6 = (~(Kxb7z6[8] & Nbziw6));
assign Kn3jw6 = (K84jw6 & R84jw6);
assign R84jw6 = (~(Pw9ov6 & Kxb7z6[8]));
assign K84jw6 = (Y84jw6 & F94jw6);
assign F94jw6 = (~(Kx9ov6 & vis_pc_o[8]));
assign Y84jw6 = (~(Gli7z6[8] & Rx9ov6));
assign Ibz7v6 = (~(M94jw6 & T94jw6));
assign T94jw6 = (~(Eji7z6[9] & C3yiw6));
assign M94jw6 = (Aa4jw6 & Ha4jw6);
assign Ha4jw6 = (~(Bhi7z6[9] & X3yiw6));
assign Aa4jw6 = (~(E4yiw6 & vis_pc_o[9]));
assign Bbz7v6 = (~(Oa4jw6 & Va4jw6));
assign Va4jw6 = (~(Eji7z6[10] & C3yiw6));
assign Oa4jw6 = (Cb4jw6 & Jb4jw6);
assign Jb4jw6 = (~(Bhi7z6[10] & X3yiw6));
assign Cb4jw6 = (~(E4yiw6 & vis_pc_o[10]));
assign Uaz7v6 = (~(Qb4jw6 & Xb4jw6));
assign Xb4jw6 = (Ec4jw6 & Lc4jw6);
assign Lc4jw6 = (Eu9ov6 | Sc4jw6);
assign Ec4jw6 = (Zc4jw6 & Gd4jw6);
assign Gd4jw6 = (~(Gv9ov6 & T1yiw6));
assign T1yiw6 = (Gninv6 ? Gli7z6[10] : Gx97z6);
assign Zc4jw6 = (~(Uv9ov6 & Gx97z6));
assign Gx97z6 = (~(Nd4jw6 & Ud4jw6));
assign Ud4jw6 = (~(Nqyiw6 & Isznv6));
assign Nd4jw6 = (Be4jw6 & Ie4jw6);
assign Ie4jw6 = (~(Pdc7z6[10] & Ouyiw6));
assign Be4jw6 = (~(Vuyiw6 & Pe4jw6));
assign Pe4jw6 = (~(We4jw6 & Df4jw6));
assign Df4jw6 = (Kf4jw6 & Rf4jw6);
assign Rf4jw6 = (Yf4jw6 & Fg4jw6);
assign Fg4jw6 = (Mg4jw6 & Ns3jw6);
assign Mg4jw6 = (~(Tg4jw6 & Uxyiw6));
assign Tg4jw6 = (Kxb7z6[10] & Ah4jw6);
assign Yf4jw6 = (Hh4jw6 & Oh4jw6);
assign Oh4jw6 = (~(Vh4jw6 & Ci4jw6));
assign Vh4jw6 = (~(Ji4jw6 & Quziw6));
assign Ji4jw6 = (Qi4jw6 & Xi4jw6);
assign Xi4jw6 = (Ah4jw6 | Ninnv6);
assign Ah4jw6 = (Ej4jw6 | Rje7z6[10]);
assign Qi4jw6 = (~(Ofnnv6 & Ej4jw6));
assign Hh4jw6 = (~(Hk3ov6 & Ug3ov6));
assign Kf4jw6 = (Lj4jw6 & Sj4jw6);
assign Sj4jw6 = (Zj4jw6 & Gk4jw6);
assign Gk4jw6 = (~(Un3ov6 & C73ov6));
assign Zj4jw6 = (~(J73ov6 & Vd3ov6));
assign Lj4jw6 = (Nk4jw6 & Uk4jw6);
assign Uk4jw6 = (~(T0ziw6 & Rje7z6[10]));
assign Nk4jw6 = (Ryfov6 | Bl4jw6);
assign We4jw6 = (Il4jw6 & Pl4jw6);
assign Pl4jw6 = (Wl4jw6 & Dm4jw6);
assign Dm4jw6 = (Km4jw6 & Rm4jw6);
assign Rm4jw6 = (~(L0g7z6[10] & J2ziw6));
assign Km4jw6 = (~(L0g7z6[26] & Q2ziw6));
assign Wl4jw6 = (Ym4jw6 & Fn4jw6);
assign Fn4jw6 = (~(O1ziw6 & Onf7z6[10]));
assign Ym4jw6 = (~(U4ziw6 & Fhc7z6[10]));
assign Il4jw6 = (Mn4jw6 & Hs2ov6);
assign Hs2ov6 = (Tn4jw6 & Ao4jw6);
assign Ao4jw6 = (~(Ho4jw6 & X9nnv6));
assign Ho4jw6 = (~(Eannv6 | Icziw6));
assign Tn4jw6 = (~(Oo4jw6 & Ubziw6));
assign Oo4jw6 = (~(X9nnv6 ^ Eannv6));
assign Eannv6 = (Vo4jw6 ^ Mennv6);
assign Vo4jw6 = (~(Cp4jw6 & Jp4jw6));
assign Jp4jw6 = (Qp4jw6 & Xp4jw6);
assign Xp4jw6 = (Eq4jw6 & Lq4jw6);
assign Lq4jw6 = (~(Yxf7z6[12] & Su0jw6));
assign Eq4jw6 = (Sq4jw6 & Zq4jw6);
assign Zq4jw6 = (~(Yxf7z6[10] & Nv0jw6));
assign Sq4jw6 = (~(Yxf7z6[11] & Uv0jw6));
assign Qp4jw6 = (Gr4jw6 & Nr4jw6);
assign Nr4jw6 = (~(Yxf7z6[13] & Pw0jw6));
assign Gr4jw6 = (Ur4jw6 | Dx0jw6);
assign Cp4jw6 = (Bs4jw6 & Is4jw6);
assign Is4jw6 = (Ps4jw6 & Ws4jw6);
assign Ws4jw6 = (~(Onf7z6[10] & My0jw6));
assign Ps4jw6 = (Dt4jw6 & Kt4jw6);
assign Kt4jw6 = (~(Hz0jw6 & Kxb7z6[10]));
assign Dt4jw6 = (~(Oz0jw6 & Fhc7z6[10]));
assign Bs4jw6 = (Rt4jw6 & Yt4jw6);
assign Yt4jw6 = (~(Onf7z6[26] & J01jw6));
assign Rt4jw6 = (~(Alf7z6[10] & Q01jw6));
assign X9nnv6 = (~(Fu4jw6 ^ Tennv6));
assign Fu4jw6 = (~(Mu4jw6 & Tu4jw6));
assign Tu4jw6 = (~(Yxf7z6[10] & Gbziw6));
assign Mu4jw6 = (~(Kxb7z6[10] & Nbziw6));
assign Mn4jw6 = (Av4jw6 & Hv4jw6);
assign Hv4jw6 = (~(Z3ziw6 & Fhc7z6[21]));
assign Av4jw6 = (~(X1mdt6 & Oztiw6));
assign Qb4jw6 = (Ov4jw6 & Vv4jw6);
assign Vv4jw6 = (~(Pw9ov6 & Kxb7z6[10]));
assign Ov4jw6 = (Cw4jw6 & Jw4jw6);
assign Jw4jw6 = (~(Kx9ov6 & vis_pc_o[10]));
assign Cw4jw6 = (~(Gli7z6[10] & Rx9ov6));
assign Naz7v6 = (~(Qw4jw6 & Xw4jw6));
assign Xw4jw6 = (~(Eji7z6[11] & C3yiw6));
assign Qw4jw6 = (Ex4jw6 & Lx4jw6);
assign Lx4jw6 = (~(Bhi7z6[11] & X3yiw6));
assign Ex4jw6 = (~(E4yiw6 & vis_pc_o[11]));
assign Gaz7v6 = (~(Sx4jw6 & Zx4jw6));
assign Zx4jw6 = (~(Eji7z6[12] & C3yiw6));
assign Sx4jw6 = (Gy4jw6 & Ny4jw6);
assign Ny4jw6 = (~(Bhi7z6[12] & X3yiw6));
assign Gy4jw6 = (~(E4yiw6 & vis_pc_o[12]));
assign Z9z7v6 = (~(Uy4jw6 & Bz4jw6));
assign Bz4jw6 = (~(Eji7z6[13] & C3yiw6));
assign Uy4jw6 = (Iz4jw6 & Pz4jw6);
assign Pz4jw6 = (~(Bhi7z6[13] & X3yiw6));
assign Iz4jw6 = (~(E4yiw6 & vis_pc_o[13]));
assign S9z7v6 = (~(Wz4jw6 & D05jw6));
assign D05jw6 = (~(Eji7z6[14] & C3yiw6));
assign Wz4jw6 = (K05jw6 & R05jw6);
assign R05jw6 = (~(Bhi7z6[14] & X3yiw6));
assign K05jw6 = (~(E4yiw6 & vis_pc_o[14]));
assign L9z7v6 = (~(Y05jw6 & F15jw6));
assign F15jw6 = (~(Eji7z6[15] & C3yiw6));
assign Y05jw6 = (M15jw6 & T15jw6);
assign T15jw6 = (~(Bhi7z6[15] & X3yiw6));
assign M15jw6 = (~(E4yiw6 & vis_pc_o[15]));
assign E9z7v6 = (~(A25jw6 & H25jw6));
assign H25jw6 = (O25jw6 & V25jw6);
assign V25jw6 = (Eu9ov6 | C35jw6);
assign O25jw6 = (J35jw6 & Q35jw6);
assign Q35jw6 = (~(Gv9ov6 & Qccov6));
assign Qccov6 = (Spyiw6 ? Kv97z6 : Gli7z6[15]);
assign J35jw6 = (~(Uv9ov6 & Kv97z6));
assign Kv97z6 = (~(X35jw6 & E45jw6));
assign E45jw6 = (~(Nqyiw6 & D8znv6));
assign X35jw6 = (L45jw6 & S45jw6);
assign S45jw6 = (~(Pdc7z6[15] & Ouyiw6));
assign L45jw6 = (~(Vuyiw6 & Z45jw6));
assign Z45jw6 = (~(G55jw6 & N55jw6));
assign N55jw6 = (U55jw6 & B65jw6);
assign B65jw6 = (I65jw6 & P65jw6);
assign P65jw6 = (W65jw6 & Ns3jw6);
assign W65jw6 = (~(D75jw6 & Uxyiw6));
assign D75jw6 = (Kxb7z6[15] & K75jw6);
assign I65jw6 = (R75jw6 & Y75jw6);
assign Y75jw6 = (~(F85jw6 & M85jw6));
assign F85jw6 = (~(T85jw6 & Quziw6));
assign T85jw6 = (A95jw6 & H95jw6);
assign H95jw6 = (K75jw6 | Ninnv6);
assign K75jw6 = (O95jw6 | Rje7z6[15]);
assign A95jw6 = (~(Ofnnv6 & O95jw6));
assign R75jw6 = (~(Ok3ov6 & Ug3ov6));
assign U55jw6 = (V95jw6 & Ca5jw6);
assign Ca5jw6 = (~(L0g7z6[15] & J2ziw6));
assign V95jw6 = (Ja5jw6 & Qa5jw6);
assign Qa5jw6 = (~(T0ziw6 & Rje7z6[15]));
assign Ja5jw6 = (Ryfov6 | Xa5jw6);
assign G55jw6 = (Eb5jw6 & Lb5jw6);
assign Lb5jw6 = (Sb5jw6 & Zb5jw6);
assign Zb5jw6 = (Gc5jw6 & Nc5jw6);
assign Nc5jw6 = (~(L0g7z6[31] & Q2ziw6));
assign Gc5jw6 = (~(O1ziw6 & Onf7z6[15]));
assign Sb5jw6 = (Uc5jw6 & Bd5jw6);
assign Bd5jw6 = (~(U4ziw6 & Fhc7z6[15]));
assign Uc5jw6 = (~(Z3ziw6 & Fhc7z6[16]));
assign Eb5jw6 = (Id5jw6 & Kp3ov6);
assign Kp3ov6 = (Pd5jw6 & Wd5jw6);
assign Wd5jw6 = (~(H8ziw6 & C73ov6));
assign Pd5jw6 = (~(J73ov6 & Y6ziw6));
assign Id5jw6 = (Eu2ov6 & De5jw6);
assign De5jw6 = (~(Irldt6 & Oztiw6));
assign Eu2ov6 = (Ke5jw6 & Re5jw6);
assign Re5jw6 = (~(Ye5jw6 & F7nnv6));
assign Ye5jw6 = (~(M7nnv6 | Icziw6));
assign Ke5jw6 = (~(Ff5jw6 & Ubziw6));
assign Ff5jw6 = (~(F7nnv6 ^ M7nnv6));
assign M7nnv6 = (Mf5jw6 ^ Mennv6);
assign Mf5jw6 = (~(Tf5jw6 & Ag5jw6));
assign Ag5jw6 = (Hg5jw6 & Og5jw6);
assign Og5jw6 = (Vg5jw6 & Ch5jw6);
assign Ch5jw6 = (~(Yxf7z6[17] & Su0jw6));
assign Vg5jw6 = (Jh5jw6 & Qh5jw6);
assign Qh5jw6 = (~(Nv0jw6 & Yxf7z6[15]));
assign Jh5jw6 = (~(Yxf7z6[16] & Uv0jw6));
assign Hg5jw6 = (Xh5jw6 & Ei5jw6);
assign Ei5jw6 = (~(Yxf7z6[18] & Pw0jw6));
assign Xh5jw6 = (~(Hz0jw6 & Kxb7z6[15]));
assign Tf5jw6 = (Li5jw6 & Si5jw6);
assign Si5jw6 = (Zi5jw6 & Gj5jw6);
assign Gj5jw6 = (~(J01jw6 & Onf7z6[31]));
assign Zi5jw6 = (Nj5jw6 & Uj5jw6);
assign Uj5jw6 = (~(Oz0jw6 & Fhc7z6[15]));
assign Nj5jw6 = (~(Onf7z6[15] & My0jw6));
assign Li5jw6 = (Bk5jw6 & Ik5jw6);
assign Ik5jw6 = (Pk5jw6 | Dx0jw6);
assign Bk5jw6 = (~(Q01jw6 & Alf7z6[15]));
assign F7nnv6 = (~(Wk5jw6 ^ Tennv6));
assign Wk5jw6 = (~(Dl5jw6 & Kl5jw6));
assign Kl5jw6 = (~(Yxf7z6[15] & Gbziw6));
assign Dl5jw6 = (~(Kxb7z6[15] & Nbziw6));
assign A25jw6 = (Rl5jw6 & Yl5jw6);
assign Yl5jw6 = (~(Pw9ov6 & Kxb7z6[15]));
assign Rl5jw6 = (Fm5jw6 & Mm5jw6);
assign Mm5jw6 = (~(Kx9ov6 & vis_pc_o[15]));
assign Fm5jw6 = (~(Gli7z6[15] & Rx9ov6));
assign X8z7v6 = (~(Tm5jw6 & An5jw6));
assign An5jw6 = (~(Eji7z6[16] & C3yiw6));
assign Tm5jw6 = (Hn5jw6 & On5jw6);
assign On5jw6 = (~(Bhi7z6[16] & X3yiw6));
assign Hn5jw6 = (~(E4yiw6 & vis_pc_o[16]));
assign Q8z7v6 = (~(Vn5jw6 & Co5jw6));
assign Co5jw6 = (~(Eji7z6[17] & C3yiw6));
assign Vn5jw6 = (Jo5jw6 & Qo5jw6);
assign Qo5jw6 = (~(Bhi7z6[17] & X3yiw6));
assign Jo5jw6 = (~(E4yiw6 & vis_pc_o[17]));
assign J8z7v6 = (~(Xo5jw6 & Ep5jw6));
assign Ep5jw6 = (~(Eji7z6[18] & C3yiw6));
assign Xo5jw6 = (Lp5jw6 & Sp5jw6);
assign Sp5jw6 = (~(Bhi7z6[18] & X3yiw6));
assign Lp5jw6 = (~(E4yiw6 & vis_pc_o[18]));
assign C8z7v6 = (~(Zp5jw6 & Gq5jw6));
assign Gq5jw6 = (Nq5jw6 & Uq5jw6);
assign Uq5jw6 = (Eu9ov6 | Br5jw6);
assign Nq5jw6 = (Ir5jw6 & Pr5jw6);
assign Pr5jw6 = (~(Gv9ov6 & Zqxiw6));
assign Zqxiw6 = (Spyiw6 ? Yw97z6 : Gli7z6[18]);
assign Ir5jw6 = (~(Uv9ov6 & Yw97z6));
assign Yw97z6 = (~(Wr5jw6 & Ds5jw6));
assign Ds5jw6 = (~(Nqyiw6 & Kuynv6));
assign Wr5jw6 = (Ks5jw6 & Rs5jw6);
assign Rs5jw6 = (~(Pdc7z6[18] & Ouyiw6));
assign Ks5jw6 = (~(Vuyiw6 & Ys5jw6));
assign Ys5jw6 = (~(Ft5jw6 & Mt5jw6));
assign Mt5jw6 = (Tt5jw6 & Au5jw6);
assign Au5jw6 = (Hu5jw6 & Ou5jw6);
assign Ou5jw6 = (Vu5jw6 & Cv5jw6);
assign Cv5jw6 = (~(Jv5jw6 & Uxyiw6));
assign Jv5jw6 = (Kxb7z6[18] & Qv5jw6);
assign Vu5jw6 = (~(Xv5jw6 & Ew5jw6));
assign Xv5jw6 = (~(Lw5jw6 & Quziw6));
assign Lw5jw6 = (Sw5jw6 & Zw5jw6);
assign Zw5jw6 = (Qv5jw6 | Ninnv6);
assign Qv5jw6 = (Gx5jw6 | Rje7z6[18]);
assign Sw5jw6 = (~(Ofnnv6 & Gx5jw6));
assign Hu5jw6 = (Nx5jw6 & Ux5jw6);
assign Ux5jw6 = (~(J73ov6 & Hk3ov6));
assign Hk3ov6 = (~(Ur4jw6 ^ Dte7z6[1]));
assign Ur4jw6 = (T3cdt6 ? Xlohw6 : Z04ov6);
assign Xlohw6 = (!V1c7z6[10]);
assign Nx5jw6 = (~(R6ziw6 & Db3ov6));
assign Tt5jw6 = (By5jw6 & Iy5jw6);
assign Iy5jw6 = (Py5jw6 & Wy5jw6);
assign Wy5jw6 = (~(F7ziw6 & Vd3ov6));
assign Py5jw6 = (~(T0ziw6 & Rje7z6[18]));
assign By5jw6 = (Dz5jw6 & Kz5jw6);
assign Kz5jw6 = (Ryfov6 | Rz5jw6);
assign Dz5jw6 = (~(L0g7z6[18] & J2ziw6));
assign Ft5jw6 = (Yz5jw6 & F06jw6);
assign F06jw6 = (M06jw6 & T06jw6);
assign T06jw6 = (A16jw6 & H16jw6);
assign H16jw6 = (~(Cqf7z6[2] & Q2ziw6));
assign A16jw6 = (~(O1ziw6 & L0g7z6[2]));
assign M06jw6 = (O16jw6 & V16jw6);
assign V16jw6 = (~(U4ziw6 & V1c7z6[18]));
assign O16jw6 = (~(Z3ziw6 & Fhc7z6[13]));
assign Yz5jw6 = (C26jw6 & Xt2ov6);
assign Xt2ov6 = (J26jw6 & Q26jw6);
assign Q26jw6 = (~(X26jw6 & P5nnv6));
assign X26jw6 = (~(W5nnv6 | Icziw6));
assign J26jw6 = (~(E36jw6 & Ubziw6));
assign E36jw6 = (~(P5nnv6 ^ W5nnv6));
assign W5nnv6 = (L36jw6 ^ Mennv6);
assign L36jw6 = (~(S36jw6 & Z36jw6));
assign Z36jw6 = (G46jw6 & N46jw6);
assign N46jw6 = (U46jw6 & B56jw6);
assign B56jw6 = (~(Yxf7z6[20] & Su0jw6));
assign U46jw6 = (I56jw6 & P56jw6);
assign P56jw6 = (~(Yxf7z6[18] & Nv0jw6));
assign I56jw6 = (~(Yxf7z6[19] & Uv0jw6));
assign G46jw6 = (W56jw6 & D66jw6);
assign D66jw6 = (~(Yxf7z6[21] & Pw0jw6));
assign W56jw6 = (~(K66jw6 & Rdziw6));
assign S36jw6 = (R66jw6 & Y66jw6);
assign Y66jw6 = (F76jw6 & M76jw6);
assign M76jw6 = (~(Onf7z6[18] & My0jw6));
assign F76jw6 = (T76jw6 & A86jw6);
assign A86jw6 = (~(Hz0jw6 & Kxb7z6[18]));
assign T76jw6 = (~(Oz0jw6 & Fhc7z6[18]));
assign R66jw6 = (H86jw6 & O86jw6);
assign O86jw6 = (~(Alf7z6[2] & J01jw6));
assign H86jw6 = (~(Alf7z6[18] & Q01jw6));
assign P5nnv6 = (~(V86jw6 ^ Tennv6));
assign V86jw6 = (~(C96jw6 & J96jw6));
assign J96jw6 = (~(Yxf7z6[2] & Laziw6));
assign C96jw6 = (Q96jw6 & X96jw6);
assign X96jw6 = (~(Yxf7z6[18] & Gbziw6));
assign Q96jw6 = (~(Kxb7z6[18] & Nbziw6));
assign C26jw6 = (T7ziw6 & Ea6jw6);
assign Ea6jw6 = (~(Zkldt6 & Oztiw6));
assign Zp5jw6 = (La6jw6 & Sa6jw6);
assign Sa6jw6 = (~(Pw9ov6 & Kxb7z6[18]));
assign La6jw6 = (Za6jw6 & Gb6jw6);
assign Gb6jw6 = (~(Kx9ov6 & vis_pc_o[18]));
assign Za6jw6 = (~(Gli7z6[18] & Rx9ov6));
assign V7z7v6 = (~(Nb6jw6 & Ub6jw6));
assign Ub6jw6 = (~(Eji7z6[19] & C3yiw6));
assign Nb6jw6 = (Bc6jw6 & Ic6jw6);
assign Ic6jw6 = (~(Bhi7z6[19] & X3yiw6));
assign Bc6jw6 = (~(E4yiw6 & vis_pc_o[19]));
assign O7z7v6 = (~(Pc6jw6 & Wc6jw6));
assign Wc6jw6 = (~(Eji7z6[20] & C3yiw6));
assign Pc6jw6 = (Dd6jw6 & Kd6jw6);
assign Kd6jw6 = (~(Bhi7z6[20] & X3yiw6));
assign Dd6jw6 = (~(E4yiw6 & vis_pc_o[20]));
assign H7z7v6 = (~(Rd6jw6 & Yd6jw6));
assign Yd6jw6 = (~(Eji7z6[21] & C3yiw6));
assign Rd6jw6 = (Fe6jw6 & Me6jw6);
assign Me6jw6 = (~(Bhi7z6[21] & X3yiw6));
assign Fe6jw6 = (~(E4yiw6 & vis_pc_o[21]));
assign A7z7v6 = (~(Te6jw6 & Af6jw6));
assign Af6jw6 = (~(Eji7z6[22] & C3yiw6));
assign Te6jw6 = (Hf6jw6 & Of6jw6);
assign Of6jw6 = (~(Bhi7z6[22] & X3yiw6));
assign Hf6jw6 = (~(E4yiw6 & vis_pc_o[22]));
assign T6z7v6 = (~(Vf6jw6 & Cg6jw6));
assign Cg6jw6 = (~(Eji7z6[23] & C3yiw6));
assign Vf6jw6 = (Jg6jw6 & Qg6jw6);
assign Qg6jw6 = (~(Bhi7z6[23] & X3yiw6));
assign Jg6jw6 = (~(E4yiw6 & vis_pc_o[23]));
assign M6z7v6 = (~(Xg6jw6 & Eh6jw6));
assign Eh6jw6 = (~(Eji7z6[24] & C3yiw6));
assign Xg6jw6 = (Lh6jw6 & Sh6jw6);
assign Sh6jw6 = (~(Bhi7z6[24] & X3yiw6));
assign Lh6jw6 = (~(E4yiw6 & vis_pc_o[24]));
assign F6z7v6 = (~(Zh6jw6 & Gi6jw6));
assign Gi6jw6 = (~(Eji7z6[25] & C3yiw6));
assign Zh6jw6 = (Ni6jw6 & Ui6jw6);
assign Ui6jw6 = (~(Bhi7z6[25] & X3yiw6));
assign Ni6jw6 = (~(E4yiw6 & vis_pc_o[25]));
assign Y5z7v6 = (~(Bj6jw6 & Ij6jw6));
assign Ij6jw6 = (Pj6jw6 & Wj6jw6);
assign Wj6jw6 = (Eu9ov6 | Dk6jw6);
assign Pj6jw6 = (Kk6jw6 & Rk6jw6);
assign Rk6jw6 = (~(Gv9ov6 & R7yiw6));
assign Kk6jw6 = (~(Uv9ov6 & Ox97z6));
assign Bj6jw6 = (Yk6jw6 & Fl6jw6);
assign Fl6jw6 = (~(Pw9ov6 & Kxb7z6[25]));
assign Yk6jw6 = (Ml6jw6 & Tl6jw6);
assign Tl6jw6 = (~(Kx9ov6 & vis_pc_o[25]));
assign Ml6jw6 = (~(Gli7z6[25] & Rx9ov6));
assign R5z7v6 = (~(Am6jw6 & Hm6jw6));
assign Hm6jw6 = (Om6jw6 & Vm6jw6);
assign Vm6jw6 = (~(H02ov6 & Ox97z6));
assign Om6jw6 = (Cn6jw6 & Jn6jw6);
assign Jn6jw6 = (C12ov6 | Kvjnv6);
assign Kvjnv6 = (Qn6jw6 & Xn6jw6);
assign Xn6jw6 = (Eo6jw6 & Lo6jw6);
assign Lo6jw6 = (So6jw6 & Zo6jw6);
assign Zo6jw6 = (Gp6jw6 & Np6jw6);
assign Np6jw6 = (~(vis_psp_o[25] & N32ov6));
assign Gp6jw6 = (~(U32ov6 & Pic7z6[25]));
assign So6jw6 = (Up6jw6 & Bq6jw6);
assign Bq6jw6 = (~(vis_msp_o[25] & P42ov6));
assign Up6jw6 = (~(vis_r12_o[25] & W42ov6));
assign Eo6jw6 = (Iq6jw6 & Pq6jw6);
assign Pq6jw6 = (Wq6jw6 & Dr6jw6);
assign Dr6jw6 = (~(vis_r11_o[25] & F62ov6));
assign Wq6jw6 = (~(vis_r10_o[25] & M62ov6));
assign Iq6jw6 = (Kr6jw6 & Rr6jw6);
assign Rr6jw6 = (~(vis_r9_o[25] & H72ov6));
assign Kr6jw6 = (~(vis_r8_o[25] & O72ov6));
assign Qn6jw6 = (Yr6jw6 & Fs6jw6);
assign Fs6jw6 = (Ms6jw6 & Ts6jw6);
assign Ts6jw6 = (At6jw6 & Ht6jw6);
assign Ht6jw6 = (~(vis_r7_o[25] & L92ov6));
assign At6jw6 = (~(vis_r6_o[25] & S92ov6));
assign Ms6jw6 = (Ot6jw6 & Vt6jw6);
assign Vt6jw6 = (~(vis_r5_o[25] & Na2ov6));
assign Ot6jw6 = (~(vis_r4_o[25] & Ua2ov6));
assign Yr6jw6 = (Cu6jw6 & Ju6jw6);
assign Ju6jw6 = (Qu6jw6 & Xu6jw6);
assign Xu6jw6 = (~(vis_r3_o[25] & Dc2ov6));
assign Qu6jw6 = (~(vis_r2_o[25] & Kc2ov6));
assign Cu6jw6 = (Ev6jw6 & Lv6jw6);
assign Lv6jw6 = (~(vis_r1_o[25] & Fd2ov6));
assign Ev6jw6 = (~(vis_r0_o[25] & Md2ov6));
assign Cn6jw6 = (~(Td2ov6 & R7yiw6));
assign R7yiw6 = (Spyiw6 ? Ox97z6 : Gli7z6[25]);
assign Ox97z6 = (~(Sv6jw6 & Zv6jw6));
assign Zv6jw6 = (~(Nqyiw6 & Xyxnv6));
assign Sv6jw6 = (Gw6jw6 & Nw6jw6);
assign Nw6jw6 = (~(Pdc7z6[25] & Ouyiw6));
assign Gw6jw6 = (~(Vuyiw6 & Uw6jw6));
assign Uw6jw6 = (~(Bx6jw6 & Ix6jw6));
assign Ix6jw6 = (Px6jw6 & Wx6jw6);
assign Wx6jw6 = (Dy6jw6 & Ky6jw6);
assign Ky6jw6 = (Ry6jw6 & Yy6jw6);
assign Yy6jw6 = (~(Fz6jw6 & Uxyiw6));
assign Fz6jw6 = (Kxb7z6[25] & Mz6jw6);
assign Ry6jw6 = (~(Tz6jw6 & A07jw6));
assign Tz6jw6 = (~(H07jw6 & Quziw6));
assign H07jw6 = (O07jw6 & V07jw6);
assign V07jw6 = (Mz6jw6 | Ninnv6);
assign Mz6jw6 = (~(C17jw6 & J17jw6));
assign C17jw6 = (!Rje7z6[25]);
assign O07jw6 = (J17jw6 | Evziw6);
assign Dy6jw6 = (Q17jw6 & X17jw6);
assign X17jw6 = (J17jw6 | Ryfov6);
assign Q17jw6 = (~(J73ov6 & Io3ov6));
assign Px6jw6 = (E27jw6 & L27jw6);
assign L27jw6 = (S27jw6 & Z27jw6);
assign Z27jw6 = (Sf3ov6 | U93ov6);
assign S27jw6 = (~(R6ziw6 & Ia3ov6));
assign E27jw6 = (G37jw6 & N37jw6);
assign N37jw6 = (~(T0ziw6 & Rje7z6[25]));
assign G37jw6 = (~(L0g7z6[25] & J2ziw6));
assign Bx6jw6 = (U37jw6 & B47jw6);
assign B47jw6 = (I47jw6 & P47jw6);
assign P47jw6 = (W47jw6 & D57jw6);
assign D57jw6 = (~(Cqf7z6[9] & Q2ziw6));
assign W47jw6 = (~(L0g7z6[9] & O1ziw6));
assign I47jw6 = (K57jw6 & R57jw6);
assign R57jw6 = (~(U4ziw6 & V1c7z6[25]));
assign K57jw6 = (~(Z3ziw6 & Fhc7z6[6]));
assign U37jw6 = (Y57jw6 & Su2ov6);
assign Su2ov6 = (F67jw6 & M67jw6);
assign M67jw6 = (~(T67jw6 & H1nnv6));
assign T67jw6 = (~(O1nnv6 | Icziw6));
assign F67jw6 = (~(A77jw6 & Ubziw6));
assign A77jw6 = (~(H1nnv6 ^ O1nnv6));
assign O1nnv6 = (H77jw6 ^ Mennv6);
assign H77jw6 = (~(O77jw6 & V77jw6));
assign V77jw6 = (C87jw6 & J87jw6);
assign J87jw6 = (Q87jw6 & X87jw6);
assign X87jw6 = (~(Yxf7z6[27] & Su0jw6));
assign Q87jw6 = (E97jw6 & L97jw6);
assign L97jw6 = (~(Yxf7z6[25] & Nv0jw6));
assign E97jw6 = (~(Yxf7z6[26] & Uv0jw6));
assign C87jw6 = (S97jw6 & Z97jw6);
assign Z97jw6 = (~(Pw0jw6 & Yxf7z6[28]));
assign S97jw6 = (~(Ga7jw6 & Rdziw6));
assign O77jw6 = (Na7jw6 & Ua7jw6);
assign Ua7jw6 = (Bb7jw6 & Ib7jw6);
assign Ib7jw6 = (~(Onf7z6[25] & My0jw6));
assign Bb7jw6 = (Pb7jw6 & Wb7jw6);
assign Wb7jw6 = (~(Hz0jw6 & Kxb7z6[25]));
assign Pb7jw6 = (~(Oz0jw6 & Fhc7z6[25]));
assign Na7jw6 = (Dc7jw6 & Kc7jw6);
assign Kc7jw6 = (~(Alf7z6[9] & J01jw6));
assign Dc7jw6 = (~(Alf7z6[25] & Q01jw6));
assign H1nnv6 = (~(Rc7jw6 ^ Tennv6));
assign Rc7jw6 = (~(Yc7jw6 & Fd7jw6));
assign Fd7jw6 = (~(Yxf7z6[9] & Laziw6));
assign Yc7jw6 = (Md7jw6 & Td7jw6);
assign Td7jw6 = (~(Yxf7z6[25] & Gbziw6));
assign Md7jw6 = (~(Kxb7z6[25] & Nbziw6));
assign Y57jw6 = (T7ziw6 & Ae7jw6);
assign Ae7jw6 = (~(E6ldt6 & Oztiw6));
assign Am6jw6 = (He7jw6 & Oe7jw6);
assign Oe7jw6 = (~(Ve2ov6 & vis_pc_o[25]));
assign He7jw6 = (~(Fhc7z6[25] & Cf2ov6));
assign K5z7v6 = (~(Ve7jw6 & Cf7jw6));
assign Cf7jw6 = (Jf7jw6 & Qf7jw6);
assign Qf7jw6 = (Eu9ov6 | Xf7jw6);
assign Jf7jw6 = (Eg7jw6 & Lg7jw6);
assign Lg7jw6 = (~(Gv9ov6 & Y7yiw6));
assign Eg7jw6 = (~(Uv9ov6 & Wx97z6));
assign Ve7jw6 = (Sg7jw6 & Zg7jw6);
assign Zg7jw6 = (~(Pw9ov6 & Kxb7z6[24]));
assign Sg7jw6 = (Gh7jw6 & Nh7jw6);
assign Nh7jw6 = (~(Kx9ov6 & vis_pc_o[24]));
assign Gh7jw6 = (~(Gli7z6[24] & Rx9ov6));
assign D5z7v6 = (~(Uh7jw6 & Bi7jw6));
assign Bi7jw6 = (Ii7jw6 & Pi7jw6);
assign Pi7jw6 = (~(H02ov6 & Wx97z6));
assign Ii7jw6 = (Wi7jw6 & Dj7jw6);
assign Dj7jw6 = (C12ov6 | Axjnv6);
assign Axjnv6 = (Kj7jw6 & Rj7jw6);
assign Rj7jw6 = (Yj7jw6 & Fk7jw6);
assign Fk7jw6 = (Mk7jw6 & Tk7jw6);
assign Tk7jw6 = (Al7jw6 & Hl7jw6);
assign Hl7jw6 = (~(vis_psp_o[24] & N32ov6));
assign Al7jw6 = (~(U32ov6 & Pic7z6[24]));
assign Mk7jw6 = (Ol7jw6 & Vl7jw6);
assign Vl7jw6 = (~(vis_msp_o[24] & P42ov6));
assign Ol7jw6 = (~(vis_r12_o[24] & W42ov6));
assign Yj7jw6 = (Cm7jw6 & Jm7jw6);
assign Jm7jw6 = (Qm7jw6 & Xm7jw6);
assign Xm7jw6 = (~(vis_r11_o[24] & F62ov6));
assign Qm7jw6 = (~(vis_r10_o[24] & M62ov6));
assign Cm7jw6 = (En7jw6 & Ln7jw6);
assign Ln7jw6 = (~(vis_r9_o[24] & H72ov6));
assign En7jw6 = (~(vis_r8_o[24] & O72ov6));
assign Kj7jw6 = (Sn7jw6 & Zn7jw6);
assign Zn7jw6 = (Go7jw6 & No7jw6);
assign No7jw6 = (Uo7jw6 & Bp7jw6);
assign Bp7jw6 = (~(vis_r7_o[24] & L92ov6));
assign Uo7jw6 = (~(vis_r6_o[24] & S92ov6));
assign Go7jw6 = (Ip7jw6 & Pp7jw6);
assign Pp7jw6 = (~(vis_r5_o[24] & Na2ov6));
assign Ip7jw6 = (~(vis_r4_o[24] & Ua2ov6));
assign Sn7jw6 = (Wp7jw6 & Dq7jw6);
assign Dq7jw6 = (Kq7jw6 & Rq7jw6);
assign Rq7jw6 = (~(vis_r3_o[24] & Dc2ov6));
assign Kq7jw6 = (~(vis_r2_o[24] & Kc2ov6));
assign Wp7jw6 = (Yq7jw6 & Fr7jw6);
assign Fr7jw6 = (~(vis_r1_o[24] & Fd2ov6));
assign Yq7jw6 = (~(vis_r0_o[24] & Md2ov6));
assign Wi7jw6 = (~(Td2ov6 & Y7yiw6));
assign Y7yiw6 = (Spyiw6 ? Wx97z6 : Gli7z6[24]);
assign Wx97z6 = (~(Mr7jw6 & Tr7jw6));
assign Tr7jw6 = (~(Nqyiw6 & M3ynv6));
assign Mr7jw6 = (As7jw6 & Hs7jw6);
assign Hs7jw6 = (~(Pdc7z6[24] & Ouyiw6));
assign As7jw6 = (~(Vuyiw6 & Os7jw6));
assign Os7jw6 = (~(Vs7jw6 & Ct7jw6));
assign Ct7jw6 = (Jt7jw6 & Qt7jw6);
assign Qt7jw6 = (Xt7jw6 & Eu7jw6);
assign Eu7jw6 = (Lu7jw6 & Su7jw6);
assign Su7jw6 = (~(Zu7jw6 & Uxyiw6));
assign Zu7jw6 = (Kxb7z6[24] & Gv7jw6);
assign Lu7jw6 = (~(Nv7jw6 & T9kov6));
assign Nv7jw6 = (~(Uv7jw6 & Quziw6));
assign Uv7jw6 = (Bw7jw6 & Iw7jw6);
assign Iw7jw6 = (Gv7jw6 | Ninnv6);
assign Gv7jw6 = (Rje7z6[24] | Pw7jw6);
assign Bw7jw6 = (~(Ofnnv6 & Pw7jw6));
assign Xt7jw6 = (Ww7jw6 & Dx7jw6);
assign Dx7jw6 = (~(J73ov6 & Bo3ov6));
assign Bo3ov6 = (~(Ww0jw6 ^ Dte7z6[1]));
assign Ww0jw6 = (T3cdt6 ? J6jnv6 : C64ov6);
assign Ww7jw6 = (~(F7ziw6 & Pa3ov6));
assign Jt7jw6 = (Kx7jw6 & Rx7jw6);
assign Rx7jw6 = (Yx7jw6 & Fy7jw6);
assign Fy7jw6 = (Zf3ov6 | Ba3ov6);
assign Yx7jw6 = (~(T0ziw6 & Rje7z6[24]));
assign Kx7jw6 = (My7jw6 & Ty7jw6);
assign Ty7jw6 = (Ryfov6 | Az7jw6);
assign My7jw6 = (~(L0g7z6[24] & J2ziw6));
assign Vs7jw6 = (Hz7jw6 & Oz7jw6);
assign Oz7jw6 = (Vz7jw6 & C08jw6);
assign C08jw6 = (J08jw6 & Q08jw6);
assign Q08jw6 = (~(Cqf7z6[8] & Q2ziw6));
assign J08jw6 = (~(L0g7z6[8] & O1ziw6));
assign Vz7jw6 = (X08jw6 & E18jw6);
assign E18jw6 = (~(U4ziw6 & V1c7z6[24]));
assign X08jw6 = (~(Z3ziw6 & Fhc7z6[7]));
assign Hz7jw6 = (L18jw6 & Lu2ov6);
assign Lu2ov6 = (S18jw6 & Z18jw6);
assign Z18jw6 = (~(G28jw6 & V1nnv6));
assign G28jw6 = (~(C2nnv6 | Icziw6));
assign S18jw6 = (~(N28jw6 & Ubziw6));
assign N28jw6 = (~(V1nnv6 ^ C2nnv6));
assign C2nnv6 = (U28jw6 ^ Mennv6);
assign U28jw6 = (~(B38jw6 & I38jw6));
assign I38jw6 = (P38jw6 & W38jw6);
assign W38jw6 = (D48jw6 & K48jw6);
assign K48jw6 = (~(Yxf7z6[26] & Su0jw6));
assign D48jw6 = (R48jw6 & Y48jw6);
assign Y48jw6 = (~(Yxf7z6[24] & Nv0jw6));
assign R48jw6 = (~(Yxf7z6[25] & Uv0jw6));
assign P38jw6 = (F58jw6 & M58jw6);
assign M58jw6 = (~(Yxf7z6[27] & Pw0jw6));
assign F58jw6 = (~(T58jw6 & Rdziw6));
assign B38jw6 = (A68jw6 & H68jw6);
assign H68jw6 = (O68jw6 & V68jw6);
assign V68jw6 = (~(Onf7z6[24] & My0jw6));
assign O68jw6 = (C78jw6 & J78jw6);
assign J78jw6 = (~(Hz0jw6 & Kxb7z6[24]));
assign C78jw6 = (~(Oz0jw6 & Fhc7z6[24]));
assign A68jw6 = (Q78jw6 & X78jw6);
assign X78jw6 = (~(Alf7z6[8] & J01jw6));
assign Q78jw6 = (~(Alf7z6[24] & Q01jw6));
assign V1nnv6 = (~(E88jw6 ^ Tennv6));
assign E88jw6 = (~(L88jw6 & S88jw6));
assign S88jw6 = (~(Yxf7z6[8] & Laziw6));
assign L88jw6 = (Z88jw6 & G98jw6);
assign G98jw6 = (~(Yxf7z6[24] & Gbziw6));
assign Z88jw6 = (~(Kxb7z6[24] & Nbziw6));
assign L18jw6 = (T7ziw6 & N98jw6);
assign N98jw6 = (~(H8ldt6 & Oztiw6));
assign Uh7jw6 = (U98jw6 & Ba8jw6);
assign Ba8jw6 = (~(Ve2ov6 & vis_pc_o[24]));
assign U98jw6 = (~(Fhc7z6[24] & Cf2ov6));
assign W4z7v6 = (~(Ia8jw6 & Pa8jw6));
assign Pa8jw6 = (Wa8jw6 & Db8jw6);
assign Db8jw6 = (Eu9ov6 | Kb8jw6);
assign Wa8jw6 = (Rb8jw6 & Yb8jw6);
assign Yb8jw6 = (~(Gv9ov6 & V9yiw6));
assign Rb8jw6 = (~(Uv9ov6 & A0a7z6));
assign Ia8jw6 = (Fc8jw6 & Mc8jw6);
assign Mc8jw6 = (~(Pw9ov6 & Kxb7z6[16]));
assign Fc8jw6 = (Tc8jw6 & Ad8jw6);
assign Ad8jw6 = (~(Kx9ov6 & vis_pc_o[16]));
assign Tc8jw6 = (~(Gli7z6[16] & Rx9ov6));
assign P4z7v6 = (~(Hd8jw6 & Od8jw6));
assign Od8jw6 = (Vd8jw6 & Ce8jw6);
assign Ce8jw6 = (~(H02ov6 & A0a7z6));
assign Vd8jw6 = (Je8jw6 & Qe8jw6);
assign Qe8jw6 = (C12ov6 | Ccknv6);
assign Ccknv6 = (Xe8jw6 & Ef8jw6);
assign Ef8jw6 = (Lf8jw6 & Sf8jw6);
assign Sf8jw6 = (Zf8jw6 & Gg8jw6);
assign Gg8jw6 = (Ng8jw6 & Ug8jw6);
assign Ug8jw6 = (~(vis_psp_o[16] & N32ov6));
assign Ng8jw6 = (~(U32ov6 & Pic7z6[16]));
assign Zf8jw6 = (Bh8jw6 & Ih8jw6);
assign Ih8jw6 = (~(vis_msp_o[16] & P42ov6));
assign Bh8jw6 = (~(vis_r12_o[16] & W42ov6));
assign Lf8jw6 = (Ph8jw6 & Wh8jw6);
assign Wh8jw6 = (Di8jw6 & Ki8jw6);
assign Ki8jw6 = (~(vis_r11_o[16] & F62ov6));
assign Di8jw6 = (~(vis_r10_o[16] & M62ov6));
assign Ph8jw6 = (Ri8jw6 & Yi8jw6);
assign Yi8jw6 = (~(vis_r9_o[16] & H72ov6));
assign Ri8jw6 = (~(vis_r8_o[16] & O72ov6));
assign Xe8jw6 = (Fj8jw6 & Mj8jw6);
assign Mj8jw6 = (Tj8jw6 & Ak8jw6);
assign Ak8jw6 = (Hk8jw6 & Ok8jw6);
assign Ok8jw6 = (~(vis_r7_o[16] & L92ov6));
assign Hk8jw6 = (~(vis_r6_o[16] & S92ov6));
assign Tj8jw6 = (Vk8jw6 & Cl8jw6);
assign Cl8jw6 = (~(vis_r5_o[16] & Na2ov6));
assign Vk8jw6 = (~(vis_r4_o[16] & Ua2ov6));
assign Fj8jw6 = (Jl8jw6 & Ql8jw6);
assign Ql8jw6 = (Xl8jw6 & Em8jw6);
assign Em8jw6 = (~(vis_r3_o[16] & Dc2ov6));
assign Xl8jw6 = (~(vis_r2_o[16] & Kc2ov6));
assign Jl8jw6 = (Lm8jw6 & Sm8jw6);
assign Sm8jw6 = (~(vis_r1_o[16] & Fd2ov6));
assign Lm8jw6 = (~(vis_r0_o[16] & Md2ov6));
assign Je8jw6 = (~(Td2ov6 & V9yiw6));
assign V9yiw6 = (Spyiw6 ? A0a7z6 : Gli7z6[16]);
assign A0a7z6 = (~(Zm8jw6 & Gn8jw6));
assign Gn8jw6 = (~(Nqyiw6 & O3znv6));
assign Zm8jw6 = (Nn8jw6 & Un8jw6);
assign Un8jw6 = (~(Pdc7z6[16] & Ouyiw6));
assign Nn8jw6 = (~(Vuyiw6 & Bo8jw6));
assign Bo8jw6 = (~(Io8jw6 & Po8jw6));
assign Po8jw6 = (Wo8jw6 & Dp8jw6);
assign Dp8jw6 = (Kp8jw6 & Rp8jw6);
assign Rp8jw6 = (Yp8jw6 & Fq8jw6);
assign Fq8jw6 = (~(Mq8jw6 & Uxyiw6));
assign Mq8jw6 = (Kxb7z6[16] & Tq8jw6);
assign Yp8jw6 = (~(Ar8jw6 & Hr8jw6));
assign Ar8jw6 = (~(Or8jw6 & Quziw6));
assign Or8jw6 = (Vr8jw6 & Cs8jw6);
assign Cs8jw6 = (Tq8jw6 | Ninnv6);
assign Tq8jw6 = (Rje7z6[16] | Js8jw6);
assign Vr8jw6 = (~(Ofnnv6 & Js8jw6));
assign Kp8jw6 = (Qs8jw6 & Xs8jw6);
assign Xs8jw6 = (~(R6ziw6 & Pa3ov6));
assign Pa3ov6 = (T58jw6 ^ Dte7z6[1]);
assign T58jw6 = (T3cdt6 ? V1c7z6[24] : T9kov6);
assign Qs8jw6 = (~(J73ov6 & Tj3ov6));
assign Tj3ov6 = (~(E54jw6 ^ Dte7z6[1]));
assign E54jw6 = (T3cdt6 ? E0phw6 : Vy3ov6);
assign Wo8jw6 = (Et8jw6 & Lt8jw6);
assign Lt8jw6 = (St8jw6 & Zt8jw6);
assign Zt8jw6 = (Sf3ov6 | Ba3ov6);
assign Ba3ov6 = (Gu8jw6 ^ Nu8jw6);
assign St8jw6 = (~(T0ziw6 & Rje7z6[16]));
assign Et8jw6 = (Uu8jw6 & Bv8jw6);
assign Bv8jw6 = (Ryfov6 | Iv8jw6);
assign Uu8jw6 = (~(L0g7z6[16] & J2ziw6));
assign Io8jw6 = (Pv8jw6 & Wv8jw6);
assign Wv8jw6 = (Dw8jw6 & Kw8jw6);
assign Kw8jw6 = (Rw8jw6 & Yw8jw6);
assign Yw8jw6 = (~(Cqf7z6[0] & Q2ziw6));
assign Rw8jw6 = (~(L0g7z6[0] & O1ziw6));
assign Dw8jw6 = (Fx8jw6 & Mx8jw6);
assign Mx8jw6 = (~(U4ziw6 & V1c7z6[16]));
assign Fx8jw6 = (~(Z3ziw6 & Fhc7z6[15]));
assign Pv8jw6 = (Tx8jw6 & Uv2ov6);
assign Uv2ov6 = (Ay8jw6 & Hy8jw6);
assign Hy8jw6 = (~(Oy8jw6 & R6nnv6));
assign Oy8jw6 = (~(Y6nnv6 | Icziw6));
assign Ay8jw6 = (~(Vy8jw6 & Ubziw6));
assign Vy8jw6 = (~(R6nnv6 ^ Y6nnv6));
assign Y6nnv6 = (Cz8jw6 ^ Mennv6);
assign Cz8jw6 = (~(Jz8jw6 & Qz8jw6));
assign Qz8jw6 = (Xz8jw6 & E09jw6);
assign E09jw6 = (L09jw6 & S09jw6);
assign S09jw6 = (~(Yxf7z6[18] & Su0jw6));
assign L09jw6 = (Z09jw6 & G19jw6);
assign G19jw6 = (~(Yxf7z6[16] & Nv0jw6));
assign Z09jw6 = (~(Yxf7z6[17] & Uv0jw6));
assign Xz8jw6 = (N19jw6 & U19jw6);
assign U19jw6 = (~(Yxf7z6[19] & Pw0jw6));
assign N19jw6 = (~(Gu8jw6 & Rdziw6));
assign Gu8jw6 = (T3cdt6 ? V1c7z6[16] : Hr8jw6);
assign Jz8jw6 = (B29jw6 & I29jw6);
assign I29jw6 = (P29jw6 & W29jw6);
assign W29jw6 = (~(Onf7z6[16] & My0jw6));
assign P29jw6 = (D39jw6 & K39jw6);
assign K39jw6 = (~(Hz0jw6 & Kxb7z6[16]));
assign D39jw6 = (~(Oz0jw6 & Fhc7z6[16]));
assign B29jw6 = (R39jw6 & Y39jw6);
assign Y39jw6 = (~(Alf7z6[0] & J01jw6));
assign R39jw6 = (~(Alf7z6[16] & Q01jw6));
assign R6nnv6 = (~(F49jw6 ^ Tennv6));
assign F49jw6 = (~(M49jw6 & T49jw6));
assign T49jw6 = (~(Yxf7z6[0] & Laziw6));
assign M49jw6 = (A59jw6 & H59jw6);
assign H59jw6 = (~(Yxf7z6[16] & Gbziw6));
assign A59jw6 = (~(Kxb7z6[16] & Nbziw6));
assign Tx8jw6 = (T7ziw6 & O59jw6);
assign O59jw6 = (~(Fpldt6 & Oztiw6));
assign Hd8jw6 = (V59jw6 & C69jw6);
assign C69jw6 = (~(Ve2ov6 & vis_pc_o[16]));
assign V59jw6 = (~(Fhc7z6[16] & Cf2ov6));
assign I4z7v6 = (~(J69jw6 & Q69jw6));
assign Q69jw6 = (X69jw6 & E79jw6);
assign E79jw6 = (Eu9ov6 | L79jw6);
assign X69jw6 = (S79jw6 & Z79jw6);
assign Z79jw6 = (~(Gv9ov6 & Lbyiw6));
assign S79jw6 = (~(Uv9ov6 & O1a7z6));
assign J69jw6 = (G89jw6 & N89jw6);
assign N89jw6 = (~(Pw9ov6 & Kxb7z6[9]));
assign G89jw6 = (U89jw6 & B99jw6);
assign B99jw6 = (~(Kx9ov6 & vis_pc_o[9]));
assign U89jw6 = (~(Gli7z6[9] & Rx9ov6));
assign B4z7v6 = (~(I99jw6 & P99jw6));
assign P99jw6 = (W99jw6 & Da9jw6);
assign Da9jw6 = (~(H02ov6 & O1a7z6));
assign W99jw6 = (Ka9jw6 & Ra9jw6);
assign Ra9jw6 = (C12ov6 | U8jnv6);
assign U8jnv6 = (Ya9jw6 & Fb9jw6);
assign Fb9jw6 = (Mb9jw6 & Tb9jw6);
assign Tb9jw6 = (Ac9jw6 & Hc9jw6);
assign Hc9jw6 = (Oc9jw6 & Vc9jw6);
assign Vc9jw6 = (~(vis_psp_o[9] & N32ov6));
assign Oc9jw6 = (~(U32ov6 & Pic7z6[9]));
assign Ac9jw6 = (Cd9jw6 & Jd9jw6);
assign Jd9jw6 = (~(vis_msp_o[9] & P42ov6));
assign Cd9jw6 = (~(vis_r12_o[9] & W42ov6));
assign Mb9jw6 = (Qd9jw6 & Xd9jw6);
assign Xd9jw6 = (Ee9jw6 & Le9jw6);
assign Le9jw6 = (~(vis_r11_o[9] & F62ov6));
assign Ee9jw6 = (~(vis_r10_o[9] & M62ov6));
assign Qd9jw6 = (Se9jw6 & Ze9jw6);
assign Ze9jw6 = (~(vis_r9_o[9] & H72ov6));
assign Se9jw6 = (~(vis_r8_o[9] & O72ov6));
assign Ya9jw6 = (Gf9jw6 & Nf9jw6);
assign Nf9jw6 = (Uf9jw6 & Bg9jw6);
assign Bg9jw6 = (Ig9jw6 & Pg9jw6);
assign Pg9jw6 = (~(vis_r7_o[9] & L92ov6));
assign Ig9jw6 = (~(vis_r6_o[9] & S92ov6));
assign Uf9jw6 = (Wg9jw6 & Dh9jw6);
assign Dh9jw6 = (~(vis_r5_o[9] & Na2ov6));
assign Wg9jw6 = (~(vis_r4_o[9] & Ua2ov6));
assign Gf9jw6 = (Kh9jw6 & Rh9jw6);
assign Rh9jw6 = (Yh9jw6 & Fi9jw6);
assign Fi9jw6 = (~(vis_r3_o[9] & Dc2ov6));
assign Yh9jw6 = (~(vis_r2_o[9] & Kc2ov6));
assign Kh9jw6 = (Mi9jw6 & Ti9jw6);
assign Ti9jw6 = (~(vis_r1_o[9] & Fd2ov6));
assign Mi9jw6 = (~(vis_r0_o[9] & Md2ov6));
assign Ka9jw6 = (~(Td2ov6 & Lbyiw6));
assign Lbyiw6 = (Spyiw6 ? O1a7z6 : Gli7z6[9]);
assign O1a7z6 = (~(Aj9jw6 & Hj9jw6));
assign Hj9jw6 = (~(Nqyiw6 & Jwznv6));
assign Aj9jw6 = (Oj9jw6 & Vj9jw6);
assign Vj9jw6 = (~(Pdc7z6[9] & Ouyiw6));
assign Oj9jw6 = (~(Vuyiw6 & Ck9jw6));
assign Ck9jw6 = (~(Jk9jw6 & Qk9jw6));
assign Qk9jw6 = (Xk9jw6 & El9jw6);
assign El9jw6 = (Ll9jw6 & Sl9jw6);
assign Sl9jw6 = (Zl9jw6 & Ns3jw6);
assign Zl9jw6 = (~(Gm9jw6 & Uxyiw6));
assign Gm9jw6 = (Kxb7z6[9] & Nm9jw6);
assign Ll9jw6 = (Um9jw6 & Bn9jw6);
assign Bn9jw6 = (~(In9jw6 & Pn9jw6));
assign In9jw6 = (~(Wn9jw6 & Quziw6));
assign Wn9jw6 = (Do9jw6 & Ko9jw6);
assign Ko9jw6 = (Nm9jw6 | Ninnv6);
assign Nm9jw6 = (Ro9jw6 | Rje7z6[9]);
assign Do9jw6 = (~(Ofnnv6 & Ro9jw6));
assign Um9jw6 = (~(Io3ov6 & C73ov6));
assign Io3ov6 = (~(Mp2jw6 ^ Dte7z6[1]));
assign Mp2jw6 = (T3cdt6 ? C6jnv6 : Hy3ov6);
assign Xk9jw6 = (Yo9jw6 & Fp9jw6);
assign Fp9jw6 = (Mp9jw6 & Tp9jw6);
assign Tp9jw6 = (~(Ak3ov6 & Ug3ov6));
assign Mp9jw6 = (~(J73ov6 & Ia3ov6));
assign Yo9jw6 = (Aq9jw6 & Hq9jw6);
assign Hq9jw6 = (~(T0ziw6 & Rje7z6[9]));
assign Aq9jw6 = (Ryfov6 | Oq9jw6);
assign Jk9jw6 = (Vq9jw6 & Cr9jw6);
assign Cr9jw6 = (Jr9jw6 & Qr9jw6);
assign Qr9jw6 = (Xr9jw6 & Es9jw6);
assign Es9jw6 = (~(L0g7z6[9] & J2ziw6));
assign Xr9jw6 = (~(L0g7z6[25] & Q2ziw6));
assign Jr9jw6 = (Ls9jw6 & Ss9jw6);
assign Ss9jw6 = (~(O1ziw6 & Onf7z6[9]));
assign Ls9jw6 = (~(U4ziw6 & Fhc7z6[9]));
assign Vq9jw6 = (Zs9jw6 & Nv2ov6);
assign Nv2ov6 = (Gt9jw6 & Nt9jw6);
assign Nt9jw6 = (~(Ut9jw6 & Ttmnv6));
assign Ut9jw6 = (~(Humnv6 | Icziw6));
assign Gt9jw6 = (~(Bu9jw6 & Ubziw6));
assign Bu9jw6 = (~(Ttmnv6 ^ Humnv6));
assign Humnv6 = (Iu9jw6 ^ Mennv6);
assign Iu9jw6 = (~(Pu9jw6 & Wu9jw6));
assign Wu9jw6 = (Dv9jw6 & Kv9jw6);
assign Kv9jw6 = (Rv9jw6 & Yv9jw6);
assign Yv9jw6 = (~(Yxf7z6[11] & Su0jw6));
assign Rv9jw6 = (Fw9jw6 & Mw9jw6);
assign Mw9jw6 = (~(Yxf7z6[9] & Nv0jw6));
assign Fw9jw6 = (~(Yxf7z6[10] & Uv0jw6));
assign Dv9jw6 = (Tw9jw6 & Ax9jw6);
assign Ax9jw6 = (~(Yxf7z6[12] & Pw0jw6));
assign Tw9jw6 = (Hx9jw6 | Dx0jw6);
assign Pu9jw6 = (Ox9jw6 & Vx9jw6);
assign Vx9jw6 = (Cy9jw6 & Jy9jw6);
assign Jy9jw6 = (~(Onf7z6[9] & My0jw6));
assign Cy9jw6 = (Qy9jw6 & Xy9jw6);
assign Xy9jw6 = (~(Hz0jw6 & Kxb7z6[9]));
assign Qy9jw6 = (~(Oz0jw6 & Fhc7z6[9]));
assign Ox9jw6 = (Ez9jw6 & Lz9jw6);
assign Lz9jw6 = (~(Onf7z6[25] & J01jw6));
assign Ez9jw6 = (~(Alf7z6[9] & Q01jw6));
assign Ttmnv6 = (~(Sz9jw6 ^ Tennv6));
assign Sz9jw6 = (~(Zz9jw6 & G0ajw6));
assign G0ajw6 = (~(Yxf7z6[9] & Gbziw6));
assign Zz9jw6 = (~(Kxb7z6[9] & Nbziw6));
assign Zs9jw6 = (N0ajw6 & U0ajw6);
assign U0ajw6 = (~(Z3ziw6 & Fhc7z6[22]));
assign N0ajw6 = (~(A4mdt6 & Oztiw6));
assign I99jw6 = (B1ajw6 & I1ajw6);
assign I1ajw6 = (~(Ve2ov6 & vis_pc_o[9]));
assign B1ajw6 = (~(Fhc7z6[9] & Cf2ov6));
assign U3z7v6 = (~(P1ajw6 & W1ajw6));
assign W1ajw6 = (D2ajw6 & K2ajw6);
assign K2ajw6 = (Eu9ov6 | R2ajw6);
assign D2ajw6 = (Y2ajw6 & F3ajw6);
assign F3ajw6 = (~(Gv9ov6 & O9yiw6));
assign Y2ajw6 = (~(Uv9ov6 & Sz97z6));
assign P1ajw6 = (M3ajw6 & T3ajw6);
assign T3ajw6 = (~(Pw9ov6 & Kxb7z6[17]));
assign M3ajw6 = (A4ajw6 & H4ajw6);
assign H4ajw6 = (~(Kx9ov6 & vis_pc_o[17]));
assign A4ajw6 = (~(Gli7z6[17] & Rx9ov6));
assign N3z7v6 = (~(O4ajw6 & V4ajw6));
assign V4ajw6 = (C5ajw6 & J5ajw6);
assign J5ajw6 = (~(H02ov6 & Sz97z6));
assign C5ajw6 = (Q5ajw6 & X5ajw6);
assign X5ajw6 = (C12ov6 | Maknv6);
assign Maknv6 = (E6ajw6 & L6ajw6);
assign L6ajw6 = (S6ajw6 & Z6ajw6);
assign Z6ajw6 = (G7ajw6 & N7ajw6);
assign N7ajw6 = (U7ajw6 & B8ajw6);
assign B8ajw6 = (~(vis_psp_o[17] & N32ov6));
assign U7ajw6 = (~(U32ov6 & Pic7z6[17]));
assign G7ajw6 = (I8ajw6 & P8ajw6);
assign P8ajw6 = (~(vis_msp_o[17] & P42ov6));
assign I8ajw6 = (~(vis_r12_o[17] & W42ov6));
assign S6ajw6 = (W8ajw6 & D9ajw6);
assign D9ajw6 = (K9ajw6 & R9ajw6);
assign R9ajw6 = (~(vis_r11_o[17] & F62ov6));
assign K9ajw6 = (~(vis_r10_o[17] & M62ov6));
assign W8ajw6 = (Y9ajw6 & Faajw6);
assign Faajw6 = (~(vis_r9_o[17] & H72ov6));
assign Y9ajw6 = (~(vis_r8_o[17] & O72ov6));
assign E6ajw6 = (Maajw6 & Taajw6);
assign Taajw6 = (Abajw6 & Hbajw6);
assign Hbajw6 = (Obajw6 & Vbajw6);
assign Vbajw6 = (~(vis_r7_o[17] & L92ov6));
assign Obajw6 = (~(vis_r6_o[17] & S92ov6));
assign Abajw6 = (Ccajw6 & Jcajw6);
assign Jcajw6 = (~(vis_r5_o[17] & Na2ov6));
assign Ccajw6 = (~(vis_r4_o[17] & Ua2ov6));
assign Maajw6 = (Qcajw6 & Xcajw6);
assign Xcajw6 = (Edajw6 & Ldajw6);
assign Ldajw6 = (~(vis_r3_o[17] & Dc2ov6));
assign Edajw6 = (~(vis_r2_o[17] & Kc2ov6));
assign Qcajw6 = (Sdajw6 & Zdajw6);
assign Zdajw6 = (~(vis_r1_o[17] & Fd2ov6));
assign Sdajw6 = (~(vis_r0_o[17] & Md2ov6));
assign Q5ajw6 = (~(Td2ov6 & O9yiw6));
assign O9yiw6 = (Spyiw6 ? Sz97z6 : Gli7z6[17]);
assign Sz97z6 = (~(Geajw6 & Neajw6));
assign Neajw6 = (~(Nqyiw6 & Zyynv6));
assign Geajw6 = (Ueajw6 & Bfajw6);
assign Bfajw6 = (~(Pdc7z6[17] & Ouyiw6));
assign Ueajw6 = (~(Vuyiw6 & Ifajw6));
assign Ifajw6 = (~(Pfajw6 & Wfajw6));
assign Wfajw6 = (Dgajw6 & Kgajw6);
assign Kgajw6 = (Rgajw6 & Ygajw6);
assign Ygajw6 = (Fhajw6 & Mhajw6);
assign Mhajw6 = (~(Thajw6 & Uxyiw6));
assign Thajw6 = (Kxb7z6[17] & Aiajw6);
assign Fhajw6 = (~(Hiajw6 & Oiajw6));
assign Hiajw6 = (~(Viajw6 & Quziw6));
assign Viajw6 = (Cjajw6 & Jjajw6);
assign Jjajw6 = (Aiajw6 | Ninnv6);
assign Aiajw6 = (Qjajw6 | Rje7z6[17]);
assign Cjajw6 = (~(Ofnnv6 & Qjajw6));
assign Rgajw6 = (Xjajw6 & Ekajw6);
assign Ekajw6 = (Zf3ov6 | U93ov6);
assign U93ov6 = (Ga7jw6 ^ Nu8jw6);
assign Ga7jw6 = (T3cdt6 ? V1c7z6[25] : A07jw6);
assign Xjajw6 = (~(J73ov6 & Ak3ov6));
assign Ak3ov6 = (~(Hx9jw6 ^ Dte7z6[1]));
assign Hx9jw6 = (T3cdt6 ? Qsohw6 : Oy3ov6);
assign Qsohw6 = (!V1c7z6[9]);
assign Dgajw6 = (Lkajw6 & Skajw6);
assign Skajw6 = (Zkajw6 & Glajw6);
assign Glajw6 = (~(F7ziw6 & Ia3ov6));
assign Ia3ov6 = (Nlajw6 ^ Dte7z6[1]);
assign Zkajw6 = (~(T0ziw6 & Rje7z6[17]));
assign Lkajw6 = (Ulajw6 & Bmajw6);
assign Bmajw6 = (Ryfov6 | Imajw6);
assign Ulajw6 = (~(L0g7z6[17] & J2ziw6));
assign Pfajw6 = (Pmajw6 & Wmajw6);
assign Wmajw6 = (Dnajw6 & Knajw6);
assign Knajw6 = (Rnajw6 & Ynajw6);
assign Ynajw6 = (~(Cqf7z6[1] & Q2ziw6));
assign Rnajw6 = (~(L0g7z6[1] & O1ziw6));
assign Dnajw6 = (Foajw6 & Moajw6);
assign Moajw6 = (~(U4ziw6 & V1c7z6[17]));
assign Foajw6 = (~(Z3ziw6 & Fhc7z6[14]));
assign Pmajw6 = (Toajw6 & Iw2ov6);
assign Iw2ov6 = (Apajw6 & Hpajw6);
assign Hpajw6 = (~(Opajw6 & D6nnv6));
assign Opajw6 = (~(K6nnv6 | Icziw6));
assign Apajw6 = (~(Vpajw6 & Ubziw6));
assign Vpajw6 = (~(D6nnv6 ^ K6nnv6));
assign K6nnv6 = (Cqajw6 ^ Mennv6);
assign Cqajw6 = (~(Jqajw6 & Qqajw6));
assign Qqajw6 = (Xqajw6 & Erajw6);
assign Erajw6 = (Lrajw6 & Srajw6);
assign Srajw6 = (~(Yxf7z6[19] & Su0jw6));
assign Lrajw6 = (Zrajw6 & Gsajw6);
assign Gsajw6 = (~(Yxf7z6[17] & Nv0jw6));
assign Zrajw6 = (~(Yxf7z6[18] & Uv0jw6));
assign Xqajw6 = (Nsajw6 & Usajw6);
assign Usajw6 = (~(Yxf7z6[20] & Pw0jw6));
assign Nsajw6 = (~(Nlajw6 & Rdziw6));
assign Nlajw6 = (T3cdt6 ? V1c7z6[17] : Oiajw6);
assign Jqajw6 = (Btajw6 & Itajw6);
assign Itajw6 = (Ptajw6 & Wtajw6);
assign Wtajw6 = (~(Onf7z6[17] & My0jw6));
assign Ptajw6 = (Duajw6 & Kuajw6);
assign Kuajw6 = (~(Hz0jw6 & Kxb7z6[17]));
assign Duajw6 = (~(Oz0jw6 & Fhc7z6[17]));
assign Btajw6 = (Ruajw6 & Yuajw6);
assign Yuajw6 = (~(Alf7z6[1] & J01jw6));
assign Ruajw6 = (~(Alf7z6[17] & Q01jw6));
assign D6nnv6 = (~(Fvajw6 ^ Tennv6));
assign Fvajw6 = (~(Mvajw6 & Tvajw6));
assign Tvajw6 = (~(Yxf7z6[1] & Laziw6));
assign Mvajw6 = (Awajw6 & Hwajw6);
assign Hwajw6 = (~(Yxf7z6[17] & Gbziw6));
assign Awajw6 = (~(Kxb7z6[17] & Nbziw6));
assign Toajw6 = (T7ziw6 & Owajw6);
assign Owajw6 = (~(Cnldt6 & Oztiw6));
assign O4ajw6 = (Vwajw6 & Cxajw6);
assign Cxajw6 = (~(Ve2ov6 & vis_pc_o[17]));
assign Vwajw6 = (~(Fhc7z6[17] & Cf2ov6));
assign G3z7v6 = (~(Jxajw6 & Qxajw6));
assign Qxajw6 = (Xxajw6 & Eyajw6);
assign Eyajw6 = (Eu9ov6 | Lyajw6);
assign Xxajw6 = (Syajw6 & Zyajw6);
assign Zyajw6 = (~(Gv9ov6 & Xayiw6));
assign Syajw6 = (~(Uv9ov6 & G1a7z6));
assign Jxajw6 = (Gzajw6 & Nzajw6);
assign Nzajw6 = (~(Pw9ov6 & Kxb7z6[11]));
assign Gzajw6 = (Uzajw6 & B0bjw6);
assign B0bjw6 = (~(Kx9ov6 & vis_pc_o[11]));
assign Uzajw6 = (~(Gli7z6[11] & Rx9ov6));
assign Z2z7v6 = (~(I0bjw6 & P0bjw6));
assign P0bjw6 = (W0bjw6 & D1bjw6);
assign D1bjw6 = (~(H02ov6 & G1a7z6));
assign W0bjw6 = (K1bjw6 & R1bjw6);
assign R1bjw6 = (~(Ktxiw6 & Lkknv6));
assign Lkknv6 = (~(Y1bjw6 & F2bjw6));
assign F2bjw6 = (M2bjw6 & T2bjw6);
assign T2bjw6 = (A3bjw6 & H3bjw6);
assign H3bjw6 = (O3bjw6 & V3bjw6);
assign V3bjw6 = (~(vis_psp_o[11] & N32ov6));
assign O3bjw6 = (~(U32ov6 & Pic7z6[11]));
assign A3bjw6 = (C4bjw6 & J4bjw6);
assign J4bjw6 = (~(vis_msp_o[11] & P42ov6));
assign C4bjw6 = (~(vis_r12_o[11] & W42ov6));
assign M2bjw6 = (Q4bjw6 & X4bjw6);
assign X4bjw6 = (E5bjw6 & L5bjw6);
assign L5bjw6 = (~(vis_r11_o[11] & F62ov6));
assign E5bjw6 = (~(vis_r10_o[11] & M62ov6));
assign Q4bjw6 = (S5bjw6 & Z5bjw6);
assign Z5bjw6 = (~(vis_r9_o[11] & H72ov6));
assign S5bjw6 = (~(vis_r8_o[11] & O72ov6));
assign Y1bjw6 = (G6bjw6 & N6bjw6);
assign N6bjw6 = (U6bjw6 & B7bjw6);
assign B7bjw6 = (I7bjw6 & P7bjw6);
assign P7bjw6 = (~(vis_r7_o[11] & L92ov6));
assign I7bjw6 = (~(vis_r6_o[11] & S92ov6));
assign U6bjw6 = (W7bjw6 & D8bjw6);
assign D8bjw6 = (~(vis_r5_o[11] & Na2ov6));
assign W7bjw6 = (~(vis_r4_o[11] & Ua2ov6));
assign G6bjw6 = (K8bjw6 & R8bjw6);
assign R8bjw6 = (Y8bjw6 & F9bjw6);
assign F9bjw6 = (~(vis_r3_o[11] & Dc2ov6));
assign Y8bjw6 = (~(vis_r2_o[11] & Kc2ov6));
assign K8bjw6 = (M9bjw6 & T9bjw6);
assign T9bjw6 = (~(vis_r1_o[11] & Fd2ov6));
assign M9bjw6 = (~(vis_r0_o[11] & Md2ov6));
assign K1bjw6 = (~(Td2ov6 & Xayiw6));
assign Xayiw6 = (Spyiw6 ? G1a7z6 : Gli7z6[11]);
assign G1a7z6 = (~(Aabjw6 & Habjw6));
assign Habjw6 = (~(Nqyiw6 & Hoznv6));
assign Aabjw6 = (Oabjw6 & Vabjw6);
assign Vabjw6 = (~(Pdc7z6[11] & Ouyiw6));
assign Oabjw6 = (~(Vuyiw6 & Cbbjw6));
assign Cbbjw6 = (~(Jbbjw6 & Qbbjw6));
assign Qbbjw6 = (Xbbjw6 & Ecbjw6);
assign Ecbjw6 = (Lcbjw6 & Scbjw6);
assign Scbjw6 = (Zcbjw6 & Ns3jw6);
assign Zcbjw6 = (~(Gdbjw6 & Uxyiw6));
assign Gdbjw6 = (Kxb7z6[11] & Ndbjw6);
assign Lcbjw6 = (Udbjw6 & Bebjw6);
assign Bebjw6 = (~(Iebjw6 & Pebjw6));
assign Iebjw6 = (~(Webjw6 & Quziw6));
assign Webjw6 = (Dfbjw6 & Kfbjw6);
assign Kfbjw6 = (Ndbjw6 | Ninnv6);
assign Ndbjw6 = (Rfbjw6 | Rje7z6[11]);
assign Dfbjw6 = (~(Ofnnv6 & Rfbjw6));
assign Udbjw6 = (~(Ri3ov6 & Ug3ov6));
assign Xbbjw6 = (Yfbjw6 & Fgbjw6);
assign Fgbjw6 = (Mgbjw6 & Tgbjw6);
assign Tgbjw6 = (~(Xl3ov6 & C73ov6));
assign Mgbjw6 = (~(J73ov6 & Hd3ov6));
assign Yfbjw6 = (Ahbjw6 & Hhbjw6);
assign Hhbjw6 = (~(T0ziw6 & Rje7z6[11]));
assign Ahbjw6 = (Ryfov6 | Ohbjw6);
assign Jbbjw6 = (Vhbjw6 & Cibjw6);
assign Cibjw6 = (Jibjw6 & Qibjw6);
assign Qibjw6 = (Xibjw6 & Ejbjw6);
assign Ejbjw6 = (~(L0g7z6[11] & J2ziw6));
assign Xibjw6 = (~(L0g7z6[27] & Q2ziw6));
assign Jibjw6 = (Ljbjw6 & Sjbjw6);
assign Sjbjw6 = (~(O1ziw6 & Onf7z6[11]));
assign Ljbjw6 = (~(U4ziw6 & Fhc7z6[11]));
assign Vhbjw6 = (Zjbjw6 & Bw2ov6);
assign Bw2ov6 = (Gkbjw6 & Nkbjw6);
assign Nkbjw6 = (~(Ukbjw6 & J9nnv6));
assign Ukbjw6 = (~(Q9nnv6 | Icziw6));
assign Gkbjw6 = (~(Blbjw6 & Ubziw6));
assign Blbjw6 = (~(J9nnv6 ^ Q9nnv6));
assign Q9nnv6 = (Ilbjw6 ^ Mennv6);
assign Ilbjw6 = (~(Plbjw6 & Wlbjw6));
assign Wlbjw6 = (Dmbjw6 & Kmbjw6);
assign Kmbjw6 = (Rmbjw6 & Ymbjw6);
assign Ymbjw6 = (~(Yxf7z6[13] & Su0jw6));
assign Rmbjw6 = (Fnbjw6 & Mnbjw6);
assign Mnbjw6 = (~(Yxf7z6[11] & Nv0jw6));
assign Fnbjw6 = (~(Yxf7z6[12] & Uv0jw6));
assign Dmbjw6 = (Tnbjw6 & Aobjw6);
assign Aobjw6 = (~(Yxf7z6[14] & Pw0jw6));
assign Tnbjw6 = (Hobjw6 | Dx0jw6);
assign Plbjw6 = (Oobjw6 & Vobjw6);
assign Vobjw6 = (Cpbjw6 & Jpbjw6);
assign Jpbjw6 = (~(Onf7z6[11] & My0jw6));
assign Cpbjw6 = (Qpbjw6 & Xpbjw6);
assign Xpbjw6 = (~(Hz0jw6 & Kxb7z6[11]));
assign Qpbjw6 = (~(Oz0jw6 & Fhc7z6[11]));
assign Oobjw6 = (Eqbjw6 & Lqbjw6);
assign Lqbjw6 = (~(Onf7z6[27] & J01jw6));
assign Eqbjw6 = (~(Alf7z6[11] & Q01jw6));
assign J9nnv6 = (~(Sqbjw6 ^ Tennv6));
assign Sqbjw6 = (~(Zqbjw6 & Grbjw6));
assign Grbjw6 = (~(Yxf7z6[11] & Gbziw6));
assign Zqbjw6 = (~(Kxb7z6[11] & Nbziw6));
assign Zjbjw6 = (Nrbjw6 & Urbjw6);
assign Urbjw6 = (~(Z3ziw6 & Fhc7z6[20]));
assign Nrbjw6 = (~(Uzldt6 & Oztiw6));
assign I0bjw6 = (Bsbjw6 & Isbjw6);
assign Isbjw6 = (~(Ve2ov6 & vis_pc_o[11]));
assign Bsbjw6 = (~(Fhc7z6[11] & Cf2ov6));
assign S2z7v6 = (~(Psbjw6 & Wsbjw6));
assign Wsbjw6 = (Dtbjw6 & Ktbjw6);
assign Ktbjw6 = (Eu9ov6 | Rtbjw6);
assign Dtbjw6 = (Ytbjw6 & Fubjw6);
assign Fubjw6 = (~(Gv9ov6 & H9yiw6));
assign Ytbjw6 = (~(Uv9ov6 & Kz97z6));
assign Psbjw6 = (Mubjw6 & Tubjw6);
assign Tubjw6 = (~(Pw9ov6 & Kxb7z6[19]));
assign Mubjw6 = (Avbjw6 & Hvbjw6);
assign Hvbjw6 = (~(Kx9ov6 & vis_pc_o[19]));
assign Avbjw6 = (~(Gli7z6[19] & Rx9ov6));
assign L2z7v6 = (~(Ovbjw6 & Vvbjw6));
assign Vvbjw6 = (Cwbjw6 & Jwbjw6);
assign Jwbjw6 = (~(H02ov6 & Kz97z6));
assign Cwbjw6 = (Qwbjw6 & Xwbjw6);
assign Xwbjw6 = (C12ov6 | G7knv6);
assign G7knv6 = (Exbjw6 & Lxbjw6);
assign Lxbjw6 = (Sxbjw6 & Zxbjw6);
assign Zxbjw6 = (Gybjw6 & Nybjw6);
assign Nybjw6 = (Uybjw6 & Bzbjw6);
assign Bzbjw6 = (~(vis_psp_o[19] & N32ov6));
assign Uybjw6 = (~(U32ov6 & Pic7z6[19]));
assign Gybjw6 = (Izbjw6 & Pzbjw6);
assign Pzbjw6 = (~(vis_msp_o[19] & P42ov6));
assign Izbjw6 = (~(vis_r12_o[19] & W42ov6));
assign Sxbjw6 = (Wzbjw6 & D0cjw6);
assign D0cjw6 = (K0cjw6 & R0cjw6);
assign R0cjw6 = (~(vis_r11_o[19] & F62ov6));
assign K0cjw6 = (~(vis_r10_o[19] & M62ov6));
assign Wzbjw6 = (Y0cjw6 & F1cjw6);
assign F1cjw6 = (~(vis_r9_o[19] & H72ov6));
assign Y0cjw6 = (~(vis_r8_o[19] & O72ov6));
assign Exbjw6 = (M1cjw6 & T1cjw6);
assign T1cjw6 = (A2cjw6 & H2cjw6);
assign H2cjw6 = (O2cjw6 & V2cjw6);
assign V2cjw6 = (~(vis_r7_o[19] & L92ov6));
assign O2cjw6 = (~(vis_r6_o[19] & S92ov6));
assign A2cjw6 = (C3cjw6 & J3cjw6);
assign J3cjw6 = (~(vis_r5_o[19] & Na2ov6));
assign C3cjw6 = (~(vis_r4_o[19] & Ua2ov6));
assign M1cjw6 = (Q3cjw6 & X3cjw6);
assign X3cjw6 = (E4cjw6 & L4cjw6);
assign L4cjw6 = (~(vis_r3_o[19] & Dc2ov6));
assign E4cjw6 = (~(vis_r2_o[19] & Kc2ov6));
assign Q3cjw6 = (S4cjw6 & Z4cjw6);
assign Z4cjw6 = (~(vis_r1_o[19] & Fd2ov6));
assign S4cjw6 = (~(vis_r0_o[19] & Md2ov6));
assign Qwbjw6 = (~(Td2ov6 & H9yiw6));
assign H9yiw6 = (Spyiw6 ? Kz97z6 : Gli7z6[19]);
assign Kz97z6 = (~(G5cjw6 & N5cjw6));
assign N5cjw6 = (~(Nqyiw6 & Vpynv6));
assign G5cjw6 = (U5cjw6 & B6cjw6);
assign B6cjw6 = (~(Pdc7z6[19] & Ouyiw6));
assign U5cjw6 = (~(Vuyiw6 & I6cjw6));
assign I6cjw6 = (~(P6cjw6 & W6cjw6));
assign W6cjw6 = (D7cjw6 & K7cjw6);
assign K7cjw6 = (R7cjw6 & Y7cjw6);
assign Y7cjw6 = (F8cjw6 & M8cjw6);
assign M8cjw6 = (~(T8cjw6 & Uxyiw6));
assign T8cjw6 = (Kxb7z6[19] & A9cjw6);
assign F8cjw6 = (~(H9cjw6 & O9cjw6));
assign H9cjw6 = (~(V9cjw6 & Quziw6));
assign V9cjw6 = (Cacjw6 & Jacjw6);
assign Jacjw6 = (A9cjw6 | Ninnv6);
assign A9cjw6 = (Qacjw6 | Rje7z6[19]);
assign Cacjw6 = (~(Ofnnv6 & Qacjw6));
assign R7cjw6 = (Xacjw6 & Ebcjw6);
assign Ebcjw6 = (~(J73ov6 & Ri3ov6));
assign Xacjw6 = (~(F7ziw6 & Hd3ov6));
assign D7cjw6 = (Lbcjw6 & Sbcjw6);
assign Sbcjw6 = (Zbcjw6 & Gccjw6);
assign Gccjw6 = (~(R6ziw6 & Ad3ov6));
assign Zbcjw6 = (~(T0ziw6 & Rje7z6[19]));
assign Lbcjw6 = (Nccjw6 & Uccjw6);
assign Uccjw6 = (Ryfov6 | Bdcjw6);
assign Nccjw6 = (~(L0g7z6[19] & J2ziw6));
assign P6cjw6 = (Idcjw6 & Pdcjw6);
assign Pdcjw6 = (Wdcjw6 & Decjw6);
assign Decjw6 = (Kecjw6 & Recjw6);
assign Recjw6 = (~(Cqf7z6[3] & Q2ziw6));
assign Kecjw6 = (~(L0g7z6[3] & O1ziw6));
assign Wdcjw6 = (Yecjw6 & Ffcjw6);
assign Ffcjw6 = (~(U4ziw6 & V1c7z6[19]));
assign Yecjw6 = (~(Z3ziw6 & Fhc7z6[12]));
assign Idcjw6 = (Mfcjw6 & My2ov6);
assign My2ov6 = (Tfcjw6 & Agcjw6);
assign Agcjw6 = (~(Hgcjw6 & B5nnv6));
assign Hgcjw6 = (~(I5nnv6 | Icziw6));
assign Tfcjw6 = (~(Ogcjw6 & Ubziw6));
assign Ogcjw6 = (~(B5nnv6 ^ I5nnv6));
assign I5nnv6 = (Vgcjw6 ^ Mennv6);
assign Vgcjw6 = (~(Chcjw6 & Jhcjw6));
assign Jhcjw6 = (Qhcjw6 & Xhcjw6);
assign Xhcjw6 = (Eicjw6 & Licjw6);
assign Licjw6 = (~(Yxf7z6[21] & Su0jw6));
assign Eicjw6 = (Sicjw6 & Zicjw6);
assign Zicjw6 = (~(Yxf7z6[19] & Nv0jw6));
assign Sicjw6 = (~(Yxf7z6[20] & Uv0jw6));
assign Qhcjw6 = (Gjcjw6 & Njcjw6);
assign Njcjw6 = (~(Yxf7z6[22] & Pw0jw6));
assign Gjcjw6 = (~(Ujcjw6 & Rdziw6));
assign Chcjw6 = (Bkcjw6 & Ikcjw6);
assign Ikcjw6 = (Pkcjw6 & Wkcjw6);
assign Wkcjw6 = (~(Onf7z6[19] & My0jw6));
assign Pkcjw6 = (Dlcjw6 & Klcjw6);
assign Klcjw6 = (~(Hz0jw6 & Kxb7z6[19]));
assign Dlcjw6 = (~(Oz0jw6 & Fhc7z6[19]));
assign Bkcjw6 = (Rlcjw6 & Ylcjw6);
assign Ylcjw6 = (~(Alf7z6[3] & J01jw6));
assign Rlcjw6 = (~(Alf7z6[19] & Q01jw6));
assign B5nnv6 = (~(Fmcjw6 ^ Tennv6));
assign Fmcjw6 = (~(Mmcjw6 & Tmcjw6));
assign Tmcjw6 = (~(Yxf7z6[3] & Laziw6));
assign Mmcjw6 = (Ikg6x6 & Pkg6x6);
assign Pkg6x6 = (~(Yxf7z6[19] & Gbziw6));
assign Ikg6x6 = (~(Kxb7z6[19] & Nbziw6));
assign Mfcjw6 = (T7ziw6 & Wkg6x6);
assign Wkg6x6 = (~(Wildt6 & Oztiw6));
assign Ovbjw6 = (Dlg6x6 & Klg6x6);
assign Klg6x6 = (~(Ve2ov6 & vis_pc_o[19]));
assign Dlg6x6 = (~(Fhc7z6[19] & Cf2ov6));
assign E2z7v6 = (~(Rlg6x6 & Ylg6x6));
assign Ylg6x6 = (Fmg6x6 & Mmg6x6);
assign Mmg6x6 = (Eu9ov6 | Tmg6x6);
assign Fmg6x6 = (Ang6x6 & Hng6x6);
assign Hng6x6 = (~(Gv9ov6 & Qayiw6));
assign Ang6x6 = (~(Uv9ov6 & Y0a7z6));
assign Rlg6x6 = (Ong6x6 & Vng6x6);
assign Vng6x6 = (~(Pw9ov6 & Kxb7z6[12]));
assign Ong6x6 = (Cog6x6 & Jog6x6);
assign Jog6x6 = (~(Kx9ov6 & vis_pc_o[12]));
assign Cog6x6 = (~(Gli7z6[12] & Rx9ov6));
assign X1z7v6 = (~(Qog6x6 & Xog6x6));
assign Xog6x6 = (Epg6x6 & Lpg6x6);
assign Lpg6x6 = (~(H02ov6 & Y0a7z6));
assign Epg6x6 = (Spg6x6 & Zpg6x6);
assign Zpg6x6 = (C12ov6 | Oiknv6);
assign Oiknv6 = (Gqg6x6 & Nqg6x6);
assign Nqg6x6 = (Uqg6x6 & Brg6x6);
assign Brg6x6 = (Irg6x6 & Prg6x6);
assign Prg6x6 = (Wrg6x6 & Dsg6x6);
assign Dsg6x6 = (~(vis_psp_o[12] & N32ov6));
assign Wrg6x6 = (~(U32ov6 & Pic7z6[12]));
assign Irg6x6 = (Ksg6x6 & Rsg6x6);
assign Rsg6x6 = (~(vis_msp_o[12] & P42ov6));
assign Ksg6x6 = (~(vis_r12_o[12] & W42ov6));
assign Uqg6x6 = (Ysg6x6 & Ftg6x6);
assign Ftg6x6 = (Mtg6x6 & Ttg6x6);
assign Ttg6x6 = (~(vis_r11_o[12] & F62ov6));
assign Mtg6x6 = (~(vis_r10_o[12] & M62ov6));
assign Ysg6x6 = (Aug6x6 & Hug6x6);
assign Hug6x6 = (~(vis_r9_o[12] & H72ov6));
assign Aug6x6 = (~(vis_r8_o[12] & O72ov6));
assign Gqg6x6 = (Oug6x6 & Vug6x6);
assign Vug6x6 = (Cvg6x6 & Jvg6x6);
assign Jvg6x6 = (Qvg6x6 & Xvg6x6);
assign Xvg6x6 = (~(vis_r7_o[12] & L92ov6));
assign Qvg6x6 = (~(vis_r6_o[12] & S92ov6));
assign Cvg6x6 = (Ewg6x6 & Lwg6x6);
assign Lwg6x6 = (~(vis_r5_o[12] & Na2ov6));
assign Ewg6x6 = (~(vis_r4_o[12] & Ua2ov6));
assign Oug6x6 = (Swg6x6 & Zwg6x6);
assign Zwg6x6 = (Gxg6x6 & Nxg6x6);
assign Nxg6x6 = (~(vis_r3_o[12] & Dc2ov6));
assign Gxg6x6 = (~(vis_r2_o[12] & Kc2ov6));
assign Swg6x6 = (Uxg6x6 & Byg6x6);
assign Byg6x6 = (~(vis_r1_o[12] & Fd2ov6));
assign Uxg6x6 = (~(vis_r0_o[12] & Md2ov6));
assign Spg6x6 = (~(Td2ov6 & Qayiw6));
assign Qayiw6 = (Spyiw6 ? Y0a7z6 : Gli7z6[12]);
assign Y0a7z6 = (~(Iyg6x6 & Pyg6x6));
assign Pyg6x6 = (~(Nqyiw6 & Gkznv6));
assign Iyg6x6 = (Wyg6x6 & Dzg6x6);
assign Dzg6x6 = (~(Pdc7z6[12] & Ouyiw6));
assign Wyg6x6 = (~(Vuyiw6 & Kzg6x6));
assign Kzg6x6 = (~(Rzg6x6 & Yzg6x6));
assign Yzg6x6 = (F0h6x6 & M0h6x6);
assign M0h6x6 = (T0h6x6 & A1h6x6);
assign A1h6x6 = (H1h6x6 & Ns3jw6);
assign H1h6x6 = (~(O1h6x6 & Uxyiw6));
assign O1h6x6 = (Kxb7z6[12] & V1h6x6);
assign T0h6x6 = (C2h6x6 & J2h6x6);
assign J2h6x6 = (~(Q2h6x6 & X2h6x6));
assign Q2h6x6 = (~(E3h6x6 & Quziw6));
assign E3h6x6 = (L3h6x6 & S3h6x6);
assign S3h6x6 = (V1h6x6 | Ninnv6);
assign V1h6x6 = (~(Z3h6x6 & G4h6x6));
assign Z3h6x6 = (!Rje7z6[12]);
assign L3h6x6 = (G4h6x6 | Evziw6);
assign C2h6x6 = (~(Em3ov6 & C73ov6));
assign F0h6x6 = (N4h6x6 & U4h6x6);
assign U4h6x6 = (B5h6x6 & I5h6x6);
assign I5h6x6 = (~(Ki3ov6 & Ug3ov6));
assign B5h6x6 = (~(J73ov6 & Od3ov6));
assign N4h6x6 = (P5h6x6 & W5h6x6);
assign W5h6x6 = (~(T0ziw6 & Rje7z6[12]));
assign P5h6x6 = (G4h6x6 | Ryfov6);
assign Rzg6x6 = (D6h6x6 & K6h6x6);
assign K6h6x6 = (R6h6x6 & Y6h6x6);
assign Y6h6x6 = (F7h6x6 & M7h6x6);
assign M7h6x6 = (~(L0g7z6[12] & J2ziw6));
assign F7h6x6 = (~(L0g7z6[28] & Q2ziw6));
assign R6h6x6 = (T7h6x6 & A8h6x6);
assign A8h6x6 = (~(O1ziw6 & Onf7z6[12]));
assign T7h6x6 = (~(U4ziw6 & Fhc7z6[12]));
assign D6h6x6 = (H8h6x6 & Fy2ov6);
assign Fy2ov6 = (O8h6x6 & V8h6x6);
assign V8h6x6 = (~(C9h6x6 & V8nnv6));
assign C9h6x6 = (~(C9nnv6 | Icziw6));
assign O8h6x6 = (~(J9h6x6 & Ubziw6));
assign J9h6x6 = (~(V8nnv6 ^ C9nnv6));
assign C9nnv6 = (Q9h6x6 ^ Mennv6);
assign Q9h6x6 = (~(X9h6x6 & Eah6x6));
assign Eah6x6 = (Lah6x6 & Sah6x6);
assign Sah6x6 = (Zah6x6 & Gbh6x6);
assign Gbh6x6 = (~(Yxf7z6[14] & Su0jw6));
assign Zah6x6 = (Nbh6x6 & Ubh6x6);
assign Ubh6x6 = (~(Yxf7z6[12] & Nv0jw6));
assign Nbh6x6 = (~(Yxf7z6[13] & Uv0jw6));
assign Lah6x6 = (Bch6x6 & Ich6x6);
assign Ich6x6 = (~(Pw0jw6 & Yxf7z6[15]));
assign Bch6x6 = (Pch6x6 | Dx0jw6);
assign X9h6x6 = (Wch6x6 & Ddh6x6);
assign Ddh6x6 = (Kdh6x6 & Rdh6x6);
assign Rdh6x6 = (~(Onf7z6[12] & My0jw6));
assign Kdh6x6 = (Ydh6x6 & Feh6x6);
assign Feh6x6 = (~(Hz0jw6 & Kxb7z6[12]));
assign Ydh6x6 = (~(Oz0jw6 & Fhc7z6[12]));
assign Wch6x6 = (Meh6x6 & Teh6x6);
assign Teh6x6 = (~(J01jw6 & Onf7z6[28]));
assign Meh6x6 = (~(Q01jw6 & Alf7z6[12]));
assign V8nnv6 = (~(Afh6x6 ^ Tennv6));
assign Afh6x6 = (~(Hfh6x6 & Ofh6x6));
assign Ofh6x6 = (~(Yxf7z6[12] & Gbziw6));
assign Hfh6x6 = (~(Kxb7z6[12] & Nbziw6));
assign H8h6x6 = (Vfh6x6 & Cgh6x6);
assign Cgh6x6 = (~(Z3ziw6 & Fhc7z6[19]));
assign Vfh6x6 = (~(Rxldt6 & Oztiw6));
assign Qog6x6 = (Jgh6x6 & Qgh6x6);
assign Qgh6x6 = (~(Ve2ov6 & vis_pc_o[12]));
assign Jgh6x6 = (~(Fhc7z6[12] & Cf2ov6));
assign Q1z7v6 = (~(Xgh6x6 & Ehh6x6));
assign Ehh6x6 = (Lhh6x6 & Shh6x6);
assign Shh6x6 = (Eu9ov6 | Zhh6x6);
assign Lhh6x6 = (Gih6x6 & Nih6x6);
assign Nih6x6 = (~(Gv9ov6 & Ncyiw6));
assign Gih6x6 = (~(Uv9ov6 & U2a7z6));
assign Xgh6x6 = (Uih6x6 & Bjh6x6);
assign Bjh6x6 = (~(Pw9ov6 & Kxb7z6[3]));
assign Uih6x6 = (Ijh6x6 & Pjh6x6);
assign Pjh6x6 = (~(Kx9ov6 & vis_pc_o[3]));
assign Ijh6x6 = (~(Gli7z6[3] & Rx9ov6));
assign J1z7v6 = (~(Wjh6x6 & Dkh6x6));
assign Dkh6x6 = (Kkh6x6 & Rkh6x6);
assign Rkh6x6 = (~(H02ov6 & U2a7z6));
assign Kkh6x6 = (Ykh6x6 & Flh6x6);
assign Flh6x6 = (C12ov6 | Mijnv6);
assign Mijnv6 = (Mlh6x6 & Tlh6x6);
assign Tlh6x6 = (Amh6x6 & Hmh6x6);
assign Hmh6x6 = (Omh6x6 & Vmh6x6);
assign Vmh6x6 = (Cnh6x6 & Jnh6x6);
assign Jnh6x6 = (~(vis_psp_o[3] & N32ov6));
assign Cnh6x6 = (~(U32ov6 & Pic7z6[3]));
assign Omh6x6 = (Qnh6x6 & Xnh6x6);
assign Xnh6x6 = (~(vis_msp_o[3] & P42ov6));
assign Qnh6x6 = (~(vis_r12_o[3] & W42ov6));
assign Amh6x6 = (Eoh6x6 & Loh6x6);
assign Loh6x6 = (Soh6x6 & Zoh6x6);
assign Zoh6x6 = (~(vis_r11_o[3] & F62ov6));
assign Soh6x6 = (~(vis_r10_o[3] & M62ov6));
assign Eoh6x6 = (Gph6x6 & Nph6x6);
assign Nph6x6 = (~(vis_r9_o[3] & H72ov6));
assign Gph6x6 = (~(vis_r8_o[3] & O72ov6));
assign Mlh6x6 = (Uph6x6 & Bqh6x6);
assign Bqh6x6 = (Iqh6x6 & Pqh6x6);
assign Pqh6x6 = (Wqh6x6 & Drh6x6);
assign Drh6x6 = (~(vis_r7_o[3] & L92ov6));
assign Wqh6x6 = (~(vis_r6_o[3] & S92ov6));
assign Iqh6x6 = (Krh6x6 & Rrh6x6);
assign Rrh6x6 = (~(vis_r5_o[3] & Na2ov6));
assign Krh6x6 = (~(vis_r4_o[3] & Ua2ov6));
assign Uph6x6 = (Yrh6x6 & Fsh6x6);
assign Fsh6x6 = (Msh6x6 & Tsh6x6);
assign Tsh6x6 = (~(vis_r3_o[3] & Dc2ov6));
assign Msh6x6 = (~(vis_r2_o[3] & Kc2ov6));
assign Yrh6x6 = (Ath6x6 & Hth6x6);
assign Hth6x6 = (~(vis_r1_o[3] & Fd2ov6));
assign Ath6x6 = (~(vis_r0_o[3] & Md2ov6));
assign Ykh6x6 = (~(Td2ov6 & Ncyiw6));
assign Ncyiw6 = (Spyiw6 ? U2a7z6 : Gli7z6[3]);
assign U2a7z6 = (~(Oth6x6 & Vth6x6));
assign Vth6x6 = (~(Nqyiw6 & Pk0ov6));
assign Oth6x6 = (Cuh6x6 & Juh6x6);
assign Juh6x6 = (~(Pdc7z6[3] & Ouyiw6));
assign Cuh6x6 = (~(Vuyiw6 & Quh6x6));
assign Quh6x6 = (~(Xuh6x6 & Evh6x6));
assign Evh6x6 = (Lvh6x6 & Svh6x6);
assign Svh6x6 = (Zvh6x6 & Gwh6x6);
assign Gwh6x6 = (Nwh6x6 & Uwh6x6);
assign Uwh6x6 = (~(Bxh6x6 & Uxyiw6));
assign Bxh6x6 = (Kxb7z6[3] & Ixh6x6);
assign Nwh6x6 = (~(Pxh6x6 & Jm0jw6));
assign Pxh6x6 = (Nob7z6[3] & Rslov6);
assign Zvh6x6 = (Wxh6x6 & Dyh6x6);
assign Dyh6x6 = (~(Kyh6x6 & Ryh6x6));
assign Kyh6x6 = (~(Yyh6x6 & Quziw6));
assign Yyh6x6 = (Fzh6x6 & Mzh6x6);
assign Mzh6x6 = (Ixh6x6 | Ninnv6);
assign Ixh6x6 = (Tzh6x6 | Rje7z6[3]);
assign Fzh6x6 = (~(Ofnnv6 & Tzh6x6));
assign Wxh6x6 = (~(Svziw6 & Wjnnv6));
assign Lvh6x6 = (A0i6x6 & H0i6x6);
assign H0i6x6 = (O0i6x6 & V0i6x6);
assign V0i6x6 = (~(Ri3ov6 & C73ov6));
assign Ri3ov6 = (~(Hobjw6 ^ Dte7z6[1]));
assign Hobjw6 = (T3cdt6 ? Ceohw6 : S04ov6);
assign O0i6x6 = (~(Ol0jw6 & Xl3ov6));
assign A0i6x6 = (C1i6x6 & J1i6x6);
assign J1i6x6 = (~(J73ov6 & Ad3ov6));
assign C1i6x6 = (~(T0ziw6 & Rje7z6[3]));
assign Xuh6x6 = (Q1i6x6 & X1i6x6);
assign X1i6x6 = (E2i6x6 & L2i6x6);
assign L2i6x6 = (S2i6x6 & Z2i6x6);
assign Z2i6x6 = (Ryfov6 | G3i6x6);
assign S2i6x6 = (~(L0g7z6[3] & J2ziw6));
assign E2i6x6 = (N3i6x6 & U3i6x6);
assign U3i6x6 = (~(L0g7z6[19] & Q2ziw6));
assign N3i6x6 = (~(O1ziw6 & Onf7z6[3]));
assign Q1i6x6 = (B4i6x6 & I4i6x6);
assign I4i6x6 = (P4i6x6 & W4i6x6);
assign W4i6x6 = (~(U4ziw6 & E3c7z6[3]));
assign P4i6x6 = (~(Z3ziw6 & Fhc7z6[28]));
assign B4i6x6 = (Az2ov6 & D5i6x6);
assign D5i6x6 = (~(Sgmdt6 & Oztiw6));
assign Az2ov6 = (K5i6x6 & R5i6x6);
assign R5i6x6 = (~(Y5i6x6 & Nxmnv6));
assign Y5i6x6 = (~(Uxmnv6 | Icziw6));
assign K5i6x6 = (~(F6i6x6 & Ubziw6));
assign F6i6x6 = (~(Nxmnv6 ^ Uxmnv6));
assign Uxmnv6 = (M6i6x6 ^ Mennv6);
assign M6i6x6 = (~(T6i6x6 & A7i6x6));
assign A7i6x6 = (H7i6x6 & O7i6x6);
assign O7i6x6 = (V7i6x6 & C8i6x6);
assign C8i6x6 = (~(Yxf7z6[5] & Su0jw6));
assign V7i6x6 = (J8i6x6 & Q8i6x6);
assign Q8i6x6 = (~(Yxf7z6[3] & Nv0jw6));
assign J8i6x6 = (~(Yxf7z6[4] & Uv0jw6));
assign H7i6x6 = (X8i6x6 & E9i6x6);
assign E9i6x6 = (~(Yxf7z6[6] & Pw0jw6));
assign X8i6x6 = (L9i6x6 | Dx0jw6);
assign T6i6x6 = (S9i6x6 & Z9i6x6);
assign Z9i6x6 = (Gai6x6 & Nai6x6);
assign Nai6x6 = (~(Onf7z6[3] & My0jw6));
assign Gai6x6 = (Uai6x6 & Bbi6x6);
assign Bbi6x6 = (~(Hz0jw6 & Kxb7z6[3]));
assign Uai6x6 = (~(Oz0jw6 & E3c7z6[3]));
assign S9i6x6 = (Ibi6x6 & Pbi6x6);
assign Pbi6x6 = (~(Onf7z6[19] & J01jw6));
assign Ibi6x6 = (~(Alf7z6[3] & Q01jw6));
assign Nxmnv6 = (~(Wbi6x6 ^ Tennv6));
assign Wbi6x6 = (~(Dci6x6 & Kci6x6));
assign Kci6x6 = (~(Yxf7z6[3] & Gbziw6));
assign Dci6x6 = (~(Kxb7z6[3] & Nbziw6));
assign Wjh6x6 = (Rci6x6 & Yci6x6);
assign Yci6x6 = (~(Ve2ov6 & vis_pc_o[3]));
assign Rci6x6 = (~(E3c7z6[3] & Cf2ov6));
assign C1z7v6 = (~(Fdi6x6 & Mdi6x6));
assign Mdi6x6 = (Tdi6x6 & Aei6x6);
assign Aei6x6 = (Eu9ov6 | Hei6x6);
assign Tdi6x6 = (Oei6x6 & Vei6x6);
assign Vei6x6 = (~(Gv9ov6 & Gcyiw6));
assign Oei6x6 = (~(Uv9ov6 & M2a7z6));
assign Fdi6x6 = (Cfi6x6 & Jfi6x6);
assign Jfi6x6 = (~(Pw9ov6 & Kxb7z6[5]));
assign Cfi6x6 = (Qfi6x6 & Xfi6x6);
assign Xfi6x6 = (~(Kx9ov6 & vis_pc_o[5]));
assign Qfi6x6 = (~(Gli7z6[5] & Rx9ov6));
assign V0z7v6 = (~(Egi6x6 & Lgi6x6));
assign Lgi6x6 = (Sgi6x6 & Zgi6x6);
assign Zgi6x6 = (~(H02ov6 & M2a7z6));
assign Sgi6x6 = (Ghi6x6 & Nhi6x6);
assign Nhi6x6 = (C12ov6 | Gfjnv6);
assign Gfjnv6 = (Uhi6x6 & Bii6x6);
assign Bii6x6 = (Iii6x6 & Pii6x6);
assign Pii6x6 = (Wii6x6 & Dji6x6);
assign Dji6x6 = (Kji6x6 & Rji6x6);
assign Rji6x6 = (~(vis_psp_o[5] & N32ov6));
assign Kji6x6 = (~(U32ov6 & Pic7z6[5]));
assign Wii6x6 = (Yji6x6 & Fki6x6);
assign Fki6x6 = (~(vis_msp_o[5] & P42ov6));
assign Yji6x6 = (~(vis_r12_o[5] & W42ov6));
assign Iii6x6 = (Mki6x6 & Tki6x6);
assign Tki6x6 = (Ali6x6 & Hli6x6);
assign Hli6x6 = (~(vis_r11_o[5] & F62ov6));
assign Ali6x6 = (~(vis_r10_o[5] & M62ov6));
assign Mki6x6 = (Oli6x6 & Vli6x6);
assign Vli6x6 = (~(vis_r9_o[5] & H72ov6));
assign Oli6x6 = (~(vis_r8_o[5] & O72ov6));
assign Uhi6x6 = (Cmi6x6 & Jmi6x6);
assign Jmi6x6 = (Qmi6x6 & Xmi6x6);
assign Xmi6x6 = (Eni6x6 & Lni6x6);
assign Lni6x6 = (~(vis_r7_o[5] & L92ov6));
assign Eni6x6 = (~(vis_r6_o[5] & S92ov6));
assign Qmi6x6 = (Sni6x6 & Zni6x6);
assign Zni6x6 = (~(vis_r5_o[5] & Na2ov6));
assign Sni6x6 = (~(vis_r4_o[5] & Ua2ov6));
assign Cmi6x6 = (Goi6x6 & Noi6x6);
assign Noi6x6 = (Uoi6x6 & Bpi6x6);
assign Bpi6x6 = (~(vis_r3_o[5] & Dc2ov6));
assign Uoi6x6 = (~(vis_r2_o[5] & Kc2ov6));
assign Goi6x6 = (Ipi6x6 & Ppi6x6);
assign Ppi6x6 = (~(vis_r1_o[5] & Fd2ov6));
assign Ipi6x6 = (~(vis_r0_o[5] & Md2ov6));
assign Ghi6x6 = (~(Td2ov6 & Gcyiw6));
assign Gcyiw6 = (Spyiw6 ? M2a7z6 : Gli7z6[5]);
assign M2a7z6 = (~(Wpi6x6 & Dqi6x6));
assign Dqi6x6 = (~(Nqyiw6 & Nc0ov6));
assign Wpi6x6 = (Kqi6x6 & Rqi6x6);
assign Rqi6x6 = (~(Pdc7z6[5] & Ouyiw6));
assign Kqi6x6 = (~(Vuyiw6 & Yqi6x6));
assign Yqi6x6 = (~(Fri6x6 & Mri6x6));
assign Mri6x6 = (Tri6x6 & Asi6x6);
assign Asi6x6 = (Hsi6x6 & Osi6x6);
assign Osi6x6 = (Vsi6x6 & Cti6x6);
assign Cti6x6 = (~(Jm0jw6 & Jti6x6));
assign Vsi6x6 = (Qti6x6 & Xti6x6);
assign Xti6x6 = (~(Eui6x6 & Uxyiw6));
assign Eui6x6 = (Kxb7z6[5] & Lui6x6);
assign Qti6x6 = (~(Xs3ov6 & Sui6x6));
assign Sui6x6 = (~(Zui6x6 & Quziw6));
assign Zui6x6 = (Gvi6x6 & Nvi6x6);
assign Nvi6x6 = (Lui6x6 | Ninnv6);
assign Lui6x6 = (Uvi6x6 | Rje7z6[5]);
assign Gvi6x6 = (~(Ofnnv6 & Uvi6x6));
assign Hsi6x6 = (Bwi6x6 & Iwi6x6);
assign Iwi6x6 = (~(Svziw6 & Bjnnv6));
assign Bjnnv6 = (Pwi6x6 & Wwi6x6);
assign Pwi6x6 = (~(Dxi6x6 | Kxi6x6));
assign Bwi6x6 = (~(J73ov6 & Rb3ov6));
assign Tri6x6 = (Rxi6x6 & Yxi6x6);
assign Yxi6x6 = (Fyi6x6 & Myi6x6);
assign Myi6x6 = (~(Yi3ov6 & C73ov6));
assign Fyi6x6 = (~(Ol0jw6 & Nn3ov6));
assign Rxi6x6 = (Tyi6x6 & Azi6x6);
assign Azi6x6 = (~(Hzi6x6 & Ppb7z6[5]));
assign Tyi6x6 = (~(T0ziw6 & Rje7z6[5]));
assign Fri6x6 = (Ozi6x6 & Vzi6x6);
assign Vzi6x6 = (C0j6x6 & J0j6x6);
assign J0j6x6 = (Q0j6x6 & X0j6x6);
assign X0j6x6 = (Ryfov6 | E1j6x6);
assign E1j6x6 = (!Uvi6x6);
assign Q0j6x6 = (~(L0g7z6[5] & J2ziw6));
assign C0j6x6 = (L1j6x6 & S1j6x6);
assign S1j6x6 = (~(L0g7z6[21] & Q2ziw6));
assign L1j6x6 = (~(O1ziw6 & Onf7z6[5]));
assign Ozi6x6 = (Z1j6x6 & G2j6x6);
assign G2j6x6 = (N2j6x6 & U2j6x6);
assign U2j6x6 = (~(U4ziw6 & Fhc7z6[5]));
assign N2j6x6 = (~(Z3ziw6 & Fhc7z6[26]));
assign Z1j6x6 = (Ty2ov6 & B3j6x6);
assign B3j6x6 = (~(Mcmdt6 & Oztiw6));
assign Ty2ov6 = (I3j6x6 & P3j6x6);
assign P3j6x6 = (~(W3j6x6 & Lwmnv6));
assign W3j6x6 = (~(Swmnv6 | Icziw6));
assign I3j6x6 = (~(D4j6x6 & Ubziw6));
assign D4j6x6 = (~(Lwmnv6 ^ Swmnv6));
assign Swmnv6 = (K4j6x6 ^ Mennv6);
assign K4j6x6 = (~(R4j6x6 & Y4j6x6));
assign Y4j6x6 = (F5j6x6 & M5j6x6);
assign M5j6x6 = (T5j6x6 & A6j6x6);
assign A6j6x6 = (~(Yxf7z6[7] & Su0jw6));
assign T5j6x6 = (H6j6x6 & O6j6x6);
assign O6j6x6 = (~(Yxf7z6[5] & Nv0jw6));
assign H6j6x6 = (~(Yxf7z6[6] & Uv0jw6));
assign F5j6x6 = (V6j6x6 & C7j6x6);
assign C7j6x6 = (~(Yxf7z6[8] & Pw0jw6));
assign V6j6x6 = (~(J7j6x6 & Rdziw6));
assign R4j6x6 = (Q7j6x6 & X7j6x6);
assign X7j6x6 = (E8j6x6 & L8j6x6);
assign L8j6x6 = (~(Onf7z6[5] & My0jw6));
assign E8j6x6 = (S8j6x6 & Z8j6x6);
assign Z8j6x6 = (~(Hz0jw6 & Kxb7z6[5]));
assign S8j6x6 = (~(Oz0jw6 & Fhc7z6[5]));
assign Q7j6x6 = (G9j6x6 & N9j6x6);
assign N9j6x6 = (~(Onf7z6[21] & J01jw6));
assign G9j6x6 = (~(Alf7z6[5] & Q01jw6));
assign Lwmnv6 = (~(U9j6x6 ^ Tennv6));
assign U9j6x6 = (~(Baj6x6 & Iaj6x6));
assign Iaj6x6 = (~(Yxf7z6[5] & Gbziw6));
assign Baj6x6 = (~(Kxb7z6[5] & Nbziw6));
assign Egi6x6 = (Paj6x6 & Waj6x6);
assign Waj6x6 = (~(Ve2ov6 & vis_pc_o[5]));
assign Paj6x6 = (~(Fhc7z6[5] & Cf2ov6));
assign O0z7v6 = (~(Dbj6x6 & Kbj6x6));
assign Kbj6x6 = (Rbj6x6 & Ybj6x6);
assign Ybj6x6 = (Eu9ov6 | Fcj6x6);
assign Rbj6x6 = (Mcj6x6 & Tcj6x6);
assign Tcj6x6 = (~(Gv9ov6 & T8yiw6));
assign Mcj6x6 = (~(Uv9ov6 & Uy97z6));
assign Dbj6x6 = (Adj6x6 & Hdj6x6);
assign Hdj6x6 = (~(Pw9ov6 & Kxb7z6[21]));
assign Adj6x6 = (Odj6x6 & Vdj6x6);
assign Vdj6x6 = (~(Kx9ov6 & vis_pc_o[21]));
assign Odj6x6 = (~(Gli7z6[21] & Rx9ov6));
assign H0z7v6 = (~(Cej6x6 & Jej6x6));
assign Jej6x6 = (Qej6x6 & Xej6x6);
assign Xej6x6 = (~(H02ov6 & Uy97z6));
assign Qej6x6 = (Efj6x6 & Lfj6x6);
assign Lfj6x6 = (C12ov6 | W1knv6);
assign W1knv6 = (Sfj6x6 & Zfj6x6);
assign Zfj6x6 = (Ggj6x6 & Ngj6x6);
assign Ngj6x6 = (Ugj6x6 & Bhj6x6);
assign Bhj6x6 = (Ihj6x6 & Phj6x6);
assign Phj6x6 = (~(vis_psp_o[21] & N32ov6));
assign Ihj6x6 = (~(U32ov6 & Pic7z6[21]));
assign Ugj6x6 = (Whj6x6 & Dij6x6);
assign Dij6x6 = (~(vis_msp_o[21] & P42ov6));
assign Whj6x6 = (~(vis_r12_o[21] & W42ov6));
assign Ggj6x6 = (Kij6x6 & Rij6x6);
assign Rij6x6 = (Yij6x6 & Fjj6x6);
assign Fjj6x6 = (~(vis_r11_o[21] & F62ov6));
assign Yij6x6 = (~(vis_r10_o[21] & M62ov6));
assign Kij6x6 = (Mjj6x6 & Tjj6x6);
assign Tjj6x6 = (~(vis_r9_o[21] & H72ov6));
assign Mjj6x6 = (~(vis_r8_o[21] & O72ov6));
assign Sfj6x6 = (Akj6x6 & Hkj6x6);
assign Hkj6x6 = (Okj6x6 & Vkj6x6);
assign Vkj6x6 = (Clj6x6 & Jlj6x6);
assign Jlj6x6 = (~(vis_r7_o[21] & L92ov6));
assign Clj6x6 = (~(vis_r6_o[21] & S92ov6));
assign Okj6x6 = (Qlj6x6 & Xlj6x6);
assign Xlj6x6 = (~(vis_r5_o[21] & Na2ov6));
assign Qlj6x6 = (~(vis_r4_o[21] & Ua2ov6));
assign Akj6x6 = (Emj6x6 & Lmj6x6);
assign Lmj6x6 = (Smj6x6 & Zmj6x6);
assign Zmj6x6 = (~(vis_r3_o[21] & Dc2ov6));
assign Smj6x6 = (~(vis_r2_o[21] & Kc2ov6));
assign Emj6x6 = (Gnj6x6 & Nnj6x6);
assign Nnj6x6 = (~(vis_r1_o[21] & Fd2ov6));
assign Gnj6x6 = (~(vis_r0_o[21] & Md2ov6));
assign Efj6x6 = (~(Td2ov6 & T8yiw6));
assign T8yiw6 = (Spyiw6 ? Uy97z6 : Gli7z6[21]);
assign Uy97z6 = (~(Unj6x6 & Boj6x6));
assign Boj6x6 = (~(Nqyiw6 & Rgynv6));
assign Unj6x6 = (Ioj6x6 & Poj6x6);
assign Poj6x6 = (~(Pdc7z6[21] & Ouyiw6));
assign Ioj6x6 = (~(Vuyiw6 & Woj6x6));
assign Woj6x6 = (~(Dpj6x6 & Kpj6x6));
assign Kpj6x6 = (Rpj6x6 & Ypj6x6);
assign Ypj6x6 = (Fqj6x6 & Mqj6x6);
assign Mqj6x6 = (Tqj6x6 & Arj6x6);
assign Arj6x6 = (~(Hrj6x6 & Uxyiw6));
assign Hrj6x6 = (Kxb7z6[21] & Orj6x6);
assign Tqj6x6 = (~(Vrj6x6 & Csj6x6));
assign Vrj6x6 = (~(Jsj6x6 & Quziw6));
assign Jsj6x6 = (Qsj6x6 & Xsj6x6);
assign Xsj6x6 = (Orj6x6 | Ninnv6);
assign Orj6x6 = (Etj6x6 | Rje7z6[21]);
assign Qsj6x6 = (~(Ofnnv6 & Etj6x6));
assign Fqj6x6 = (Ltj6x6 & Stj6x6);
assign Stj6x6 = (~(R6ziw6 & Rb3ov6));
assign Rb3ov6 = (Ph1jw6 ^ Dte7z6[1]);
assign Ph1jw6 = (T3cdt6 ? V1c7z6[29] : Lt3ov6);
assign Ltj6x6 = (~(J73ov6 & Yi3ov6));
assign Rpj6x6 = (Ztj6x6 & Guj6x6);
assign Guj6x6 = (Nuj6x6 & Uuj6x6);
assign Uuj6x6 = (~(F7ziw6 & Kb3ov6));
assign Nuj6x6 = (~(T0ziw6 & Rje7z6[21]));
assign Ztj6x6 = (Bvj6x6 & Ivj6x6);
assign Ivj6x6 = (Ryfov6 | Pvj6x6);
assign Bvj6x6 = (~(L0g7z6[21] & J2ziw6));
assign Dpj6x6 = (Wvj6x6 & Dwj6x6);
assign Dwj6x6 = (Kwj6x6 & Rwj6x6);
assign Rwj6x6 = (Ywj6x6 & Fxj6x6);
assign Fxj6x6 = (~(Cqf7z6[5] & Q2ziw6));
assign Ywj6x6 = (~(L0g7z6[5] & O1ziw6));
assign Kwj6x6 = (Mxj6x6 & Txj6x6);
assign Txj6x6 = (~(U4ziw6 & V1c7z6[21]));
assign Mxj6x6 = (~(Z3ziw6 & Fhc7z6[10]));
assign Wvj6x6 = (Ayj6x6 & C03ov6);
assign C03ov6 = (Hyj6x6 & Oyj6x6);
assign Oyj6x6 = (~(Vyj6x6 & L3nnv6));
assign Vyj6x6 = (~(S3nnv6 | Icziw6));
assign Hyj6x6 = (~(Czj6x6 & Ubziw6));
assign Czj6x6 = (~(L3nnv6 ^ S3nnv6));
assign S3nnv6 = (Jzj6x6 ^ Mennv6);
assign Jzj6x6 = (~(Qzj6x6 & Xzj6x6));
assign Xzj6x6 = (E0k6x6 & L0k6x6);
assign L0k6x6 = (S0k6x6 & Z0k6x6);
assign Z0k6x6 = (~(Yxf7z6[23] & Su0jw6));
assign S0k6x6 = (G1k6x6 & N1k6x6);
assign N1k6x6 = (~(Yxf7z6[21] & Nv0jw6));
assign G1k6x6 = (~(Yxf7z6[22] & Uv0jw6));
assign E0k6x6 = (U1k6x6 & B2k6x6);
assign B2k6x6 = (~(Yxf7z6[24] & Pw0jw6));
assign U1k6x6 = (~(I2k6x6 & Rdziw6));
assign Qzj6x6 = (P2k6x6 & W2k6x6);
assign W2k6x6 = (D3k6x6 & K3k6x6);
assign K3k6x6 = (~(Onf7z6[21] & My0jw6));
assign D3k6x6 = (R3k6x6 & Y3k6x6);
assign Y3k6x6 = (~(Hz0jw6 & Kxb7z6[21]));
assign R3k6x6 = (~(Oz0jw6 & Fhc7z6[21]));
assign P2k6x6 = (F4k6x6 & M4k6x6);
assign M4k6x6 = (~(Alf7z6[5] & J01jw6));
assign F4k6x6 = (~(Alf7z6[21] & Q01jw6));
assign L3nnv6 = (~(T4k6x6 ^ Tennv6));
assign T4k6x6 = (~(A5k6x6 & H5k6x6));
assign H5k6x6 = (~(Yxf7z6[5] & Laziw6));
assign A5k6x6 = (O5k6x6 & V5k6x6);
assign V5k6x6 = (~(Yxf7z6[21] & Gbziw6));
assign O5k6x6 = (~(Kxb7z6[21] & Nbziw6));
assign Ayj6x6 = (T7ziw6 & C6k6x6);
assign C6k6x6 = (~(Qeldt6 & Oztiw6));
assign Cej6x6 = (J6k6x6 & Q6k6x6);
assign Q6k6x6 = (~(Ve2ov6 & vis_pc_o[21]));
assign J6k6x6 = (~(Fhc7z6[21] & Cf2ov6));
assign A0z7v6 = (~(X6k6x6 & E7k6x6));
assign E7k6x6 = (L7k6x6 & S7k6x6);
assign S7k6x6 = (Eu9ov6 | Z7k6x6);
assign L7k6x6 = (G8k6x6 & N8k6x6);
assign N8k6x6 = (~(Gv9ov6 & Jayiw6));
assign G8k6x6 = (~(Uv9ov6 & Q0a7z6));
assign X6k6x6 = (U8k6x6 & B9k6x6);
assign B9k6x6 = (~(Pw9ov6 & Kxb7z6[13]));
assign U8k6x6 = (I9k6x6 & P9k6x6);
assign P9k6x6 = (~(Kx9ov6 & vis_pc_o[13]));
assign I9k6x6 = (~(Gli7z6[13] & Rx9ov6));
assign Tzy7v6 = (~(W9k6x6 & Dak6x6));
assign Dak6x6 = (Kak6x6 & Rak6x6);
assign Rak6x6 = (~(H02ov6 & Q0a7z6));
assign Kak6x6 = (Yak6x6 & Fbk6x6);
assign Fbk6x6 = (C12ov6 | Ygknv6);
assign Ygknv6 = (Mbk6x6 & Tbk6x6);
assign Tbk6x6 = (Ack6x6 & Hck6x6);
assign Hck6x6 = (Ock6x6 & Vck6x6);
assign Vck6x6 = (Cdk6x6 & Jdk6x6);
assign Jdk6x6 = (~(vis_psp_o[13] & N32ov6));
assign Cdk6x6 = (~(U32ov6 & Pic7z6[13]));
assign Ock6x6 = (Qdk6x6 & Xdk6x6);
assign Xdk6x6 = (~(vis_msp_o[13] & P42ov6));
assign Qdk6x6 = (~(vis_r12_o[13] & W42ov6));
assign Ack6x6 = (Eek6x6 & Lek6x6);
assign Lek6x6 = (Sek6x6 & Zek6x6);
assign Zek6x6 = (~(vis_r11_o[13] & F62ov6));
assign Sek6x6 = (~(vis_r10_o[13] & M62ov6));
assign Eek6x6 = (Gfk6x6 & Nfk6x6);
assign Nfk6x6 = (~(vis_r9_o[13] & H72ov6));
assign Gfk6x6 = (~(vis_r8_o[13] & O72ov6));
assign Mbk6x6 = (Ufk6x6 & Bgk6x6);
assign Bgk6x6 = (Igk6x6 & Pgk6x6);
assign Pgk6x6 = (Wgk6x6 & Dhk6x6);
assign Dhk6x6 = (~(vis_r7_o[13] & L92ov6));
assign Wgk6x6 = (~(vis_r6_o[13] & S92ov6));
assign Igk6x6 = (Khk6x6 & Rhk6x6);
assign Rhk6x6 = (~(vis_r5_o[13] & Na2ov6));
assign Khk6x6 = (~(vis_r4_o[13] & Ua2ov6));
assign Ufk6x6 = (Yhk6x6 & Fik6x6);
assign Fik6x6 = (Mik6x6 & Tik6x6);
assign Tik6x6 = (~(vis_r3_o[13] & Dc2ov6));
assign Mik6x6 = (~(vis_r2_o[13] & Kc2ov6));
assign Yhk6x6 = (Ajk6x6 & Hjk6x6);
assign Hjk6x6 = (~(vis_r1_o[13] & Fd2ov6));
assign Ajk6x6 = (~(vis_r0_o[13] & Md2ov6));
assign Yak6x6 = (~(Td2ov6 & Jayiw6));
assign Jayiw6 = (Spyiw6 ? Q0a7z6 : Gli7z6[13]);
assign Q0a7z6 = (~(Ojk6x6 & Vjk6x6));
assign Vjk6x6 = (~(Nqyiw6 & Fgznv6));
assign Ojk6x6 = (Ckk6x6 & Jkk6x6);
assign Jkk6x6 = (~(Pdc7z6[13] & Ouyiw6));
assign Ckk6x6 = (~(Vuyiw6 & Qkk6x6));
assign Qkk6x6 = (~(Xkk6x6 & Elk6x6));
assign Elk6x6 = (Llk6x6 & Slk6x6);
assign Slk6x6 = (Zlk6x6 & Gmk6x6);
assign Gmk6x6 = (Nmk6x6 & Ns3jw6);
assign Nmk6x6 = (~(Umk6x6 & Uxyiw6));
assign Umk6x6 = (Kxb7z6[13] & Bnk6x6);
assign Zlk6x6 = (Ink6x6 & Pnk6x6);
assign Pnk6x6 = (~(Wnk6x6 & Dok6x6));
assign Wnk6x6 = (~(Kok6x6 & Quziw6));
assign Kok6x6 = (Rok6x6 & Yok6x6);
assign Yok6x6 = (Bnk6x6 | Ninnv6);
assign Bnk6x6 = (Fpk6x6 | Rje7z6[13]);
assign Rok6x6 = (~(Ofnnv6 & Fpk6x6));
assign Ink6x6 = (~(Yi3ov6 & Ug3ov6));
assign Yi3ov6 = (Mpk6x6 ^ Dte7z6[1]);
assign Llk6x6 = (Tpk6x6 & Aqk6x6);
assign Aqk6x6 = (Hqk6x6 & Oqk6x6);
assign Oqk6x6 = (~(Nn3ov6 & C73ov6));
assign Nn3ov6 = (J7j6x6 ^ Dte7z6[1]);
assign J7j6x6 = (T3cdt6 ? V1c7z6[5] : Xs3ov6);
assign Hqk6x6 = (~(J73ov6 & Kb3ov6));
assign Kb3ov6 = (I2k6x6 ^ Dte7z6[1]);
assign I2k6x6 = (T3cdt6 ? V1c7z6[21] : Csj6x6);
assign Tpk6x6 = (Vqk6x6 & Crk6x6);
assign Crk6x6 = (~(T0ziw6 & Rje7z6[13]));
assign Vqk6x6 = (Ryfov6 | Jrk6x6);
assign Xkk6x6 = (Qrk6x6 & Xrk6x6);
assign Xrk6x6 = (Esk6x6 & Lsk6x6);
assign Lsk6x6 = (Ssk6x6 & Zsk6x6);
assign Zsk6x6 = (~(L0g7z6[13] & J2ziw6));
assign Ssk6x6 = (~(L0g7z6[29] & Q2ziw6));
assign Esk6x6 = (Gtk6x6 & Ntk6x6);
assign Ntk6x6 = (~(O1ziw6 & Onf7z6[13]));
assign Gtk6x6 = (~(U4ziw6 & Fhc7z6[13]));
assign Qrk6x6 = (Utk6x6 & Vz2ov6);
assign Vz2ov6 = (Buk6x6 & Iuk6x6);
assign Iuk6x6 = (~(Puk6x6 & H8nnv6));
assign Puk6x6 = (~(O8nnv6 | Icziw6));
assign Buk6x6 = (~(Wuk6x6 & Ubziw6));
assign Wuk6x6 = (~(H8nnv6 ^ O8nnv6));
assign O8nnv6 = (Dvk6x6 ^ Mennv6);
assign Dvk6x6 = (~(Kvk6x6 & Rvk6x6));
assign Rvk6x6 = (Yvk6x6 & Fwk6x6);
assign Fwk6x6 = (Mwk6x6 & Twk6x6);
assign Twk6x6 = (~(Su0jw6 & Yxf7z6[15]));
assign Mwk6x6 = (Axk6x6 & Hxk6x6);
assign Hxk6x6 = (~(Yxf7z6[13] & Nv0jw6));
assign Axk6x6 = (~(Yxf7z6[14] & Uv0jw6));
assign Yvk6x6 = (Oxk6x6 & Vxk6x6);
assign Vxk6x6 = (~(Yxf7z6[16] & Pw0jw6));
assign Oxk6x6 = (~(Mpk6x6 & Rdziw6));
assign Mpk6x6 = (T3cdt6 ? V1c7z6[13] : Dok6x6);
assign Kvk6x6 = (Cyk6x6 & Jyk6x6);
assign Jyk6x6 = (Qyk6x6 & Xyk6x6);
assign Xyk6x6 = (~(Onf7z6[13] & My0jw6));
assign Qyk6x6 = (Ezk6x6 & Lzk6x6);
assign Lzk6x6 = (~(Hz0jw6 & Kxb7z6[13]));
assign Ezk6x6 = (~(Oz0jw6 & Fhc7z6[13]));
assign Cyk6x6 = (Szk6x6 & Zzk6x6);
assign Zzk6x6 = (~(Onf7z6[29] & J01jw6));
assign Szk6x6 = (~(Alf7z6[13] & Q01jw6));
assign H8nnv6 = (~(G0l6x6 ^ Tennv6));
assign G0l6x6 = (~(N0l6x6 & U0l6x6));
assign U0l6x6 = (~(Yxf7z6[13] & Gbziw6));
assign N0l6x6 = (~(Kxb7z6[13] & Nbziw6));
assign Utk6x6 = (B1l6x6 & I1l6x6);
assign I1l6x6 = (~(Z3ziw6 & Fhc7z6[18]));
assign B1l6x6 = (~(Ovldt6 & Oztiw6));
assign W9k6x6 = (P1l6x6 & W1l6x6);
assign W1l6x6 = (~(Ve2ov6 & vis_pc_o[13]));
assign P1l6x6 = (~(Fhc7z6[13] & Cf2ov6));
assign Mzy7v6 = (~(D2l6x6 & K2l6x6));
assign K2l6x6 = (R2l6x6 & Y2l6x6);
assign Y2l6x6 = (Eu9ov6 | F3l6x6);
assign R2l6x6 = (M3l6x6 & T3l6x6);
assign T3l6x6 = (~(Gv9ov6 & Zbyiw6));
assign M3l6x6 = (~(Uv9ov6 & E2a7z6));
assign D2l6x6 = (A4l6x6 & H4l6x6);
assign H4l6x6 = (~(Pw9ov6 & Kxb7z6[6]));
assign A4l6x6 = (O4l6x6 & V4l6x6);
assign V4l6x6 = (~(Kx9ov6 & vis_pc_o[6]));
assign O4l6x6 = (~(Gli7z6[6] & Rx9ov6));
assign Fzy7v6 = (~(C5l6x6 & J5l6x6));
assign J5l6x6 = (Q5l6x6 & X5l6x6);
assign X5l6x6 = (~(H02ov6 & E2a7z6));
assign Q5l6x6 = (E6l6x6 & L6l6x6);
assign L6l6x6 = (C12ov6 | Qdjnv6);
assign Qdjnv6 = (S6l6x6 & Z6l6x6);
assign Z6l6x6 = (G7l6x6 & N7l6x6);
assign N7l6x6 = (U7l6x6 & B8l6x6);
assign B8l6x6 = (I8l6x6 & P8l6x6);
assign P8l6x6 = (~(vis_psp_o[6] & N32ov6));
assign I8l6x6 = (~(U32ov6 & Pic7z6[6]));
assign U7l6x6 = (W8l6x6 & D9l6x6);
assign D9l6x6 = (~(vis_msp_o[6] & P42ov6));
assign W8l6x6 = (~(vis_r12_o[6] & W42ov6));
assign G7l6x6 = (K9l6x6 & R9l6x6);
assign R9l6x6 = (Y9l6x6 & Fal6x6);
assign Fal6x6 = (~(vis_r11_o[6] & F62ov6));
assign Y9l6x6 = (~(vis_r10_o[6] & M62ov6));
assign K9l6x6 = (Mal6x6 & Tal6x6);
assign Tal6x6 = (~(vis_r9_o[6] & H72ov6));
assign Mal6x6 = (~(vis_r8_o[6] & O72ov6));
assign S6l6x6 = (Abl6x6 & Hbl6x6);
assign Hbl6x6 = (Obl6x6 & Vbl6x6);
assign Vbl6x6 = (Ccl6x6 & Jcl6x6);
assign Jcl6x6 = (~(vis_r7_o[6] & L92ov6));
assign Ccl6x6 = (~(vis_r6_o[6] & S92ov6));
assign Obl6x6 = (Qcl6x6 & Xcl6x6);
assign Xcl6x6 = (~(vis_r5_o[6] & Na2ov6));
assign Qcl6x6 = (~(vis_r4_o[6] & Ua2ov6));
assign Abl6x6 = (Edl6x6 & Ldl6x6);
assign Ldl6x6 = (Sdl6x6 & Zdl6x6);
assign Zdl6x6 = (~(vis_r3_o[6] & Dc2ov6));
assign Sdl6x6 = (~(vis_r2_o[6] & Kc2ov6));
assign Edl6x6 = (Gel6x6 & Nel6x6);
assign Nel6x6 = (~(vis_r1_o[6] & Fd2ov6));
assign Gel6x6 = (~(vis_r0_o[6] & Md2ov6));
assign E6l6x6 = (~(Td2ov6 & Zbyiw6));
assign Zbyiw6 = (Spyiw6 ? E2a7z6 : Gli7z6[6]);
assign E2a7z6 = (~(Uel6x6 & Bfl6x6));
assign Bfl6x6 = (~(Nqyiw6 & M80ov6));
assign Uel6x6 = (Ifl6x6 & Pfl6x6);
assign Pfl6x6 = (~(Pdc7z6[6] & Ouyiw6));
assign Ifl6x6 = (~(Vuyiw6 & Wfl6x6));
assign Wfl6x6 = (~(Dgl6x6 & Kgl6x6));
assign Kgl6x6 = (Rgl6x6 & Ygl6x6);
assign Ygl6x6 = (Fhl6x6 & Mhl6x6);
assign Mhl6x6 = (Thl6x6 & Ail6x6);
assign Ail6x6 = (~(Hil6x6 & Uxyiw6));
assign Hil6x6 = (Kxb7z6[6] & Oil6x6);
assign Thl6x6 = (~(Vil6x6 & Jm0jw6));
assign Vil6x6 = (Nob7z6[6] & Rslov6);
assign Fhl6x6 = (Cjl6x6 & Jjl6x6);
assign Jjl6x6 = (~(Nu3ov6 & Qjl6x6));
assign Qjl6x6 = (~(Xjl6x6 & Quziw6));
assign Xjl6x6 = (Ekl6x6 & Lkl6x6);
assign Lkl6x6 = (Oil6x6 | Ninnv6);
assign Oil6x6 = (Skl6x6 | Rje7z6[6]);
assign Ekl6x6 = (~(Ofnnv6 & Skl6x6));
assign Cjl6x6 = (~(Ol0jw6 & Ql3ov6));
assign Ol0jw6 = (Gg3ov6 & Zkl6x6);
assign Zkl6x6 = (Gll6x6 | Nll6x6);
assign Rgl6x6 = (Ull6x6 & Bml6x6);
assign Bml6x6 = (Iml6x6 & Pml6x6);
assign Pml6x6 = (~(Di3ov6 & C73ov6));
assign Iml6x6 = (~(Hzi6x6 & Ppb7z6[6]));
assign Ull6x6 = (Wml6x6 & Dnl6x6);
assign Dnl6x6 = (~(T0ziw6 & Rje7z6[6]));
assign Wml6x6 = (Ryfov6 | Knl6x6);
assign Dgl6x6 = (Rnl6x6 & Ynl6x6);
assign Ynl6x6 = (Fol6x6 & Mol6x6);
assign Mol6x6 = (Tol6x6 & Apl6x6);
assign Apl6x6 = (~(J73ov6 & Je3ov6));
assign Tol6x6 = (~(L0g7z6[6] & J2ziw6));
assign Fol6x6 = (Hpl6x6 & Opl6x6);
assign Opl6x6 = (~(L0g7z6[22] & Q2ziw6));
assign Hpl6x6 = (~(O1ziw6 & Onf7z6[6]));
assign Rnl6x6 = (Vpl6x6 & Cql6x6);
assign Cql6x6 = (Jql6x6 & Qql6x6);
assign Qql6x6 = (~(U4ziw6 & Fhc7z6[6]));
assign Jql6x6 = (~(Z3ziw6 & Fhc7z6[25]));
assign Vpl6x6 = (Q03ov6 & Xql6x6);
assign Xql6x6 = (~(Jamdt6 & Oztiw6));
assign Q03ov6 = (Erl6x6 & Lrl6x6);
assign Lrl6x6 = (~(Srl6x6 & Xvmnv6));
assign Srl6x6 = (~(Ewmnv6 | Icziw6));
assign Erl6x6 = (~(Zrl6x6 & Ubziw6));
assign Zrl6x6 = (~(Xvmnv6 ^ Ewmnv6));
assign Ewmnv6 = (Gsl6x6 ^ Mennv6);
assign Gsl6x6 = (~(Nsl6x6 & Usl6x6));
assign Usl6x6 = (Btl6x6 & Itl6x6);
assign Itl6x6 = (Ptl6x6 & Wtl6x6);
assign Wtl6x6 = (~(Yxf7z6[8] & Su0jw6));
assign Ptl6x6 = (Dul6x6 & Kul6x6);
assign Kul6x6 = (~(Yxf7z6[6] & Nv0jw6));
assign Dul6x6 = (~(Yxf7z6[7] & Uv0jw6));
assign Btl6x6 = (Rul6x6 & Yul6x6);
assign Yul6x6 = (~(Yxf7z6[9] & Pw0jw6));
assign Rul6x6 = (~(Fvl6x6 & Rdziw6));
assign Nsl6x6 = (Mvl6x6 & Tvl6x6);
assign Tvl6x6 = (Awl6x6 & Hwl6x6);
assign Hwl6x6 = (~(Onf7z6[6] & My0jw6));
assign Awl6x6 = (Owl6x6 & Vwl6x6);
assign Vwl6x6 = (~(Hz0jw6 & Kxb7z6[6]));
assign Owl6x6 = (~(Oz0jw6 & Fhc7z6[6]));
assign Mvl6x6 = (Cxl6x6 & Jxl6x6);
assign Jxl6x6 = (~(Onf7z6[22] & J01jw6));
assign Cxl6x6 = (~(Alf7z6[6] & Q01jw6));
assign Xvmnv6 = (~(Qxl6x6 ^ Tennv6));
assign Qxl6x6 = (~(Xxl6x6 & Eyl6x6));
assign Eyl6x6 = (~(Yxf7z6[6] & Gbziw6));
assign Xxl6x6 = (~(Kxb7z6[6] & Nbziw6));
assign C5l6x6 = (Lyl6x6 & Syl6x6);
assign Syl6x6 = (~(Ve2ov6 & vis_pc_o[6]));
assign Lyl6x6 = (~(Fhc7z6[6] & Cf2ov6));
assign Yyy7v6 = (~(Zyl6x6 & Gzl6x6));
assign Gzl6x6 = (Nzl6x6 & Uzl6x6);
assign Uzl6x6 = (Eu9ov6 | B0m6x6);
assign Nzl6x6 = (I0m6x6 & P0m6x6);
assign P0m6x6 = (~(Gv9ov6 & M8yiw6));
assign I0m6x6 = (~(Uv9ov6 & My97z6));
assign Zyl6x6 = (W0m6x6 & D1m6x6);
assign D1m6x6 = (~(Pw9ov6 & Kxb7z6[22]));
assign W0m6x6 = (K1m6x6 & R1m6x6);
assign R1m6x6 = (~(Kx9ov6 & vis_pc_o[22]));
assign K1m6x6 = (~(Gli7z6[22] & Rx9ov6));
assign Ryy7v6 = (~(Y1m6x6 & F2m6x6));
assign F2m6x6 = (M2m6x6 & T2m6x6);
assign T2m6x6 = (~(H02ov6 & My97z6));
assign M2m6x6 = (A3m6x6 & H3m6x6);
assign H3m6x6 = (C12ov6 | G0knv6);
assign G0knv6 = (O3m6x6 & V3m6x6);
assign V3m6x6 = (C4m6x6 & J4m6x6);
assign J4m6x6 = (Q4m6x6 & X4m6x6);
assign X4m6x6 = (E5m6x6 & L5m6x6);
assign L5m6x6 = (~(vis_psp_o[22] & N32ov6));
assign E5m6x6 = (~(U32ov6 & Pic7z6[22]));
assign Q4m6x6 = (S5m6x6 & Z5m6x6);
assign Z5m6x6 = (~(vis_msp_o[22] & P42ov6));
assign S5m6x6 = (~(vis_r12_o[22] & W42ov6));
assign C4m6x6 = (G6m6x6 & N6m6x6);
assign N6m6x6 = (U6m6x6 & B7m6x6);
assign B7m6x6 = (~(vis_r11_o[22] & F62ov6));
assign U6m6x6 = (~(vis_r10_o[22] & M62ov6));
assign G6m6x6 = (I7m6x6 & P7m6x6);
assign P7m6x6 = (~(vis_r9_o[22] & H72ov6));
assign I7m6x6 = (~(vis_r8_o[22] & O72ov6));
assign O3m6x6 = (W7m6x6 & D8m6x6);
assign D8m6x6 = (K8m6x6 & R8m6x6);
assign R8m6x6 = (Y8m6x6 & F9m6x6);
assign F9m6x6 = (~(vis_r7_o[22] & L92ov6));
assign Y8m6x6 = (~(vis_r6_o[22] & S92ov6));
assign K8m6x6 = (M9m6x6 & T9m6x6);
assign T9m6x6 = (~(vis_r5_o[22] & Na2ov6));
assign M9m6x6 = (~(vis_r4_o[22] & Ua2ov6));
assign W7m6x6 = (Aam6x6 & Ham6x6);
assign Ham6x6 = (Oam6x6 & Vam6x6);
assign Vam6x6 = (~(vis_r3_o[22] & Dc2ov6));
assign Oam6x6 = (~(vis_r2_o[22] & Kc2ov6));
assign Aam6x6 = (Cbm6x6 & Jbm6x6);
assign Jbm6x6 = (~(vis_r1_o[22] & Fd2ov6));
assign Cbm6x6 = (~(vis_r0_o[22] & Md2ov6));
assign A3m6x6 = (~(Td2ov6 & M8yiw6));
assign M8yiw6 = (Spyiw6 ? My97z6 : Gli7z6[22]);
assign My97z6 = (~(Qbm6x6 & Xbm6x6));
assign Xbm6x6 = (~(Nqyiw6 & Ccynv6));
assign Qbm6x6 = (Ecm6x6 & Lcm6x6);
assign Lcm6x6 = (~(Pdc7z6[22] & Ouyiw6));
assign Ecm6x6 = (~(Vuyiw6 & Scm6x6));
assign Scm6x6 = (~(Zcm6x6 & Gdm6x6));
assign Gdm6x6 = (Ndm6x6 & Udm6x6);
assign Udm6x6 = (Bem6x6 & Iem6x6);
assign Iem6x6 = (Pem6x6 & Wem6x6);
assign Wem6x6 = (~(Dfm6x6 & Uxyiw6));
assign Dfm6x6 = (Kxb7z6[22] & Kfm6x6);
assign Pem6x6 = (~(Rfm6x6 & Yfm6x6));
assign Rfm6x6 = (~(Fgm6x6 & Quziw6));
assign Fgm6x6 = (Mgm6x6 & Tgm6x6);
assign Tgm6x6 = (Kfm6x6 | Ninnv6);
assign Kfm6x6 = (Ahm6x6 | Rje7z6[22]);
assign Mgm6x6 = (~(Ofnnv6 & Ahm6x6));
assign Bem6x6 = (Hhm6x6 & Ohm6x6);
assign Ohm6x6 = (~(J73ov6 & Di3ov6));
assign Hhm6x6 = (~(T0ziw6 & Rje7z6[22]));
assign Ndm6x6 = (Vhm6x6 & Cim6x6);
assign Cim6x6 = (Jim6x6 & Qim6x6);
assign Qim6x6 = (Ryfov6 | Xim6x6);
assign Jim6x6 = (~(L0g7z6[22] & J2ziw6));
assign Vhm6x6 = (Ejm6x6 & Ljm6x6);
assign Ljm6x6 = (~(R6ziw6 & Je3ov6));
assign Ejm6x6 = (~(F7ziw6 & Qe3ov6));
assign Zcm6x6 = (Sjm6x6 & Zjm6x6);
assign Zjm6x6 = (Gkm6x6 & Nkm6x6);
assign Nkm6x6 = (Ukm6x6 & Blm6x6);
assign Blm6x6 = (~(Cqf7z6[6] & Q2ziw6));
assign Ukm6x6 = (~(L0g7z6[6] & O1ziw6));
assign Gkm6x6 = (Ilm6x6 & Plm6x6);
assign Plm6x6 = (~(U4ziw6 & V1c7z6[22]));
assign Ilm6x6 = (~(Z3ziw6 & Fhc7z6[9]));
assign Sjm6x6 = (Wlm6x6 & J03ov6);
assign J03ov6 = (Dmm6x6 & Kmm6x6);
assign Kmm6x6 = (~(Rmm6x6 & X2nnv6));
assign Rmm6x6 = (~(E3nnv6 | Icziw6));
assign Dmm6x6 = (~(Ymm6x6 & Ubziw6));
assign Ymm6x6 = (~(X2nnv6 ^ E3nnv6));
assign E3nnv6 = (Fnm6x6 ^ Mennv6);
assign Fnm6x6 = (~(Mnm6x6 & Tnm6x6));
assign Tnm6x6 = (Aom6x6 & Hom6x6);
assign Hom6x6 = (Oom6x6 & Vom6x6);
assign Vom6x6 = (~(Yxf7z6[24] & Su0jw6));
assign Oom6x6 = (Cpm6x6 & Jpm6x6);
assign Jpm6x6 = (~(Yxf7z6[22] & Nv0jw6));
assign Cpm6x6 = (~(Yxf7z6[23] & Uv0jw6));
assign Aom6x6 = (Qpm6x6 & Xpm6x6);
assign Xpm6x6 = (~(Yxf7z6[25] & Pw0jw6));
assign Qpm6x6 = (~(Eqm6x6 & Rdziw6));
assign Mnm6x6 = (Lqm6x6 & Sqm6x6);
assign Sqm6x6 = (Zqm6x6 & Grm6x6);
assign Grm6x6 = (~(Onf7z6[22] & My0jw6));
assign Zqm6x6 = (Nrm6x6 & Urm6x6);
assign Urm6x6 = (~(Hz0jw6 & Kxb7z6[22]));
assign Nrm6x6 = (~(Oz0jw6 & Fhc7z6[22]));
assign Lqm6x6 = (Bsm6x6 & Ism6x6);
assign Ism6x6 = (~(Alf7z6[6] & J01jw6));
assign Bsm6x6 = (~(Alf7z6[22] & Q01jw6));
assign X2nnv6 = (~(Psm6x6 ^ Tennv6));
assign Psm6x6 = (~(Wsm6x6 & Dtm6x6));
assign Dtm6x6 = (~(Yxf7z6[6] & Laziw6));
assign Wsm6x6 = (Ktm6x6 & Rtm6x6);
assign Rtm6x6 = (~(Yxf7z6[22] & Gbziw6));
assign Ktm6x6 = (~(Kxb7z6[22] & Nbziw6));
assign Wlm6x6 = (T7ziw6 & Ytm6x6);
assign Ytm6x6 = (~(Ncldt6 & Oztiw6));
assign Y1m6x6 = (Fum6x6 & Mum6x6);
assign Mum6x6 = (~(Ve2ov6 & vis_pc_o[22]));
assign Fum6x6 = (~(Fhc7z6[22] & Cf2ov6));
assign Kyy7v6 = (~(Tum6x6 & Avm6x6));
assign Avm6x6 = (Hvm6x6 & Ovm6x6);
assign Ovm6x6 = (Eu9ov6 | Vvm6x6);
assign Hvm6x6 = (Cwm6x6 & Jwm6x6);
assign Jwm6x6 = (~(Gv9ov6 & Cayiw6));
assign Cwm6x6 = (~(Uv9ov6 & I0a7z6));
assign Tum6x6 = (Qwm6x6 & Xwm6x6);
assign Xwm6x6 = (~(Pw9ov6 & Kxb7z6[14]));
assign Qwm6x6 = (Exm6x6 & Lxm6x6);
assign Lxm6x6 = (~(Kx9ov6 & vis_pc_o[14]));
assign Exm6x6 = (~(Gli7z6[14] & Rx9ov6));
assign Dyy7v6 = (~(Sxm6x6 & Zxm6x6));
assign Zxm6x6 = (Gym6x6 & Nym6x6);
assign Nym6x6 = (~(H02ov6 & I0a7z6));
assign Gym6x6 = (Uym6x6 & Bzm6x6);
assign Bzm6x6 = (C12ov6 | Ifknv6);
assign Ifknv6 = (Izm6x6 & Pzm6x6);
assign Pzm6x6 = (Wzm6x6 & D0n6x6);
assign D0n6x6 = (K0n6x6 & R0n6x6);
assign R0n6x6 = (Y0n6x6 & F1n6x6);
assign F1n6x6 = (~(vis_psp_o[14] & N32ov6));
assign Y0n6x6 = (~(U32ov6 & Pic7z6[14]));
assign K0n6x6 = (M1n6x6 & T1n6x6);
assign T1n6x6 = (~(vis_msp_o[14] & P42ov6));
assign M1n6x6 = (~(vis_r12_o[14] & W42ov6));
assign Wzm6x6 = (A2n6x6 & H2n6x6);
assign H2n6x6 = (O2n6x6 & V2n6x6);
assign V2n6x6 = (~(vis_r11_o[14] & F62ov6));
assign O2n6x6 = (~(vis_r10_o[14] & M62ov6));
assign A2n6x6 = (C3n6x6 & J3n6x6);
assign J3n6x6 = (~(vis_r9_o[14] & H72ov6));
assign C3n6x6 = (~(vis_r8_o[14] & O72ov6));
assign Izm6x6 = (Q3n6x6 & X3n6x6);
assign X3n6x6 = (E4n6x6 & L4n6x6);
assign L4n6x6 = (S4n6x6 & Z4n6x6);
assign Z4n6x6 = (~(vis_r7_o[14] & L92ov6));
assign S4n6x6 = (~(vis_r6_o[14] & S92ov6));
assign E4n6x6 = (G5n6x6 & N5n6x6);
assign N5n6x6 = (~(vis_r5_o[14] & Na2ov6));
assign G5n6x6 = (~(vis_r4_o[14] & Ua2ov6));
assign Q3n6x6 = (U5n6x6 & B6n6x6);
assign B6n6x6 = (I6n6x6 & P6n6x6);
assign P6n6x6 = (~(vis_r3_o[14] & Dc2ov6));
assign I6n6x6 = (~(vis_r2_o[14] & Kc2ov6));
assign U5n6x6 = (W6n6x6 & D7n6x6);
assign D7n6x6 = (~(vis_r1_o[14] & Fd2ov6));
assign W6n6x6 = (~(vis_r0_o[14] & Md2ov6));
assign Uym6x6 = (~(Td2ov6 & Cayiw6));
assign Cayiw6 = (Spyiw6 ? I0a7z6 : Gli7z6[14]);
assign I0a7z6 = (~(K7n6x6 & R7n6x6));
assign R7n6x6 = (~(Nqyiw6 & Ecznv6));
assign K7n6x6 = (Y7n6x6 & F8n6x6);
assign F8n6x6 = (~(Pdc7z6[14] & Ouyiw6));
assign Y7n6x6 = (~(Vuyiw6 & M8n6x6));
assign M8n6x6 = (~(T8n6x6 & A9n6x6));
assign A9n6x6 = (H9n6x6 & O9n6x6);
assign O9n6x6 = (V9n6x6 & Can6x6);
assign Can6x6 = (Jan6x6 & Ns3jw6);
assign Jan6x6 = (~(Qan6x6 & Uxyiw6));
assign Qan6x6 = (Kxb7z6[14] & Xan6x6);
assign V9n6x6 = (Ebn6x6 & Lbn6x6);
assign Lbn6x6 = (~(Sbn6x6 & Zbn6x6));
assign Sbn6x6 = (~(Gcn6x6 & Quziw6));
assign Gcn6x6 = (Ncn6x6 & Ucn6x6);
assign Ucn6x6 = (Xan6x6 | Ninnv6);
assign Xan6x6 = (Bdn6x6 | Rje7z6[14]);
assign Ncn6x6 = (~(Ofnnv6 & Bdn6x6));
assign Ebn6x6 = (~(Di3ov6 & Ug3ov6));
assign Di3ov6 = (Idn6x6 ^ Dte7z6[1]);
assign H9n6x6 = (Pdn6x6 & Wdn6x6);
assign Wdn6x6 = (Den6x6 & Ken6x6);
assign Ken6x6 = (~(Ql3ov6 & C73ov6));
assign Den6x6 = (~(T0ziw6 & Rje7z6[14]));
assign Pdn6x6 = (Ren6x6 & Yen6x6);
assign Yen6x6 = (Ryfov6 | Ffn6x6);
assign Ren6x6 = (~(J73ov6 & Qe3ov6));
assign T8n6x6 = (Mfn6x6 & Tfn6x6);
assign Tfn6x6 = (Agn6x6 & Hgn6x6);
assign Hgn6x6 = (Ogn6x6 & Vgn6x6);
assign Vgn6x6 = (~(L0g7z6[14] & J2ziw6));
assign Ogn6x6 = (~(L0g7z6[30] & Q2ziw6));
assign Agn6x6 = (Chn6x6 & Jhn6x6);
assign Jhn6x6 = (~(O1ziw6 & Onf7z6[14]));
assign Chn6x6 = (~(U4ziw6 & Fhc7z6[14]));
assign Mfn6x6 = (Qhn6x6 & G23ov6);
assign G23ov6 = (Xhn6x6 & Ein6x6);
assign Ein6x6 = (~(Lin6x6 & T7nnv6));
assign Lin6x6 = (~(A8nnv6 | Icziw6));
assign Xhn6x6 = (~(Sin6x6 & Ubziw6));
assign Sin6x6 = (~(T7nnv6 ^ A8nnv6));
assign A8nnv6 = (Zin6x6 ^ Mennv6);
assign Zin6x6 = (~(Gjn6x6 & Njn6x6));
assign Njn6x6 = (Ujn6x6 & Bkn6x6);
assign Bkn6x6 = (Ikn6x6 & Pkn6x6);
assign Pkn6x6 = (~(Yxf7z6[16] & Su0jw6));
assign Ikn6x6 = (Wkn6x6 & Dln6x6);
assign Dln6x6 = (~(Yxf7z6[14] & Nv0jw6));
assign Wkn6x6 = (~(Uv0jw6 & Yxf7z6[15]));
assign Ujn6x6 = (Kln6x6 & Rln6x6);
assign Rln6x6 = (~(Yxf7z6[17] & Pw0jw6));
assign Kln6x6 = (~(Idn6x6 & Rdziw6));
assign Idn6x6 = (T3cdt6 ? V1c7z6[14] : Zbn6x6);
assign Gjn6x6 = (Yln6x6 & Fmn6x6);
assign Fmn6x6 = (Mmn6x6 & Tmn6x6);
assign Tmn6x6 = (~(Onf7z6[14] & My0jw6));
assign Mmn6x6 = (Ann6x6 & Hnn6x6);
assign Hnn6x6 = (~(Hz0jw6 & Kxb7z6[14]));
assign Ann6x6 = (~(Oz0jw6 & Fhc7z6[14]));
assign Yln6x6 = (Onn6x6 & Vnn6x6);
assign Vnn6x6 = (~(Onf7z6[30] & J01jw6));
assign Onn6x6 = (~(Alf7z6[14] & Q01jw6));
assign T7nnv6 = (~(Con6x6 ^ Tennv6));
assign Con6x6 = (~(Jon6x6 & Qon6x6));
assign Qon6x6 = (~(Yxf7z6[14] & Gbziw6));
assign Jon6x6 = (~(Kxb7z6[14] & Nbziw6));
assign Qhn6x6 = (Xon6x6 & Epn6x6);
assign Epn6x6 = (~(Z3ziw6 & Fhc7z6[17]));
assign Xon6x6 = (~(Ltldt6 & Oztiw6));
assign Sxm6x6 = (Lpn6x6 & Spn6x6);
assign Spn6x6 = (~(Ve2ov6 & vis_pc_o[14]));
assign Lpn6x6 = (~(Fhc7z6[14] & Cf2ov6));
assign Wxy7v6 = (~(Zpn6x6 & Gqn6x6));
assign Gqn6x6 = (Nqn6x6 & Uqn6x6);
assign Uqn6x6 = (Eu9ov6 | Brn6x6);
assign Nqn6x6 = (Irn6x6 & Prn6x6);
assign Prn6x6 = (~(Gv9ov6 & Sbyiw6));
assign Irn6x6 = (~(Uv9ov6 & W1a7z6));
assign Zpn6x6 = (Wrn6x6 & Dsn6x6);
assign Dsn6x6 = (~(Pw9ov6 & Kxb7z6[7]));
assign Wrn6x6 = (Ksn6x6 & Rsn6x6);
assign Rsn6x6 = (~(Kx9ov6 & vis_pc_o[7]));
assign Ksn6x6 = (~(Gli7z6[7] & Rx9ov6));
assign Pxy7v6 = (~(Ysn6x6 & Ftn6x6));
assign Ftn6x6 = (Mtn6x6 & Ttn6x6);
assign Ttn6x6 = (~(Cuziw6 & C6bov6));
assign Mtn6x6 = (~(J6bov6 & Alf7z6[0]));
assign Ysn6x6 = (Aun6x6 & Hun6x6);
assign Hun6x6 = (~(L0g7z6[16] & E7bov6));
assign Aun6x6 = (~(L0g7z6[0] & L7bov6));
assign Ixy7v6 = (~(Oun6x6 & Vun6x6));
assign Vun6x6 = (Cvn6x6 & Jvn6x6);
assign Jvn6x6 = (~(H02ov6 & W1a7z6));
assign Cvn6x6 = (Qvn6x6 & Xvn6x6);
assign Xvn6x6 = (C12ov6 | Acjnv6);
assign Acjnv6 = (Ewn6x6 & Lwn6x6);
assign Lwn6x6 = (Swn6x6 & Zwn6x6);
assign Zwn6x6 = (Gxn6x6 & Nxn6x6);
assign Nxn6x6 = (Uxn6x6 & Byn6x6);
assign Byn6x6 = (~(vis_psp_o[7] & N32ov6));
assign Uxn6x6 = (~(U32ov6 & Pic7z6[7]));
assign Gxn6x6 = (Iyn6x6 & Pyn6x6);
assign Pyn6x6 = (~(vis_msp_o[7] & P42ov6));
assign Iyn6x6 = (~(vis_r12_o[7] & W42ov6));
assign Swn6x6 = (Wyn6x6 & Dzn6x6);
assign Dzn6x6 = (Kzn6x6 & Rzn6x6);
assign Rzn6x6 = (~(vis_r11_o[7] & F62ov6));
assign Kzn6x6 = (~(vis_r10_o[7] & M62ov6));
assign Wyn6x6 = (Yzn6x6 & F0o6x6);
assign F0o6x6 = (~(vis_r9_o[7] & H72ov6));
assign Yzn6x6 = (~(vis_r8_o[7] & O72ov6));
assign Ewn6x6 = (M0o6x6 & T0o6x6);
assign T0o6x6 = (A1o6x6 & H1o6x6);
assign H1o6x6 = (O1o6x6 & V1o6x6);
assign V1o6x6 = (~(vis_r7_o[7] & L92ov6));
assign O1o6x6 = (~(vis_r6_o[7] & S92ov6));
assign A1o6x6 = (C2o6x6 & J2o6x6);
assign J2o6x6 = (~(vis_r5_o[7] & Na2ov6));
assign C2o6x6 = (~(vis_r4_o[7] & Ua2ov6));
assign M0o6x6 = (Q2o6x6 & X2o6x6);
assign X2o6x6 = (E3o6x6 & L3o6x6);
assign L3o6x6 = (~(vis_r3_o[7] & Dc2ov6));
assign E3o6x6 = (~(vis_r2_o[7] & Kc2ov6));
assign Q2o6x6 = (S3o6x6 & Z3o6x6);
assign Z3o6x6 = (~(vis_r1_o[7] & Fd2ov6));
assign S3o6x6 = (~(vis_r0_o[7] & Md2ov6));
assign Qvn6x6 = (~(Td2ov6 & Sbyiw6));
assign Sbyiw6 = (Spyiw6 ? W1a7z6 : Gli7z6[7]);
assign W1a7z6 = (~(G4o6x6 & N4o6x6));
assign N4o6x6 = (~(Nqyiw6 & L40ov6));
assign G4o6x6 = (U4o6x6 & B5o6x6);
assign B5o6x6 = (~(Pdc7z6[7] & Ouyiw6));
assign U4o6x6 = (~(Vuyiw6 & I5o6x6));
assign I5o6x6 = (~(P5o6x6 & W5o6x6));
assign W5o6x6 = (D6o6x6 & K6o6x6);
assign K6o6x6 = (R6o6x6 & Y6o6x6);
assign Y6o6x6 = (F7o6x6 & M7o6x6);
assign M7o6x6 = (~(T7o6x6 & Uxyiw6));
assign T7o6x6 = (Kxb7z6[7] & A8o6x6);
assign F7o6x6 = (~(Bv3ov6 & H8o6x6));
assign H8o6x6 = (~(O8o6x6 & Quziw6));
assign O8o6x6 = (V8o6x6 & C9o6x6);
assign C9o6x6 = (A8o6x6 | Ninnv6);
assign A8o6x6 = (J9o6x6 | Rje7z6[7]);
assign V8o6x6 = (~(Ofnnv6 & J9o6x6));
assign R6o6x6 = (Q9o6x6 & X9o6x6);
assign X9o6x6 = (~(Hzi6x6 & Ppb7z6[7]));
assign Hzi6x6 = (Eao6x6 & C1gov6);
assign C1gov6 = (Lao6x6 & Dte7z6[16]);
assign Lao6x6 = (Sao6x6 & Msziw6);
assign Eao6x6 = (~(Zao6x6 | Gbo6x6));
assign Q9o6x6 = (~(Ok3ov6 & C73ov6));
assign C73ov6 = (~(Zf3ov6 & Nbo6x6));
assign Nbo6x6 = (Ubo6x6 | Bi2ov6);
assign D6o6x6 = (Bco6x6 & Ico6x6);
assign Ico6x6 = (Pco6x6 & Wco6x6);
assign Wco6x6 = (~(Jm0jw6 & Ddo6x6));
assign Jm0jw6 = (Kdo6x6 & Dte7z6[14]);
assign Pco6x6 = (~(T0ziw6 & Rje7z6[7]));
assign Bco6x6 = (Rdo6x6 & Ydo6x6);
assign Ydo6x6 = (Ryfov6 | Feo6x6);
assign Feo6x6 = (!J9o6x6);
assign Rdo6x6 = (~(L0g7z6[7] & J2ziw6));
assign P5o6x6 = (Meo6x6 & Teo6x6);
assign Teo6x6 = (Afo6x6 & Hfo6x6);
assign Hfo6x6 = (Ofo6x6 & Vfo6x6);
assign Vfo6x6 = (~(L0g7z6[23] & Q2ziw6));
assign Ofo6x6 = (~(O1ziw6 & Onf7z6[7]));
assign Afo6x6 = (Cgo6x6 & Jgo6x6);
assign Jgo6x6 = (~(U4ziw6 & Fhc7z6[7]));
assign Cgo6x6 = (~(Z3ziw6 & Fhc7z6[24]));
assign Meo6x6 = (Qgo6x6 & Wo3ov6);
assign Wo3ov6 = (Xgo6x6 & Eho6x6);
assign Eho6x6 = (~(J73ov6 & M7ziw6));
assign Xgo6x6 = (Lho6x6 & Ns3jw6);
assign Ns3jw6 = (~(Nll6x6 & H8ziw6));
assign Lho6x6 = (~(H8ziw6 & Gll6x6));
assign Gll6x6 = (Ug3ov6 | Ubo6x6);
assign Ug3ov6 = (~(Sf3ov6 & Sho6x6));
assign Sho6x6 = (~(Zho6x6 & Ubo6x6));
assign Sf3ov6 = (!F7ziw6);
assign Qgo6x6 = (Z13ov6 & Gio6x6);
assign Gio6x6 = (~(G8mdt6 & Oztiw6));
assign Z13ov6 = (Nio6x6 & Uio6x6);
assign Uio6x6 = (~(Bjo6x6 & Jvmnv6));
assign Bjo6x6 = (~(Qvmnv6 | Icziw6));
assign Nio6x6 = (~(Ijo6x6 & Ubziw6));
assign Ijo6x6 = (~(Jvmnv6 ^ Qvmnv6));
assign Qvmnv6 = (Pjo6x6 ^ Mennv6);
assign Pjo6x6 = (~(Wjo6x6 & Dko6x6));
assign Dko6x6 = (Kko6x6 & Rko6x6);
assign Rko6x6 = (Yko6x6 & Flo6x6);
assign Flo6x6 = (~(Yxf7z6[9] & Su0jw6));
assign Yko6x6 = (Mlo6x6 & Tlo6x6);
assign Tlo6x6 = (~(Yxf7z6[7] & Nv0jw6));
assign Mlo6x6 = (~(Yxf7z6[8] & Uv0jw6));
assign Kko6x6 = (Amo6x6 & Hmo6x6);
assign Hmo6x6 = (~(Yxf7z6[10] & Pw0jw6));
assign Amo6x6 = (~(Hz0jw6 & Kxb7z6[7]));
assign Wjo6x6 = (Omo6x6 & Vmo6x6);
assign Vmo6x6 = (Cno6x6 & Jno6x6);
assign Jno6x6 = (~(Onf7z6[23] & J01jw6));
assign Cno6x6 = (Qno6x6 & Xno6x6);
assign Xno6x6 = (~(Oz0jw6 & Fhc7z6[7]));
assign Qno6x6 = (~(Onf7z6[7] & My0jw6));
assign Omo6x6 = (Eoo6x6 & Loo6x6);
assign Loo6x6 = (~(Soo6x6 & Rdziw6));
assign Eoo6x6 = (~(Alf7z6[7] & Q01jw6));
assign Jvmnv6 = (~(Zoo6x6 ^ Tennv6));
assign Zoo6x6 = (~(Gpo6x6 & Npo6x6));
assign Npo6x6 = (~(Yxf7z6[7] & Gbziw6));
assign Gpo6x6 = (~(Kxb7z6[7] & Nbziw6));
assign Oun6x6 = (Upo6x6 & Bqo6x6);
assign Bqo6x6 = (~(Ve2ov6 & vis_pc_o[7]));
assign Upo6x6 = (~(Fhc7z6[7] & Cf2ov6));
assign Bxy7v6 = (~(Iqo6x6 & Pqo6x6));
assign Pqo6x6 = (Wqo6x6 & Dro6x6);
assign Dro6x6 = (~(St3ov6 & C6bov6));
assign Wqo6x6 = (~(J6bov6 & Alf7z6[27]));
assign Iqo6x6 = (Kro6x6 & Rro6x6);
assign Rro6x6 = (~(Cqf7z6[11] & E7bov6));
assign Kro6x6 = (~(L0g7z6[27] & L7bov6));
assign Uwy7v6 = (~(Yro6x6 & Fso6x6));
assign Fso6x6 = (Mso6x6 & Tso6x6);
assign Tso6x6 = (~(Qs3ov6 & C6bov6));
assign Mso6x6 = (~(J6bov6 & Alf7z6[26]));
assign Yro6x6 = (Ato6x6 & Hto6x6);
assign Hto6x6 = (~(Cqf7z6[10] & E7bov6));
assign Ato6x6 = (~(L0g7z6[26] & L7bov6));
assign Nwy7v6 = (~(Oto6x6 & Vto6x6));
assign Vto6x6 = (Cuo6x6 & Juo6x6);
assign Juo6x6 = (Eu9ov6 | Quo6x6);
assign Cuo6x6 = (Xuo6x6 & Evo6x6);
assign Evo6x6 = (~(Gv9ov6 & F8yiw6));
assign Xuo6x6 = (~(Uv9ov6 & Ey97z6));
assign Oto6x6 = (Lvo6x6 & Svo6x6);
assign Svo6x6 = (~(Pw9ov6 & Kxb7z6[23]));
assign Lvo6x6 = (Zvo6x6 & Gwo6x6);
assign Gwo6x6 = (~(Kx9ov6 & vis_pc_o[23]));
assign Zvo6x6 = (~(Gli7z6[23] & Rx9ov6));
assign Gwy7v6 = (~(Nwo6x6 & Uwo6x6));
assign Uwo6x6 = (Bxo6x6 & Ixo6x6);
assign Ixo6x6 = (~(H02ov6 & Ey97z6));
assign Bxo6x6 = (Pxo6x6 & Wxo6x6);
assign Wxo6x6 = (C12ov6 | Qyjnv6);
assign Qyjnv6 = (Dyo6x6 & Kyo6x6);
assign Kyo6x6 = (Ryo6x6 & Yyo6x6);
assign Yyo6x6 = (Fzo6x6 & Mzo6x6);
assign Mzo6x6 = (Tzo6x6 & A0p6x6);
assign A0p6x6 = (~(vis_psp_o[23] & N32ov6));
assign Tzo6x6 = (~(U32ov6 & Pic7z6[23]));
assign Fzo6x6 = (H0p6x6 & O0p6x6);
assign O0p6x6 = (~(vis_msp_o[23] & P42ov6));
assign H0p6x6 = (~(vis_r12_o[23] & W42ov6));
assign Ryo6x6 = (V0p6x6 & C1p6x6);
assign C1p6x6 = (J1p6x6 & Q1p6x6);
assign Q1p6x6 = (~(vis_r11_o[23] & F62ov6));
assign J1p6x6 = (~(vis_r10_o[23] & M62ov6));
assign V0p6x6 = (X1p6x6 & E2p6x6);
assign E2p6x6 = (~(vis_r9_o[23] & H72ov6));
assign X1p6x6 = (~(vis_r8_o[23] & O72ov6));
assign Dyo6x6 = (L2p6x6 & S2p6x6);
assign S2p6x6 = (Z2p6x6 & G3p6x6);
assign G3p6x6 = (N3p6x6 & U3p6x6);
assign U3p6x6 = (~(vis_r7_o[23] & L92ov6));
assign N3p6x6 = (~(vis_r6_o[23] & S92ov6));
assign Z2p6x6 = (B4p6x6 & I4p6x6);
assign I4p6x6 = (~(vis_r5_o[23] & Na2ov6));
assign B4p6x6 = (~(vis_r4_o[23] & Ua2ov6));
assign L2p6x6 = (P4p6x6 & W4p6x6);
assign W4p6x6 = (D5p6x6 & K5p6x6);
assign K5p6x6 = (~(vis_r3_o[23] & Dc2ov6));
assign D5p6x6 = (~(vis_r2_o[23] & Kc2ov6));
assign P4p6x6 = (R5p6x6 & Y5p6x6);
assign Y5p6x6 = (~(vis_r1_o[23] & Fd2ov6));
assign R5p6x6 = (~(vis_r0_o[23] & Md2ov6));
assign Pxo6x6 = (~(Td2ov6 & F8yiw6));
assign F8yiw6 = (Spyiw6 ? Ey97z6 : Gli7z6[23]);
assign Ey97z6 = (~(F6p6x6 & M6p6x6));
assign M6p6x6 = (~(Nqyiw6 & N7ynv6));
assign F6p6x6 = (T6p6x6 & A7p6x6);
assign A7p6x6 = (~(Pdc7z6[23] & Ouyiw6));
assign T6p6x6 = (~(Vuyiw6 & H7p6x6));
assign H7p6x6 = (~(O7p6x6 & V7p6x6));
assign V7p6x6 = (C8p6x6 & J8p6x6);
assign J8p6x6 = (Q8p6x6 & X8p6x6);
assign X8p6x6 = (E9p6x6 & L9p6x6);
assign L9p6x6 = (~(S9p6x6 & Uxyiw6));
assign S9p6x6 = (Kxb7z6[23] & Z9p6x6);
assign E9p6x6 = (~(Gap6x6 & Nap6x6));
assign Gap6x6 = (~(Uap6x6 & Quziw6));
assign Uap6x6 = (Bbp6x6 & Ibp6x6);
assign Ibp6x6 = (Z9p6x6 | Ninnv6);
assign Z9p6x6 = (Pbp6x6 | Rje7z6[23]);
assign Bbp6x6 = (~(Ofnnv6 & Pbp6x6));
assign Q8p6x6 = (Wbp6x6 & Dcp6x6);
assign Dcp6x6 = (~(T0ziw6 & Rje7z6[23]));
assign Wbp6x6 = (Ryfov6 | Kcp6x6);
assign C8p6x6 = (Rcp6x6 & Ycp6x6);
assign Ycp6x6 = (~(Cqf7z6[7] & Q2ziw6));
assign Rcp6x6 = (Fdp6x6 & Mdp6x6);
assign Mdp6x6 = (~(J73ov6 & Ok3ov6));
assign Fdp6x6 = (~(L0g7z6[23] & J2ziw6));
assign O7p6x6 = (Tdp6x6 & Aep6x6);
assign Aep6x6 = (Hep6x6 & Oep6x6);
assign Oep6x6 = (~(Z3ziw6 & Fhc7z6[8]));
assign Hep6x6 = (Vep6x6 & Cfp6x6);
assign Cfp6x6 = (~(L0g7z6[7] & O1ziw6));
assign Vep6x6 = (~(U4ziw6 & V1c7z6[23]));
assign Tdp6x6 = (Jfp6x6 & Dp3ov6);
assign Dp3ov6 = (Qfp6x6 & T7ziw6);
assign Qfp6x6 = (Xfp6x6 & Egp6x6);
assign Egp6x6 = (~(F7ziw6 & Y6ziw6));
assign Y6ziw6 = (~(Lgp6x6 ^ Nu8jw6));
assign Xfp6x6 = (~(R6ziw6 & M7ziw6));
assign M7ziw6 = (Kdziw6 ^ Dte7z6[1]);
assign Kdziw6 = (Kvbov6 ? Wx1ov6 : V1c7z6[31]);
assign Wx1ov6 = (Dte7z6[12] ? S7gdt6 : V5bov6);
assign Jfp6x6 = (U23ov6 & Sgp6x6);
assign Sgp6x6 = (~(Kaldt6 & Oztiw6));
assign U23ov6 = (Zgp6x6 & Ghp6x6);
assign Ghp6x6 = (~(Nhp6x6 & J2nnv6));
assign Nhp6x6 = (~(Q2nnv6 | Icziw6));
assign Zgp6x6 = (~(Uhp6x6 & Ubziw6));
assign Uhp6x6 = (~(J2nnv6 ^ Q2nnv6));
assign Q2nnv6 = (Bip6x6 ^ Mennv6);
assign Bip6x6 = (~(Iip6x6 & Pip6x6));
assign Pip6x6 = (Wip6x6 & Djp6x6);
assign Djp6x6 = (Kjp6x6 & Rjp6x6);
assign Rjp6x6 = (~(Yxf7z6[25] & Su0jw6));
assign Kjp6x6 = (Yjp6x6 & Fkp6x6);
assign Fkp6x6 = (~(Yxf7z6[23] & Nv0jw6));
assign Yjp6x6 = (~(Yxf7z6[24] & Uv0jw6));
assign Wip6x6 = (Mkp6x6 & Tkp6x6);
assign Tkp6x6 = (~(Yxf7z6[26] & Pw0jw6));
assign Mkp6x6 = (~(Lgp6x6 & Rdziw6));
assign Lgp6x6 = (T3cdt6 ? V1c7z6[23] : Nap6x6);
assign Iip6x6 = (Alp6x6 & Hlp6x6);
assign Hlp6x6 = (Olp6x6 & Vlp6x6);
assign Vlp6x6 = (~(Onf7z6[23] & My0jw6));
assign Olp6x6 = (Cmp6x6 & Jmp6x6);
assign Jmp6x6 = (~(Hz0jw6 & Kxb7z6[23]));
assign Cmp6x6 = (~(Oz0jw6 & Fhc7z6[23]));
assign Alp6x6 = (Qmp6x6 & Xmp6x6);
assign Xmp6x6 = (~(Alf7z6[7] & J01jw6));
assign Qmp6x6 = (~(Alf7z6[23] & Q01jw6));
assign J2nnv6 = (~(Enp6x6 ^ Tennv6));
assign Enp6x6 = (~(Lnp6x6 & Snp6x6));
assign Snp6x6 = (~(Yxf7z6[7] & Laziw6));
assign Lnp6x6 = (Znp6x6 & Gop6x6);
assign Gop6x6 = (~(Yxf7z6[23] & Gbziw6));
assign Znp6x6 = (~(Kxb7z6[23] & Nbziw6));
assign Nwo6x6 = (Nop6x6 & Uop6x6);
assign Uop6x6 = (~(Ve2ov6 & vis_pc_o[23]));
assign Nop6x6 = (~(Fhc7z6[23] & Cf2ov6));
assign Zvy7v6 = (~(Bpp6x6 & Ipp6x6));
assign Ipp6x6 = (Ppp6x6 & Wpp6x6);
assign Wpp6x6 = (Eu9ov6 | Dqp6x6);
assign Ppp6x6 = (Kqp6x6 & Rqp6x6);
assign Rqp6x6 = (~(Gv9ov6 & A9yiw6));
assign Kqp6x6 = (~(Uv9ov6 & Cz97z6));
assign Bpp6x6 = (Yqp6x6 & Frp6x6);
assign Frp6x6 = (~(Pw9ov6 & Kxb7z6[20]));
assign Yqp6x6 = (Mrp6x6 & Trp6x6);
assign Trp6x6 = (~(Kx9ov6 & vis_pc_o[20]));
assign Mrp6x6 = (~(Gli7z6[20] & Rx9ov6));
assign Svy7v6 = (~(Asp6x6 & Hsp6x6));
assign Hsp6x6 = (Osp6x6 & Vsp6x6);
assign Vsp6x6 = (~(Td2ov6 & A9yiw6));
assign A9yiw6 = (Spyiw6 ? Cz97z6 : Gli7z6[20]);
assign Td2ov6 = (~(Ctp6x6 | Jtp6x6));
assign Ctp6x6 = (Cf2ov6 | Mbihw6);
assign Osp6x6 = (Qtp6x6 & Xtp6x6);
assign Xtp6x6 = (~(H02ov6 & Cz97z6));
assign Cz97z6 = (~(Eup6x6 & Lup6x6));
assign Lup6x6 = (~(Nqyiw6 & Glynv6));
assign Eup6x6 = (Sup6x6 & Zup6x6);
assign Zup6x6 = (~(Pdc7z6[20] & Ouyiw6));
assign Sup6x6 = (~(Vuyiw6 & Gvp6x6));
assign Gvp6x6 = (~(Nvp6x6 & Uvp6x6));
assign Uvp6x6 = (Bwp6x6 & Iwp6x6);
assign Iwp6x6 = (Pwp6x6 & Wwp6x6);
assign Wwp6x6 = (Dxp6x6 & Kxp6x6);
assign Kxp6x6 = (~(Rxp6x6 & Uxyiw6));
assign Rxp6x6 = (Kxb7z6[20] & Yxp6x6);
assign Dxp6x6 = (~(Fyp6x6 & Myp6x6));
assign Fyp6x6 = (~(Typ6x6 & Quziw6));
assign Typ6x6 = (Azp6x6 & Hzp6x6);
assign Hzp6x6 = (Yxp6x6 | Ninnv6);
assign Yxp6x6 = (Ozp6x6 | Rje7z6[20]);
assign Azp6x6 = (~(Ofnnv6 & Ozp6x6));
assign Pwp6x6 = (Vzp6x6 & C0q6x6);
assign C0q6x6 = (~(J73ov6 & Ki3ov6));
assign Ki3ov6 = (~(Pch6x6 ^ Dte7z6[1]));
assign Pch6x6 = (T3cdt6 ? J0q6x6 : N14ov6);
assign Vzp6x6 = (~(F7ziw6 & Od3ov6));
assign Bwp6x6 = (Q0q6x6 & X0q6x6);
assign X0q6x6 = (E1q6x6 & L1q6x6);
assign L1q6x6 = (~(R6ziw6 & Xe3ov6));
assign E1q6x6 = (~(T0ziw6 & Rje7z6[20]));
assign Q0q6x6 = (S1q6x6 & Z1q6x6);
assign Z1q6x6 = (Ryfov6 | G2q6x6);
assign S1q6x6 = (~(L0g7z6[20] & J2ziw6));
assign Nvp6x6 = (N2q6x6 & U2q6x6);
assign U2q6x6 = (B3q6x6 & I3q6x6);
assign I3q6x6 = (P3q6x6 & W3q6x6);
assign W3q6x6 = (~(Cqf7z6[4] & Q2ziw6));
assign P3q6x6 = (~(L0g7z6[4] & O1ziw6));
assign B3q6x6 = (D4q6x6 & K4q6x6);
assign K4q6x6 = (~(U4ziw6 & V1c7z6[20]));
assign D4q6x6 = (~(Z3ziw6 & Fhc7z6[11]));
assign N2q6x6 = (R4q6x6 & N23ov6);
assign N23ov6 = (Y4q6x6 & F5q6x6);
assign F5q6x6 = (~(M5q6x6 & Z3nnv6));
assign M5q6x6 = (~(G4nnv6 | Icziw6));
assign Y4q6x6 = (~(T5q6x6 & Ubziw6));
assign T5q6x6 = (~(Z3nnv6 ^ G4nnv6));
assign G4nnv6 = (A6q6x6 ^ Mennv6);
assign A6q6x6 = (~(H6q6x6 & O6q6x6));
assign O6q6x6 = (V6q6x6 & C7q6x6);
assign C7q6x6 = (J7q6x6 & Q7q6x6);
assign Q7q6x6 = (~(Yxf7z6[22] & Su0jw6));
assign J7q6x6 = (X7q6x6 & E8q6x6);
assign E8q6x6 = (~(Yxf7z6[20] & Nv0jw6));
assign X7q6x6 = (~(Yxf7z6[21] & Uv0jw6));
assign V6q6x6 = (L8q6x6 & S8q6x6);
assign S8q6x6 = (~(Yxf7z6[23] & Pw0jw6));
assign L8q6x6 = (~(Z8q6x6 & Rdziw6));
assign H6q6x6 = (G9q6x6 & N9q6x6);
assign N9q6x6 = (U9q6x6 & Baq6x6);
assign Baq6x6 = (~(Onf7z6[20] & My0jw6));
assign U9q6x6 = (Iaq6x6 & Paq6x6);
assign Paq6x6 = (~(Hz0jw6 & Kxb7z6[20]));
assign Iaq6x6 = (~(Oz0jw6 & Fhc7z6[20]));
assign G9q6x6 = (Waq6x6 & Dbq6x6);
assign Dbq6x6 = (~(Alf7z6[4] & J01jw6));
assign Waq6x6 = (~(Alf7z6[20] & Q01jw6));
assign Z3nnv6 = (~(Kbq6x6 ^ Tennv6));
assign Kbq6x6 = (~(Rbq6x6 & Ybq6x6));
assign Ybq6x6 = (~(Yxf7z6[4] & Laziw6));
assign Rbq6x6 = (Fcq6x6 & Mcq6x6);
assign Mcq6x6 = (~(Yxf7z6[20] & Gbziw6));
assign Fcq6x6 = (~(Kxb7z6[20] & Nbziw6));
assign R4q6x6 = (T7ziw6 & Tcq6x6);
assign Tcq6x6 = (~(Tgldt6 & Oztiw6));
assign H02ov6 = (Adq6x6 & C3yiw6);
assign Adq6x6 = (Hdq6x6 & Mbihw6);
assign Qtp6x6 = (C12ov6 | M3knv6);
assign M3knv6 = (Odq6x6 & Vdq6x6);
assign Vdq6x6 = (Ceq6x6 & Jeq6x6);
assign Jeq6x6 = (Qeq6x6 & Xeq6x6);
assign Xeq6x6 = (Efq6x6 & Lfq6x6);
assign Lfq6x6 = (~(vis_psp_o[20] & N32ov6));
assign N32ov6 = (~(Y3ihw6 | Sfq6x6));
assign Efq6x6 = (~(U32ov6 & Pic7z6[20]));
assign U32ov6 = (Yzriw6 & Zfq6x6);
assign Qeq6x6 = (Ggq6x6 & Ngq6x6);
assign Ngq6x6 = (~(vis_msp_o[20] & P42ov6));
assign P42ov6 = (~(Zfq6x6 | Y3ihw6));
assign Ggq6x6 = (~(vis_r12_o[20] & W42ov6));
assign W42ov6 = (Sfq6x6 & Yzriw6);
assign Ceq6x6 = (Ugq6x6 & Bhq6x6);
assign Bhq6x6 = (Ihq6x6 & Phq6x6);
assign Phq6x6 = (~(vis_r11_o[20] & F62ov6));
assign F62ov6 = (Whq6x6 & Diq6x6);
assign Ihq6x6 = (~(vis_r10_o[20] & M62ov6));
assign M62ov6 = (Kiq6x6 & Diq6x6);
assign Ugq6x6 = (Riq6x6 & Yiq6x6);
assign Yiq6x6 = (~(vis_r9_o[20] & H72ov6));
assign H72ov6 = (Whq6x6 & Fjq6x6);
assign Whq6x6 = (Nfihw6 & Zeihw6);
assign Riq6x6 = (~(vis_r8_o[20] & O72ov6));
assign O72ov6 = (Kiq6x6 & Fjq6x6);
assign Kiq6x6 = (Mjq6x6 & Nfihw6);
assign Odq6x6 = (Tjq6x6 & Akq6x6);
assign Akq6x6 = (Hkq6x6 & Okq6x6);
assign Okq6x6 = (Vkq6x6 & Clq6x6);
assign Clq6x6 = (~(vis_r7_o[20] & L92ov6));
assign L92ov6 = (Jlq6x6 & Qlq6x6);
assign Vkq6x6 = (~(vis_r6_o[20] & S92ov6));
assign S92ov6 = (Jlq6x6 & Xlq6x6);
assign Jlq6x6 = (Zfq6x6 & Xdihw6);
assign Hkq6x6 = (Emq6x6 & Lmq6x6);
assign Lmq6x6 = (~(vis_r5_o[20] & Na2ov6));
assign Na2ov6 = (Smq6x6 & Qlq6x6);
assign Emq6x6 = (~(vis_r4_o[20] & Ua2ov6));
assign Ua2ov6 = (Smq6x6 & Xlq6x6);
assign Smq6x6 = (Sfq6x6 & Xdihw6);
assign Tjq6x6 = (Zmq6x6 & Gnq6x6);
assign Gnq6x6 = (Nnq6x6 & Unq6x6);
assign Unq6x6 = (~(vis_r3_o[20] & Dc2ov6));
assign Dc2ov6 = (Qlq6x6 & Diq6x6);
assign Nnq6x6 = (~(vis_r2_o[20] & Kc2ov6));
assign Kc2ov6 = (Xlq6x6 & Diq6x6);
assign Diq6x6 = (~(Xdihw6 | Sfq6x6));
assign Zmq6x6 = (Boq6x6 & Ioq6x6);
assign Ioq6x6 = (~(vis_r1_o[20] & Fd2ov6));
assign Fd2ov6 = (Qlq6x6 & Fjq6x6);
assign Qlq6x6 = (~(Nfihw6 | Mjq6x6));
assign Boq6x6 = (~(vis_r0_o[20] & Md2ov6));
assign Md2ov6 = (Xlq6x6 & Fjq6x6);
assign Fjq6x6 = (~(Zfq6x6 | Xdihw6));
assign Xlq6x6 = (~(Nfihw6 | Zeihw6));
assign C12ov6 = (!Ktxiw6);
assign Ktxiw6 = (Poq6x6 & Hdq6x6);
assign Poq6x6 = (Jtp6x6 & Bmknv6);
assign Bmknv6 = (!Mbihw6);
assign Jtp6x6 = (~(Woq6x6 & Dpq6x6));
assign Dpq6x6 = (Kpq6x6 & Rpq6x6);
assign Rpq6x6 = (Ylyiw6 ^ Sfq6x6);
assign Sfq6x6 = (!Zfq6x6);
assign Zfq6x6 = (~(Ypq6x6 & Fqq6x6));
assign Fqq6x6 = (~(Mqq6x6 & Tqq6x6));
assign Kpq6x6 = (Liyiw6 & Arq6x6);
assign Arq6x6 = (Zeihw6 ^ Bkyiw6);
assign Woq6x6 = (Hrq6x6 & Orq6x6);
assign Orq6x6 = (Mlziw6 ^ Nfihw6);
assign Hrq6x6 = (Coyiw6 ^ Xdihw6);
assign Asp6x6 = (Vrq6x6 & Csq6x6);
assign Csq6x6 = (~(Ve2ov6 & vis_pc_o[20]));
assign Ve2ov6 = (Jsq6x6 & Hdq6x6);
assign Hdq6x6 = (!Cf2ov6);
assign Jsq6x6 = (Mbihw6 & Qsq6x6);
assign Mbihw6 = (Mqq6x6 & F4ihw6);
assign Mqq6x6 = (!Y3ihw6);
assign Y3ihw6 = (~(Xsq6x6 & Nfihw6));
assign Xsq6x6 = (Xdihw6 & Zeihw6);
assign Vrq6x6 = (~(Fhc7z6[20] & Cf2ov6));
assign Cf2ov6 = (~(Etq6x6 & Ltq6x6));
assign Lvy7v6 = (Z6jhw6 ? D5f7z6[3] : Wjnnv6);
assign Wjnnv6 = (Ua0jw6 | P40jw6);
assign Evy7v6 = (~(Stq6x6 & Ztq6x6));
assign Ztq6x6 = (Guq6x6 & Nuq6x6);
assign Nuq6x6 = (~(Myp6x6 & C6bov6));
assign Guq6x6 = (~(J6bov6 & Alf7z6[20]));
assign Stq6x6 = (Uuq6x6 & Bvq6x6);
assign Bvq6x6 = (~(Cqf7z6[4] & E7bov6));
assign Uuq6x6 = (~(L0g7z6[20] & L7bov6));
assign Xuy7v6 = (~(Ivq6x6 & Pvq6x6));
assign Pvq6x6 = (Wvq6x6 & Dwq6x6);
assign Dwq6x6 = (~(Lt3ov6 & C6bov6));
assign Wvq6x6 = (~(J6bov6 & Alf7z6[29]));
assign Ivq6x6 = (Kwq6x6 & Rwq6x6);
assign Rwq6x6 = (~(Cqf7z6[13] & E7bov6));
assign Kwq6x6 = (~(L0g7z6[29] & L7bov6));
assign Quy7v6 = (~(Ywq6x6 & Fxq6x6));
assign Fxq6x6 = (Mxq6x6 & Txq6x6);
assign Txq6x6 = (~(Uu3ov6 & C6bov6));
assign Mxq6x6 = (~(J6bov6 & Alf7z6[28]));
assign Ywq6x6 = (Ayq6x6 & Hyq6x6);
assign Hyq6x6 = (~(Cqf7z6[12] & E7bov6));
assign Ayq6x6 = (~(L0g7z6[28] & L7bov6));
assign Juy7v6 = (~(Oyq6x6 & Vyq6x6));
assign Vyq6x6 = (Czq6x6 & Jzq6x6);
assign Jzq6x6 = (~(M85jw6 & C6bov6));
assign Czq6x6 = (~(J6bov6 & Alf7z6[15]));
assign Oyq6x6 = (Qzq6x6 & Xzq6x6);
assign Xzq6x6 = (~(L0g7z6[31] & E7bov6));
assign Qzq6x6 = (~(L0g7z6[15] & L7bov6));
assign Cuy7v6 = (~(E0r6x6 & L0r6x6));
assign L0r6x6 = (S0r6x6 & Z0r6x6);
assign Z0r6x6 = (~(Nap6x6 & C6bov6));
assign S0r6x6 = (~(J6bov6 & Alf7z6[23]));
assign E0r6x6 = (G1r6x6 & N1r6x6);
assign N1r6x6 = (~(Cqf7z6[7] & E7bov6));
assign G1r6x6 = (~(L0g7z6[23] & L7bov6));
assign Vty7v6 = (~(U1r6x6 & B2r6x6));
assign B2r6x6 = (I2r6x6 & P2r6x6);
assign P2r6x6 = (~(Bv3ov6 & C6bov6));
assign I2r6x6 = (~(J6bov6 & Alf7z6[7]));
assign U1r6x6 = (W2r6x6 & D3r6x6);
assign D3r6x6 = (~(L0g7z6[23] & E7bov6));
assign W2r6x6 = (~(L0g7z6[7] & L7bov6));
assign Oty7v6 = (~(K3r6x6 & R3r6x6));
assign R3r6x6 = (Y3r6x6 & F4r6x6);
assign F4r6x6 = (~(Zbn6x6 & C6bov6));
assign Y3r6x6 = (~(J6bov6 & Alf7z6[14]));
assign K3r6x6 = (M4r6x6 & T4r6x6);
assign T4r6x6 = (~(L0g7z6[30] & E7bov6));
assign M4r6x6 = (~(L0g7z6[14] & L7bov6));
assign Hty7v6 = (~(A5r6x6 & H5r6x6));
assign H5r6x6 = (O5r6x6 & V5r6x6);
assign V5r6x6 = (~(Yfm6x6 & C6bov6));
assign O5r6x6 = (~(J6bov6 & Alf7z6[22]));
assign A5r6x6 = (C6r6x6 & J6r6x6);
assign J6r6x6 = (~(Cqf7z6[6] & E7bov6));
assign C6r6x6 = (~(L0g7z6[22] & L7bov6));
assign Aty7v6 = (~(Q6r6x6 & X6r6x6));
assign X6r6x6 = (E7r6x6 & L7r6x6);
assign L7r6x6 = (~(Nu3ov6 & C6bov6));
assign E7r6x6 = (~(J6bov6 & Alf7z6[6]));
assign Q6r6x6 = (S7r6x6 & Z7r6x6);
assign Z7r6x6 = (~(L0g7z6[22] & E7bov6));
assign S7r6x6 = (~(L0g7z6[6] & L7bov6));
assign Tsy7v6 = (~(G8r6x6 & N8r6x6));
assign N8r6x6 = (U8r6x6 & B9r6x6);
assign B9r6x6 = (~(Dok6x6 & C6bov6));
assign U8r6x6 = (~(J6bov6 & Alf7z6[13]));
assign G8r6x6 = (I9r6x6 & P9r6x6);
assign P9r6x6 = (~(L0g7z6[29] & E7bov6));
assign I9r6x6 = (~(L0g7z6[13] & L7bov6));
assign Msy7v6 = (~(W9r6x6 & Dar6x6));
assign Dar6x6 = (Kar6x6 & Rar6x6);
assign Rar6x6 = (~(Csj6x6 & C6bov6));
assign Kar6x6 = (~(J6bov6 & Alf7z6[21]));
assign W9r6x6 = (Yar6x6 & Fbr6x6);
assign Fbr6x6 = (~(Cqf7z6[5] & E7bov6));
assign Yar6x6 = (~(L0g7z6[21] & L7bov6));
assign Fsy7v6 = (~(Mbr6x6 & Tbr6x6));
assign Tbr6x6 = (Acr6x6 & Hcr6x6);
assign Hcr6x6 = (~(Xs3ov6 & C6bov6));
assign Acr6x6 = (~(J6bov6 & Alf7z6[5]));
assign Mbr6x6 = (Ocr6x6 & Vcr6x6);
assign Vcr6x6 = (~(L0g7z6[21] & E7bov6));
assign Ocr6x6 = (~(L0g7z6[5] & L7bov6));
assign Yry7v6 = (~(Cdr6x6 & Jdr6x6));
assign Jdr6x6 = (Qdr6x6 & Xdr6x6);
assign Xdr6x6 = (~(Et3ov6 & C6bov6));
assign Qdr6x6 = (~(J6bov6 & Alf7z6[4]));
assign Cdr6x6 = (Eer6x6 & Ler6x6);
assign Ler6x6 = (~(L0g7z6[20] & E7bov6));
assign Eer6x6 = (~(L0g7z6[4] & L7bov6));
assign Rry7v6 = (~(Ser6x6 & Zer6x6));
assign Zer6x6 = (Gfr6x6 & Nfr6x6);
assign Nfr6x6 = (~(Ryh6x6 & C6bov6));
assign Gfr6x6 = (~(J6bov6 & Alf7z6[3]));
assign Ser6x6 = (Ufr6x6 & Bgr6x6);
assign Bgr6x6 = (~(L0g7z6[19] & E7bov6));
assign Ufr6x6 = (~(L0g7z6[3] & L7bov6));
assign Kry7v6 = (~(Igr6x6 & Pgr6x6));
assign Pgr6x6 = (Wgr6x6 & Dhr6x6);
assign Dhr6x6 = (~(X2h6x6 & C6bov6));
assign Wgr6x6 = (~(J6bov6 & Alf7z6[12]));
assign Igr6x6 = (Khr6x6 & Rhr6x6);
assign Rhr6x6 = (~(L0g7z6[28] & E7bov6));
assign Khr6x6 = (~(L0g7z6[12] & L7bov6));
assign Dry7v6 = (~(Yhr6x6 & Fir6x6));
assign Fir6x6 = (Mir6x6 & Tir6x6);
assign Tir6x6 = (~(O9cjw6 & C6bov6));
assign Mir6x6 = (~(J6bov6 & Alf7z6[19]));
assign Yhr6x6 = (Ajr6x6 & Hjr6x6);
assign Hjr6x6 = (~(Cqf7z6[3] & E7bov6));
assign Ajr6x6 = (~(L0g7z6[19] & L7bov6));
assign Wqy7v6 = (~(Ojr6x6 & Vjr6x6));
assign Vjr6x6 = (Ckr6x6 & Jkr6x6);
assign Jkr6x6 = (~(Pebjw6 & C6bov6));
assign Ckr6x6 = (~(J6bov6 & Alf7z6[11]));
assign Ojr6x6 = (Qkr6x6 & Xkr6x6);
assign Xkr6x6 = (~(L0g7z6[27] & E7bov6));
assign Qkr6x6 = (~(L0g7z6[11] & L7bov6));
assign Pqy7v6 = (~(Elr6x6 & Llr6x6));
assign Llr6x6 = (Slr6x6 & Zlr6x6);
assign Zlr6x6 = (~(Oiajw6 & C6bov6));
assign Slr6x6 = (~(J6bov6 & Alf7z6[17]));
assign Elr6x6 = (Gmr6x6 & Nmr6x6);
assign Nmr6x6 = (~(Cqf7z6[1] & E7bov6));
assign Gmr6x6 = (~(L0g7z6[17] & L7bov6));
assign Iqy7v6 = (~(Umr6x6 & Bnr6x6));
assign Bnr6x6 = (Inr6x6 & Pnr6x6);
assign Pnr6x6 = (~(Pn9jw6 & C6bov6));
assign Inr6x6 = (~(J6bov6 & Alf7z6[9]));
assign Umr6x6 = (Wnr6x6 & Dor6x6);
assign Dor6x6 = (~(L0g7z6[25] & E7bov6));
assign Wnr6x6 = (~(L0g7z6[9] & L7bov6));
assign Bqy7v6 = (~(Kor6x6 & Ror6x6));
assign Ror6x6 = (Yor6x6 & Fpr6x6);
assign Fpr6x6 = (~(Ku3jw6 & C6bov6));
assign Yor6x6 = (~(J6bov6 & Alf7z6[8]));
assign Kor6x6 = (Mpr6x6 & Tpr6x6);
assign Tpr6x6 = (~(L0g7z6[24] & E7bov6));
assign Mpr6x6 = (~(L0g7z6[8] & L7bov6));
assign Upy7v6 = (~(Aqr6x6 & Hqr6x6));
assign Hqr6x6 = (Oqr6x6 & Vqr6x6);
assign Vqr6x6 = (~(Hr8jw6 & C6bov6));
assign Oqr6x6 = (~(J6bov6 & Alf7z6[16]));
assign Aqr6x6 = (Crr6x6 & Jrr6x6);
assign Jrr6x6 = (~(Cqf7z6[0] & E7bov6));
assign Crr6x6 = (~(L0g7z6[16] & L7bov6));
assign Npy7v6 = (~(Qrr6x6 & Xrr6x6));
assign Xrr6x6 = (Esr6x6 & Lsr6x6);
assign Lsr6x6 = (~(A07jw6 & C6bov6));
assign Esr6x6 = (~(J6bov6 & Alf7z6[25]));
assign Qrr6x6 = (Ssr6x6 & Zsr6x6);
assign Zsr6x6 = (~(Cqf7z6[9] & E7bov6));
assign Ssr6x6 = (~(L0g7z6[25] & L7bov6));
assign Gpy7v6 = (~(Gtr6x6 & Ntr6x6));
assign Ntr6x6 = (~(Eji7z6[26] & C3yiw6));
assign Gtr6x6 = (Utr6x6 & Bur6x6);
assign Bur6x6 = (~(Bhi7z6[26] & X3yiw6));
assign Utr6x6 = (~(E4yiw6 & vis_pc_o[26]));
assign Zoy7v6 = (~(Iur6x6 & Pur6x6));
assign Pur6x6 = (~(Eji7z6[27] & C3yiw6));
assign Iur6x6 = (Wur6x6 & Dvr6x6);
assign Dvr6x6 = (~(Bhi7z6[27] & X3yiw6));
assign Wur6x6 = (~(E4yiw6 & vis_pc_o[27]));
assign Soy7v6 = (~(Kvr6x6 & Rvr6x6));
assign Rvr6x6 = (~(Eji7z6[28] & C3yiw6));
assign Kvr6x6 = (Yvr6x6 & Fwr6x6);
assign Fwr6x6 = (~(Bhi7z6[28] & X3yiw6));
assign Yvr6x6 = (~(E4yiw6 & vis_pc_o[28]));
assign Loy7v6 = (~(Mwr6x6 & Twr6x6));
assign Twr6x6 = (~(Eji7z6[29] & C3yiw6));
assign Mwr6x6 = (Axr6x6 & Hxr6x6);
assign Hxr6x6 = (~(Bhi7z6[29] & X3yiw6));
assign Axr6x6 = (~(E4yiw6 & vis_pc_o[29]));
assign Eoy7v6 = (~(Oxr6x6 & Vxr6x6));
assign Vxr6x6 = (~(Eji7z6[30] & C3yiw6));
assign Oxr6x6 = (Cyr6x6 & Jyr6x6);
assign Jyr6x6 = (~(Bhi7z6[30] & X3yiw6));
assign Cyr6x6 = (~(E4yiw6 & vis_pc_o[30]));
assign Xny7v6 = (~(Qyr6x6 & Xyr6x6));
assign Xyr6x6 = (~(Eji7z6[31] & C3yiw6));
assign Qyr6x6 = (Ezr6x6 & Lzr6x6);
assign Lzr6x6 = (~(Bhi7z6[31] & X3yiw6));
assign X3yiw6 = (~(E4yiw6 | C3yiw6));
assign Ezr6x6 = (~(E4yiw6 & vis_pc_o[31]));
assign E4yiw6 = (~(Ut2jw6 | C3yiw6));
assign Qny7v6 = (~(Szr6x6 & Zzr6x6));
assign Zzr6x6 = (G0s6x6 & N0s6x6);
assign N0s6x6 = (Eu9ov6 | U0s6x6);
assign G0s6x6 = (B1s6x6 & I1s6x6);
assign I1s6x6 = (~(Gv9ov6 & W7xiw6));
assign W7xiw6 = (Gninv6 ? Gli7z6[26] : Qw97z6);
assign B1s6x6 = (~(Uv9ov6 & Qw97z6));
assign Qw97z6 = (~(P1s6x6 & W1s6x6));
assign W1s6x6 = (~(Nqyiw6 & Iuxnv6));
assign P1s6x6 = (D2s6x6 & K2s6x6);
assign K2s6x6 = (~(Pdc7z6[26] & Ouyiw6));
assign D2s6x6 = (~(Vuyiw6 & R2s6x6));
assign R2s6x6 = (~(Y2s6x6 & F3s6x6));
assign F3s6x6 = (M3s6x6 & T3s6x6);
assign T3s6x6 = (A4s6x6 & H4s6x6);
assign H4s6x6 = (O4s6x6 & V4s6x6);
assign V4s6x6 = (~(C5s6x6 & Uxyiw6));
assign C5s6x6 = (Kxb7z6[26] & J5s6x6);
assign O4s6x6 = (~(Qs3ov6 & Q5s6x6));
assign Q5s6x6 = (~(X5s6x6 & Quziw6));
assign X5s6x6 = (E6s6x6 & L6s6x6);
assign L6s6x6 = (J5s6x6 | Ninnv6);
assign J5s6x6 = (S6s6x6 | Rje7z6[26]);
assign E6s6x6 = (~(Ofnnv6 & S6s6x6));
assign A4s6x6 = (Z6s6x6 & G7s6x6);
assign G7s6x6 = (~(J73ov6 & Un3ov6));
assign Un3ov6 = (~(M42jw6 ^ Dte7z6[1]));
assign M42jw6 = (T3cdt6 ? N7s6x6 : Fx3ov6);
assign Z6s6x6 = (~(F7ziw6 & Db3ov6));
assign Db3ov6 = (U7s6x6 ^ Dte7z6[1]);
assign M3s6x6 = (B8s6x6 & I8s6x6);
assign I8s6x6 = (P8s6x6 & W8s6x6);
assign W8s6x6 = (~(R6ziw6 & Vd3ov6));
assign Vd3ov6 = (K66jw6 ^ Dte7z6[1]);
assign K66jw6 = (T3cdt6 ? V1c7z6[18] : Ew5jw6);
assign P8s6x6 = (~(T0ziw6 & Rje7z6[26]));
assign B8s6x6 = (D9s6x6 & K9s6x6);
assign K9s6x6 = (Ryfov6 | R9s6x6);
assign R9s6x6 = (!S6s6x6);
assign D9s6x6 = (~(L0g7z6[26] & J2ziw6));
assign Y2s6x6 = (Y9s6x6 & Fas6x6);
assign Fas6x6 = (Mas6x6 & Tas6x6);
assign Tas6x6 = (Abs6x6 & Hbs6x6);
assign Hbs6x6 = (~(Cqf7z6[10] & Q2ziw6));
assign Abs6x6 = (~(L0g7z6[10] & O1ziw6));
assign Mas6x6 = (Obs6x6 & Vbs6x6);
assign Vbs6x6 = (~(U4ziw6 & V1c7z6[26]));
assign Obs6x6 = (~(Z3ziw6 & Fhc7z6[5]));
assign Y9s6x6 = (Ccs6x6 & W33ov6);
assign W33ov6 = (Jcs6x6 & Qcs6x6);
assign Qcs6x6 = (~(Xcs6x6 & T0nnv6));
assign Xcs6x6 = (~(A1nnv6 | Icziw6));
assign Jcs6x6 = (~(Eds6x6 & Ubziw6));
assign Eds6x6 = (~(T0nnv6 ^ A1nnv6));
assign A1nnv6 = (Lds6x6 ^ Mennv6);
assign Lds6x6 = (~(Sds6x6 & Zds6x6));
assign Zds6x6 = (Ges6x6 & Nes6x6);
assign Nes6x6 = (Ues6x6 & Bfs6x6);
assign Bfs6x6 = (~(Su0jw6 & Yxf7z6[28]));
assign Ues6x6 = (Ifs6x6 & Pfs6x6);
assign Pfs6x6 = (~(Yxf7z6[26] & Nv0jw6));
assign Ifs6x6 = (~(Yxf7z6[27] & Uv0jw6));
assign Ges6x6 = (Wfs6x6 & Dgs6x6);
assign Dgs6x6 = (~(Pw0jw6 & Yxf7z6[29]));
assign Wfs6x6 = (~(U7s6x6 & Rdziw6));
assign U7s6x6 = (T3cdt6 ? V1c7z6[26] : Qs3ov6);
assign Sds6x6 = (Kgs6x6 & Rgs6x6);
assign Rgs6x6 = (Ygs6x6 & Fhs6x6);
assign Fhs6x6 = (~(Onf7z6[26] & My0jw6));
assign Ygs6x6 = (Mhs6x6 & Ths6x6);
assign Ths6x6 = (~(Hz0jw6 & Kxb7z6[26]));
assign Mhs6x6 = (~(Oz0jw6 & Fhc7z6[26]));
assign Kgs6x6 = (Ais6x6 & His6x6);
assign His6x6 = (~(Alf7z6[10] & J01jw6));
assign Ais6x6 = (~(Alf7z6[26] & Q01jw6));
assign T0nnv6 = (~(Ois6x6 ^ Tennv6));
assign Ois6x6 = (~(Vis6x6 & Cjs6x6));
assign Cjs6x6 = (~(Yxf7z6[10] & Laziw6));
assign Vis6x6 = (Jjs6x6 & Qjs6x6);
assign Qjs6x6 = (~(Yxf7z6[26] & Gbziw6));
assign Jjs6x6 = (~(Kxb7z6[26] & Nbziw6));
assign Ccs6x6 = (T7ziw6 & Xjs6x6);
assign Xjs6x6 = (~(B4ldt6 & Oztiw6));
assign Szr6x6 = (Eks6x6 & Lks6x6);
assign Lks6x6 = (~(Pw9ov6 & Kxb7z6[26]));
assign Eks6x6 = (Sks6x6 & Zks6x6);
assign Zks6x6 = (~(Kx9ov6 & vis_pc_o[26]));
assign Sks6x6 = (~(Gli7z6[26] & Rx9ov6));
assign Jny7v6 = (~(Gls6x6 & Nls6x6));
assign Nls6x6 = (Uls6x6 & Bms6x6);
assign Bms6x6 = (~(Kp1jw6 & C6bov6));
assign Uls6x6 = (~(J6bov6 & Alf7z6[2]));
assign Gls6x6 = (Ims6x6 & Pms6x6);
assign Pms6x6 = (~(L0g7z6[18] & E7bov6));
assign Ims6x6 = (~(L0g7z6[2] & L7bov6));
assign Cny7v6 = (~(Wms6x6 & Dns6x6));
assign Dns6x6 = (Kns6x6 & Rns6x6);
assign Rns6x6 = (~(Ci4jw6 & C6bov6));
assign Kns6x6 = (~(J6bov6 & Alf7z6[10]));
assign Wms6x6 = (Yns6x6 & Fos6x6);
assign Fos6x6 = (~(L0g7z6[26] & E7bov6));
assign Yns6x6 = (~(L0g7z6[10] & L7bov6));
assign Vmy7v6 = (~(Mos6x6 & Tos6x6));
assign Tos6x6 = (Aps6x6 & Hps6x6);
assign Hps6x6 = (~(Ew5jw6 & C6bov6));
assign Aps6x6 = (~(J6bov6 & Alf7z6[18]));
assign Mos6x6 = (Ops6x6 & Vps6x6);
assign Vps6x6 = (~(Cqf7z6[2] & E7bov6));
assign Ops6x6 = (~(L0g7z6[18] & L7bov6));
assign Omy7v6 = (~(Cqs6x6 & Jqs6x6));
assign Jqs6x6 = (Qqs6x6 & Xqs6x6);
assign Xqs6x6 = (Eu9ov6 | Ers6x6);
assign Qqs6x6 = (Lrs6x6 & Srs6x6);
assign Srs6x6 = (~(Gv9ov6 & S2gov6));
assign S2gov6 = (Gninv6 ? Gli7z6[27] : Sv97z6);
assign Lrs6x6 = (~(Uv9ov6 & Sv97z6));
assign Sv97z6 = (~(Zrs6x6 & Gss6x6));
assign Gss6x6 = (~(Nqyiw6 & Tpxnv6));
assign Zrs6x6 = (Nss6x6 & Uss6x6);
assign Uss6x6 = (~(Pdc7z6[27] & Ouyiw6));
assign Nss6x6 = (~(Vuyiw6 & Bts6x6));
assign Bts6x6 = (~(Its6x6 & Pts6x6));
assign Pts6x6 = (Wts6x6 & Dus6x6);
assign Dus6x6 = (Kus6x6 & Rus6x6);
assign Rus6x6 = (Yus6x6 & Fvs6x6);
assign Fvs6x6 = (~(Mvs6x6 & Uxyiw6));
assign Mvs6x6 = (Kxb7z6[27] & Tvs6x6);
assign Yus6x6 = (~(St3ov6 & Aws6x6));
assign Aws6x6 = (~(Hws6x6 & Quziw6));
assign Hws6x6 = (Ows6x6 & Vws6x6);
assign Vws6x6 = (Tvs6x6 | Ninnv6);
assign Tvs6x6 = (Cxs6x6 | Rje7z6[27]);
assign Ows6x6 = (~(Ofnnv6 & Cxs6x6));
assign Kus6x6 = (Jxs6x6 & Qxs6x6);
assign Qxs6x6 = (~(J73ov6 & Xl3ov6));
assign Xl3ov6 = (~(L9i6x6 ^ Dte7z6[1]));
assign L9i6x6 = (T3cdt6 ? G8phw6 : Ay3ov6);
assign Jxs6x6 = (~(R6ziw6 & Hd3ov6));
assign Hd3ov6 = (Ujcjw6 ^ Dte7z6[1]);
assign Ujcjw6 = (T3cdt6 ? V1c7z6[19] : O9cjw6);
assign Wts6x6 = (Xxs6x6 & Eys6x6);
assign Eys6x6 = (Lys6x6 & Sys6x6);
assign Sys6x6 = (~(F7ziw6 & Ad3ov6));
assign Ad3ov6 = (Zys6x6 ^ Dte7z6[1]);
assign Lys6x6 = (~(T0ziw6 & Rje7z6[27]));
assign Xxs6x6 = (Gzs6x6 & Nzs6x6);
assign Nzs6x6 = (Ryfov6 | Uzs6x6);
assign Uzs6x6 = (!Cxs6x6);
assign Gzs6x6 = (~(L0g7z6[27] & J2ziw6));
assign Its6x6 = (B0t6x6 & I0t6x6);
assign I0t6x6 = (P0t6x6 & W0t6x6);
assign W0t6x6 = (D1t6x6 & K1t6x6);
assign K1t6x6 = (~(Cqf7z6[11] & Q2ziw6));
assign D1t6x6 = (~(L0g7z6[11] & O1ziw6));
assign P0t6x6 = (R1t6x6 & Y1t6x6);
assign Y1t6x6 = (~(U4ziw6 & V1c7z6[27]));
assign R1t6x6 = (~(B5ziw6 & Lsfdt6));
assign B0t6x6 = (F2t6x6 & M2t6x6);
assign M2t6x6 = (T2t6x6 & A3t6x6);
assign A3t6x6 = (~(Z3ziw6 & E3c7z6[4]));
assign T2t6x6 = (~(Y1ldt6 & Oztiw6));
assign F2t6x6 = (P33ov6 & T7ziw6);
assign P33ov6 = (H3t6x6 & O3t6x6);
assign O3t6x6 = (~(V3t6x6 & F0nnv6));
assign V3t6x6 = (~(M0nnv6 | Icziw6));
assign H3t6x6 = (~(C4t6x6 & Ubziw6));
assign C4t6x6 = (~(F0nnv6 ^ M0nnv6));
assign M0nnv6 = (J4t6x6 ^ Mennv6);
assign J4t6x6 = (~(Q4t6x6 & X4t6x6));
assign X4t6x6 = (E5t6x6 & L5t6x6);
assign L5t6x6 = (S5t6x6 & Z5t6x6);
assign Z5t6x6 = (~(Su0jw6 & Yxf7z6[29]));
assign S5t6x6 = (G6t6x6 & N6t6x6);
assign N6t6x6 = (~(Yxf7z6[27] & Nv0jw6));
assign G6t6x6 = (~(Uv0jw6 & Yxf7z6[28]));
assign E5t6x6 = (U6t6x6 & B7t6x6);
assign B7t6x6 = (~(Pw0jw6 & Yxf7z6[30]));
assign U6t6x6 = (~(Zys6x6 & Rdziw6));
assign Zys6x6 = (T3cdt6 ? V1c7z6[27] : St3ov6);
assign Q4t6x6 = (I7t6x6 & P7t6x6);
assign P7t6x6 = (W7t6x6 & D8t6x6);
assign D8t6x6 = (~(Onf7z6[27] & My0jw6));
assign W7t6x6 = (K8t6x6 & R8t6x6);
assign R8t6x6 = (~(Hz0jw6 & Kxb7z6[27]));
assign K8t6x6 = (~(Oz0jw6 & Fhc7z6[27]));
assign I7t6x6 = (Y8t6x6 & F9t6x6);
assign F9t6x6 = (~(Alf7z6[11] & J01jw6));
assign Y8t6x6 = (~(Alf7z6[27] & Q01jw6));
assign F0nnv6 = (~(M9t6x6 ^ Tennv6));
assign M9t6x6 = (~(T9t6x6 & Aat6x6));
assign Aat6x6 = (~(Yxf7z6[11] & Laziw6));
assign T9t6x6 = (Hat6x6 & Oat6x6);
assign Oat6x6 = (~(Yxf7z6[27] & Gbziw6));
assign Hat6x6 = (~(Kxb7z6[27] & Nbziw6));
assign Cqs6x6 = (Vat6x6 & Cbt6x6);
assign Cbt6x6 = (~(Pw9ov6 & Kxb7z6[27]));
assign Vat6x6 = (Jbt6x6 & Qbt6x6);
assign Qbt6x6 = (~(Kx9ov6 & vis_pc_o[27]));
assign Jbt6x6 = (~(Gli7z6[27] & Rx9ov6));
assign Hmy7v6 = (~(Xbt6x6 & Ect6x6));
assign Ect6x6 = (Lct6x6 & Sct6x6);
assign Sct6x6 = (Eu9ov6 | Zct6x6);
assign Lct6x6 = (Gdt6x6 & Ndt6x6);
assign Ndt6x6 = (~(Gv9ov6 & C7aov6));
assign C7aov6 = (Gninv6 ? Gli7z6[28] : Uu97z6);
assign Gdt6x6 = (~(Uv9ov6 & Uu97z6));
assign Uu97z6 = (~(Udt6x6 & Bet6x6));
assign Bet6x6 = (~(Nqyiw6 & Elxnv6));
assign Udt6x6 = (Iet6x6 & Pet6x6);
assign Pet6x6 = (~(Pdc7z6[28] & Ouyiw6));
assign Iet6x6 = (~(Vuyiw6 & Wet6x6));
assign Wet6x6 = (~(Dft6x6 & Kft6x6));
assign Kft6x6 = (Rft6x6 & Yft6x6);
assign Yft6x6 = (Fgt6x6 & Mgt6x6);
assign Mgt6x6 = (Tgt6x6 & Aht6x6);
assign Aht6x6 = (~(Hht6x6 & Uxyiw6));
assign Hht6x6 = (Kxb7z6[28] & Oht6x6);
assign Tgt6x6 = (~(Uu3ov6 & Vht6x6));
assign Vht6x6 = (~(Cit6x6 & Quziw6));
assign Cit6x6 = (Jit6x6 & Qit6x6);
assign Qit6x6 = (Oht6x6 | Ninnv6);
assign Oht6x6 = (Rje7z6[28] | Xit6x6);
assign Jit6x6 = (~(Ofnnv6 & Xit6x6));
assign Fgt6x6 = (Ejt6x6 & Ljt6x6);
assign Ljt6x6 = (~(J73ov6 & Em3ov6));
assign Em3ov6 = (Ue3jw6 ^ Dte7z6[1]);
assign Ue3jw6 = (T3cdt6 ? V1c7z6[4] : Et3ov6);
assign Ejt6x6 = (~(R6ziw6 & Od3ov6));
assign Od3ov6 = (Z8q6x6 ^ Dte7z6[1]);
assign Z8q6x6 = (T3cdt6 ? V1c7z6[20] : Myp6x6);
assign Rft6x6 = (Sjt6x6 & Zjt6x6);
assign Zjt6x6 = (Gkt6x6 & Nkt6x6);
assign Nkt6x6 = (~(F7ziw6 & Xe3ov6));
assign Xe3ov6 = (Ukt6x6 ^ Dte7z6[1]);
assign Gkt6x6 = (~(T0ziw6 & Rje7z6[28]));
assign Sjt6x6 = (Blt6x6 & Ilt6x6);
assign Ilt6x6 = (Ryfov6 | Plt6x6);
assign Blt6x6 = (~(L0g7z6[28] & J2ziw6));
assign Dft6x6 = (Wlt6x6 & Dmt6x6);
assign Dmt6x6 = (Kmt6x6 & Rmt6x6);
assign Rmt6x6 = (Ymt6x6 & Fnt6x6);
assign Fnt6x6 = (~(Cqf7z6[12] & Q2ziw6));
assign Ymt6x6 = (~(L0g7z6[12] & O1ziw6));
assign Kmt6x6 = (Mnt6x6 & Tnt6x6);
assign Tnt6x6 = (~(U4ziw6 & V1c7z6[28]));
assign Mnt6x6 = (~(B5ziw6 & H9gdt6));
assign Wlt6x6 = (Aot6x6 & Hot6x6);
assign Hot6x6 = (Oot6x6 & Vot6x6);
assign Vot6x6 = (~(Z3ziw6 & E3c7z6[3]));
assign Oot6x6 = (~(Vzkdt6 & Oztiw6));
assign Aot6x6 = (D43ov6 & T7ziw6);
assign D43ov6 = (Cpt6x6 & Jpt6x6);
assign Jpt6x6 = (~(Qpt6x6 & Rzmnv6));
assign Qpt6x6 = (~(Yzmnv6 | Icziw6));
assign Cpt6x6 = (~(Xpt6x6 & Ubziw6));
assign Xpt6x6 = (~(Rzmnv6 ^ Yzmnv6));
assign Yzmnv6 = (Eqt6x6 ^ Mennv6);
assign Eqt6x6 = (~(Lqt6x6 & Sqt6x6));
assign Sqt6x6 = (Zqt6x6 & Grt6x6);
assign Grt6x6 = (Nrt6x6 & Urt6x6);
assign Urt6x6 = (~(Yxf7z6[30] & Su0jw6));
assign Nrt6x6 = (Bst6x6 & Ist6x6);
assign Ist6x6 = (~(Yxf7z6[28] & Nv0jw6));
assign Bst6x6 = (~(Yxf7z6[29] & Uv0jw6));
assign Zqt6x6 = (Pst6x6 & Wst6x6);
assign Wst6x6 = (~(Pw0jw6 & Yxf7z6[31]));
assign Pst6x6 = (~(Ukt6x6 & Rdziw6));
assign Ukt6x6 = (T3cdt6 ? V1c7z6[28] : Uu3ov6);
assign Lqt6x6 = (Dtt6x6 & Ktt6x6);
assign Ktt6x6 = (Rtt6x6 & Ytt6x6);
assign Ytt6x6 = (~(Onf7z6[28] & My0jw6));
assign Rtt6x6 = (Fut6x6 & Mut6x6);
assign Mut6x6 = (~(Hz0jw6 & Kxb7z6[28]));
assign Fut6x6 = (~(Oz0jw6 & Fhc7z6[28]));
assign Dtt6x6 = (Tut6x6 & Avt6x6);
assign Avt6x6 = (~(Alf7z6[12] & J01jw6));
assign Tut6x6 = (~(Alf7z6[28] & Q01jw6));
assign Rzmnv6 = (~(Hvt6x6 ^ Tennv6));
assign Tennv6 = (!Dte7z6[0]);
assign Hvt6x6 = (~(Ovt6x6 & Vvt6x6));
assign Vvt6x6 = (~(Yxf7z6[12] & Laziw6));
assign Ovt6x6 = (Cwt6x6 & Jwt6x6);
assign Jwt6x6 = (~(Yxf7z6[28] & Gbziw6));
assign Cwt6x6 = (~(Kxb7z6[28] & Nbziw6));
assign Xbt6x6 = (Qwt6x6 & Xwt6x6);
assign Xwt6x6 = (~(Pw9ov6 & Kxb7z6[28]));
assign Qwt6x6 = (Ext6x6 & Lxt6x6);
assign Lxt6x6 = (~(Kx9ov6 & vis_pc_o[28]));
assign Ext6x6 = (~(Gli7z6[28] & Rx9ov6));
assign Amy7v6 = (~(Sxt6x6 & Zxt6x6));
assign Zxt6x6 = (Gyt6x6 & Nyt6x6);
assign Nyt6x6 = (~(Kx9ov6 & vis_pc_o[30]));
assign Kx9ov6 = (Uyt6x6 & Qsq6x6);
assign Gyt6x6 = (Bzt6x6 & Izt6x6);
assign Izt6x6 = (~(Uv9ov6 & Eu97z6));
assign Uv9ov6 = (Uyt6x6 & C3yiw6);
assign C3yiw6 = (!Qsq6x6);
assign Qsq6x6 = (~(Pzt6x6 & Gt2jw6));
assign Pzt6x6 = (Wzt6x6 & D0u6x6);
assign Uyt6x6 = (K0u6x6 & R0u6x6);
assign K0u6x6 = (Ut2jw6 & Y0u6x6);
assign Bzt6x6 = (Eu9ov6 | F1u6x6);
assign Eu9ov6 = (~(M1u6x6 & T1u6x6));
assign M1u6x6 = (Y0u6x6 & A2u6x6);
assign Sxt6x6 = (H2u6x6 & O2u6x6);
assign O2u6x6 = (~(Pw9ov6 & Kxb7z6[30]));
assign H2u6x6 = (V2u6x6 & C3u6x6);
assign C3u6x6 = (~(Rx9ov6 & Gli7z6[30]));
assign Rx9ov6 = (~(J3u6x6 | Ut2jw6));
assign Ut2jw6 = (~(Q3u6x6 & Vs9ov6));
assign Q3u6x6 = (~(X3u6x6 & E4u6x6));
assign E4u6x6 = (L4u6x6 & S4u6x6);
assign S4u6x6 = (~(Ffadt6 | Tuddt6));
assign L4u6x6 = (Rihov6 & Z4u6x6);
assign Z4u6x6 = (~(G5u6x6 & N5u6x6));
assign N5u6x6 = (U5u6x6 & Kkmhw6);
assign G5u6x6 = (B6u6x6 & Ijmhw6);
assign Ijmhw6 = (!C9mov6);
assign C9mov6 = (I6u6x6 & Nneet6);
assign I6u6x6 = (O5a7z6 & P6u6x6);
assign B6u6x6 = (~(W6u6x6 & D7u6x6));
assign X3u6x6 = (K7u6x6 & Mlmhw6);
assign Mlmhw6 = (R7u6x6 & E1wnv6);
assign R7u6x6 = (Ldo7v6 & S2onv6);
assign K7u6x6 = (Zhbdt6 & Y7u6x6);
assign J3u6x6 = (~(R0u6x6 & Y0u6x6));
assign V2u6x6 = (~(Gv9ov6 & Fi4ov6));
assign Fi4ov6 = (Gninv6 ? Gli7z6[30] : Eu97z6);
assign Eu97z6 = (~(F8u6x6 & M8u6x6));
assign M8u6x6 = (~(Nqyiw6 & Acxnv6));
assign Nqyiw6 = (!Z11jw6);
assign F8u6x6 = (T8u6x6 & A9u6x6);
assign A9u6x6 = (~(Pdc7z6[30] & Ouyiw6));
assign T8u6x6 = (~(Vuyiw6 & H9u6x6));
assign H9u6x6 = (~(O9u6x6 & V9u6x6));
assign V9u6x6 = (Cau6x6 & Jau6x6);
assign Jau6x6 = (Qau6x6 & Xau6x6);
assign Xau6x6 = (Ebu6x6 & Lbu6x6);
assign Lbu6x6 = (~(Sbu6x6 & Uxyiw6));
assign Sbu6x6 = (Kxb7z6[30] & Zbu6x6);
assign Ebu6x6 = (~(Iv3ov6 & Gcu6x6));
assign Gcu6x6 = (~(Ncu6x6 & Quziw6));
assign Quziw6 = (Kzyiw6 & Ucu6x6);
assign Ucu6x6 = (Rw3ov6 | Bdu6x6);
assign Kzyiw6 = (Wdu6x6 ? Pdu6x6 : Idu6x6);
assign Pdu6x6 = (~(Deu6x6 & Fzfov6));
assign Idu6x6 = (Mzfov6 | Uinnv6);
assign Mzfov6 = (~(Mrbdt6 & Keu6x6));
assign Keu6x6 = (!Reu6x6);
assign Ncu6x6 = (Yeu6x6 & Ffu6x6);
assign Ffu6x6 = (Zbu6x6 | Ninnv6);
assign Zbu6x6 = (Rje7z6[30] | F0ziw6);
assign Yeu6x6 = (~(F0ziw6 & Ofnnv6));
assign Qau6x6 = (Mfu6x6 & Tfu6x6);
assign Tfu6x6 = (Ryfov6 | Agu6x6);
assign Ryfov6 = (~(Hgu6x6 & Wdu6x6));
assign Wdu6x6 = (!V5bov6);
assign Hgu6x6 = (~(Uinnv6 | Deu6x6));
assign Deu6x6 = (Ogu6x6 & Vgu6x6);
assign Vgu6x6 = (Chu6x6 & Jhu6x6);
assign Jhu6x6 = (Qhu6x6 & Xhu6x6);
assign Xhu6x6 = (Eiu6x6 & Liu6x6);
assign Liu6x6 = (Siu6x6 & Ziu6x6);
assign Ziu6x6 = (~(Rje7z6[0] & Cuziw6));
assign Siu6x6 = (~(Rje7z6[2] & Kp1jw6));
assign Eiu6x6 = (Gju6x6 & Nju6x6);
assign Nju6x6 = (~(Rje7z6[3] & Ryh6x6));
assign Gju6x6 = (~(Rje7z6[4] & Et3ov6));
assign Qhu6x6 = (Uju6x6 & Bku6x6);
assign Bku6x6 = (Iku6x6 & Pku6x6);
assign Pku6x6 = (~(Rje7z6[5] & Xs3ov6));
assign Iku6x6 = (~(Rje7z6[8] & Ku3jw6));
assign Uju6x6 = (Wku6x6 & Dlu6x6);
assign Dlu6x6 = (~(Rje7z6[9] & Pn9jw6));
assign Wku6x6 = (~(Rje7z6[10] & Ci4jw6));
assign Chu6x6 = (Klu6x6 & Rlu6x6);
assign Rlu6x6 = (Ylu6x6 & Fmu6x6);
assign Fmu6x6 = (Mmu6x6 & Tmu6x6);
assign Tmu6x6 = (~(Rje7z6[11] & Pebjw6));
assign Mmu6x6 = (~(Rje7z6[12] & X2h6x6));
assign Ylu6x6 = (Anu6x6 & Hnu6x6);
assign Hnu6x6 = (~(Rje7z6[13] & Dok6x6));
assign Anu6x6 = (~(Rje7z6[14] & Zbn6x6));
assign Klu6x6 = (Onu6x6 & Vnu6x6);
assign Vnu6x6 = (Cou6x6 & Jou6x6);
assign Jou6x6 = (~(Rje7z6[16] & Hr8jw6));
assign Cou6x6 = (~(Rje7z6[17] & Oiajw6));
assign Onu6x6 = (Qou6x6 & Xou6x6);
assign Xou6x6 = (~(Rje7z6[18] & Ew5jw6));
assign Qou6x6 = (~(Rje7z6[19] & O9cjw6));
assign Ogu6x6 = (Epu6x6 & Lpu6x6);
assign Lpu6x6 = (Spu6x6 & Zpu6x6);
assign Zpu6x6 = (Gqu6x6 & Nqu6x6);
assign Nqu6x6 = (Uqu6x6 & Bru6x6);
assign Bru6x6 = (~(Rje7z6[20] & Myp6x6));
assign Uqu6x6 = (~(Rje7z6[21] & Csj6x6));
assign Gqu6x6 = (Iru6x6 & Pru6x6);
assign Pru6x6 = (~(Rje7z6[23] & Nap6x6));
assign Iru6x6 = (~(Rje7z6[24] & T9kov6));
assign Spu6x6 = (Wru6x6 & Dsu6x6);
assign Dsu6x6 = (Ksu6x6 & Rsu6x6);
assign Rsu6x6 = (~(Rje7z6[25] & A07jw6));
assign Ksu6x6 = (~(Rje7z6[26] & Qs3ov6));
assign Wru6x6 = (Ysu6x6 & Ftu6x6);
assign Ftu6x6 = (~(Rje7z6[27] & St3ov6));
assign Ysu6x6 = (~(Rje7z6[29] & Lt3ov6));
assign Epu6x6 = (Mtu6x6 & Ttu6x6);
assign Ttu6x6 = (Auu6x6 & Huu6x6);
assign Huu6x6 = (Ouu6x6 & Vuu6x6);
assign Vuu6x6 = (~(Rje7z6[28] & Uu3ov6));
assign Ouu6x6 = (~(Rje7z6[6] & Nu3ov6));
assign Auu6x6 = (Cvu6x6 & Jvu6x6);
assign Jvu6x6 = (~(Rje7z6[22] & Yfm6x6));
assign Cvu6x6 = (~(Rje7z6[30] & Iv3ov6));
assign Mtu6x6 = (Qvu6x6 & Xvu6x6);
assign Xvu6x6 = (~(Rje7z6[1] & Se2jw6));
assign Qvu6x6 = (Ewu6x6 & Lwu6x6);
assign Lwu6x6 = (~(Rje7z6[7] & Bv3ov6));
assign Ewu6x6 = (~(Rje7z6[15] & M85jw6));
assign Mfu6x6 = (~(T0ziw6 & Rje7z6[30]));
assign T0ziw6 = (Swu6x6 & Zwu6x6);
assign Zwu6x6 = (~(Gxu6x6 & Evziw6));
assign Gxu6x6 = (~(Nxu6x6 & Mrbdt6));
assign Nxu6x6 = (Reu6x6 & V5bov6);
assign V5bov6 = (~(Uxu6x6 & Byu6x6));
assign Uxu6x6 = (~(Yvbov6 & Iyu6x6));
assign Iyu6x6 = (~(Pyu6x6 & Wyu6x6));
assign Wyu6x6 = (Dzu6x6 | Ntbov6);
assign Yvbov6 = (~(Kzu6x6 & Rzu6x6));
assign Rzu6x6 = (Yzu6x6 & F0v6x6);
assign F0v6x6 = (M0v6x6 | T0v6x6);
assign Yzu6x6 = (A1v6x6 | H1v6x6);
assign Kzu6x6 = (O1v6x6 & V1v6x6);
assign V1v6x6 = (C2v6x6 | J2v6x6);
assign O1v6x6 = (Q2v6x6 | X2v6x6);
assign Reu6x6 = (~(E3v6x6 & L3v6x6));
assign L3v6x6 = (S3v6x6 & Z3v6x6);
assign Z3v6x6 = (G4v6x6 & N4v6x6);
assign N4v6x6 = (U4v6x6 & B5v6x6);
assign B5v6x6 = (I5v6x6 & P5v6x6);
assign P5v6x6 = (~(Fx3ov6 & Fq1jw6));
assign Fx3ov6 = (!Kp1jw6);
assign Kp1jw6 = (~(W5v6x6 & D6v6x6));
assign D6v6x6 = (~(K6v6x6 & R6v6x6));
assign R6v6x6 = (~(Y6v6x6 & F7v6x6));
assign F7v6x6 = (M7v6x6 & T7v6x6);
assign T7v6x6 = (C2v6x6 | A8v6x6);
assign M7v6x6 = (M0v6x6 | J2v6x6);
assign Y6v6x6 = (H8v6x6 & O8v6x6);
assign O8v6x6 = (A1v6x6 | V8v6x6);
assign H8v6x6 = (Q2v6x6 | C9v6x6);
assign K6v6x6 = (~(Dzu6x6 ^ J9v6x6));
assign W5v6x6 = (~(Xrbov6 & Q9v6x6));
assign Q9v6x6 = (Dzu6x6 | J9v6x6);
assign J9v6x6 = (X9v6x6 & Eav6x6);
assign X9v6x6 = (Zav6x6 ? Sav6x6 : Lav6x6);
assign I5v6x6 = (~(Yw3ov6 & J17jw6));
assign J17jw6 = (~(Js8jw6 & Gbv6x6));
assign Yw3ov6 = (!A07jw6);
assign A07jw6 = (~(Nbv6x6 & Ubv6x6));
assign Ubv6x6 = (~(Bcv6x6 & Icv6x6));
assign Icv6x6 = (~(Pcv6x6 & Wcv6x6));
assign Wcv6x6 = (Ddv6x6 & Kdv6x6);
assign Kdv6x6 = (A1v6x6 | Rdv6x6);
assign Ddv6x6 = (Q2v6x6 | Ydv6x6);
assign Pcv6x6 = (Fev6x6 & Mev6x6);
assign Mev6x6 = (C2v6x6 | Tev6x6);
assign Fev6x6 = (M0v6x6 | Afv6x6);
assign Bcv6x6 = (~(Dzu6x6 ^ Hfv6x6));
assign Nbv6x6 = (~(Xrbov6 & Ofv6x6));
assign Ofv6x6 = (Dzu6x6 | Hfv6x6);
assign Hfv6x6 = (Vfv6x6 & Cgv6x6);
assign Cgv6x6 = (Jgv6x6 | Qgv6x6);
assign U4v6x6 = (Xgv6x6 & Ehv6x6);
assign Ehv6x6 = (Iv3ov6 | F0ziw6);
assign Xgv6x6 = (~(Hy3ov6 & Rh2jw6));
assign Rh2jw6 = (!Uf2jw6);
assign Uf2jw6 = (~(Fq1jw6 & Lhv6x6));
assign Lhv6x6 = (~(M0ziw6 & Lvziw6));
assign Fq1jw6 = (!Vr1jw6);
assign Vr1jw6 = (C53jw6 | Shv6x6);
assign Hy3ov6 = (!Se2jw6);
assign G4v6x6 = (Zhv6x6 & Giv6x6);
assign Giv6x6 = (Niv6x6 & Uiv6x6);
assign Uiv6x6 = (~(Ay3ov6 & G3i6x6));
assign G3i6x6 = (!Tzh6x6);
assign Tzh6x6 = (~(P83jw6 & Bjv6x6));
assign Bjv6x6 = (~(Shv6x6 & M0ziw6));
assign P83jw6 = (!C53jw6);
assign Ay3ov6 = (!Ryh6x6);
assign Ryh6x6 = (~(Ijv6x6 & Pjv6x6));
assign Pjv6x6 = (~(Wjv6x6 & Dkv6x6));
assign Dkv6x6 = (~(Kkv6x6 & Rkv6x6));
assign Rkv6x6 = (Ykv6x6 & Flv6x6);
assign Flv6x6 = (Q2v6x6 | A8v6x6);
assign Ykv6x6 = (C2v6x6 | Mlv6x6);
assign Kkv6x6 = (Tlv6x6 & Amv6x6);
assign Amv6x6 = (A1v6x6 | C9v6x6);
assign Tlv6x6 = (M0v6x6 | V8v6x6);
assign Wjv6x6 = (~(Dzu6x6 ^ Hmv6x6));
assign Ijv6x6 = (~(Xrbov6 & Omv6x6));
assign Omv6x6 = (Dzu6x6 | Hmv6x6);
assign Hmv6x6 = (Vmv6x6 & Eav6x6);
assign Vmv6x6 = (Zav6x6 ? Jnv6x6 : Cnv6x6);
assign Niv6x6 = (C53jw6 | Et3ov6);
assign Et3ov6 = (Xnv6x6 ? Xrbov6 : Qnv6x6);
assign Xnv6x6 = (Eov6x6 & Lov6x6);
assign Lov6x6 = (~(Sov6x6 & Cnv6x6));
assign Qnv6x6 = (~(Zov6x6 & Gpv6x6));
assign Gpv6x6 = (Npv6x6 & Upv6x6);
assign Upv6x6 = (A1v6x6 | A8v6x6);
assign Npv6x6 = (Q2v6x6 | Mlv6x6);
assign Zov6x6 = (Bqv6x6 & Iqv6x6);
assign Iqv6x6 = (C2v6x6 | Pqv6x6);
assign Bqv6x6 = (M0v6x6 | C9v6x6);
assign C53jw6 = (~(Zy3jw6 & Wqv6x6));
assign Wqv6x6 = (~(Drv6x6 & Lvziw6));
assign Zhv6x6 = (Krv6x6 & Rrv6x6);
assign Rrv6x6 = (Uvi6x6 | Xs3ov6);
assign Xs3ov6 = (Fsv6x6 ? Xrbov6 : Yrv6x6);
assign Fsv6x6 = (Eov6x6 & Msv6x6);
assign Msv6x6 = (~(Sov6x6 & Lav6x6));
assign Yrv6x6 = (~(Tsv6x6 & Atv6x6));
assign Atv6x6 = (Htv6x6 & Otv6x6);
assign Otv6x6 = (M0v6x6 | A8v6x6);
assign A8v6x6 = (Vtv6x6 & Cuv6x6);
assign Cuv6x6 = (Juv6x6 | Quv6x6);
assign Vtv6x6 = (Xuv6x6 & Evv6x6);
assign Evv6x6 = (Lvv6x6 | Svv6x6);
assign Xuv6x6 = (~(Zvv6x6 & Gwv6x6));
assign Htv6x6 = (A1v6x6 | Mlv6x6);
assign Tsv6x6 = (Nwv6x6 & Uwv6x6);
assign Uwv6x6 = (Q2v6x6 | Pqv6x6);
assign Nwv6x6 = (C2v6x6 | Bxv6x6);
assign Uvi6x6 = (~(Knl6x6 & Ixv6x6));
assign Ixv6x6 = (~(Pxv6x6 & Lvziw6));
assign Knl6x6 = (!Skl6x6);
assign Krv6x6 = (Skl6x6 | Nu3ov6);
assign Skl6x6 = (~(Zy3jw6 & Wxv6x6));
assign Wxv6x6 = (~(Shv6x6 & Drv6x6));
assign S3v6x6 = (Dyv6x6 & Kyv6x6);
assign Kyv6x6 = (Ryv6x6 & Yyv6x6);
assign Yyv6x6 = (Fzv6x6 & Mzv6x6);
assign Mzv6x6 = (J9o6x6 | Bv3ov6);
assign J9o6x6 = (~(Zy3jw6 & Tzv6x6));
assign Tzv6x6 = (~(Pxv6x6 & Shv6x6));
assign Fzv6x6 = (~(Vy3ov6 & Zy3jw6));
assign Zy3jw6 = (!Mv3jw6);
assign Vy3ov6 = (!Ku3jw6);
assign Ku3jw6 = (~(A0w6x6 & H0w6x6));
assign H0w6x6 = (~(O0w6x6 & V0w6x6));
assign V0w6x6 = (~(C1w6x6 & J1w6x6));
assign J1w6x6 = (Q1w6x6 & X1w6x6);
assign X1w6x6 = (M0v6x6 | Bxv6x6);
assign Q1w6x6 = (E2w6x6 & L2w6x6);
assign E2w6x6 = (C2v6x6 | S2w6x6);
assign C1w6x6 = (Z2w6x6 & G3w6x6);
assign G3w6x6 = (A1v6x6 | N3w6x6);
assign Z2w6x6 = (Q2v6x6 | U3w6x6);
assign O0w6x6 = (P4w6x6 ? I4w6x6 : B4w6x6);
assign A0w6x6 = (P4w6x6 | Byu6x6);
assign Ryv6x6 = (W4w6x6 & D5w6x6);
assign D5w6x6 = (~(Oy3ov6 & Oq9jw6));
assign Oq9jw6 = (!Ro9jw6);
assign Ro9jw6 = (~(Iv8jw6 & K5w6x6));
assign K5w6x6 = (~(Gbv6x6 & Lvziw6));
assign Gbv6x6 = (R5w6x6 & Y5w6x6);
assign Y5w6x6 = (~(F6w6x6 & M6w6x6));
assign F6w6x6 = (T6w6x6 & A7w6x6);
assign Oy3ov6 = (!Pn9jw6);
assign Pn9jw6 = (~(H7w6x6 & O7w6x6));
assign O7w6x6 = (~(V7w6x6 & C8w6x6));
assign C8w6x6 = (~(J8w6x6 & Q8w6x6));
assign Q8w6x6 = (X8w6x6 & E9w6x6);
assign E9w6x6 = (C2v6x6 | L9w6x6);
assign X8w6x6 = (S9w6x6 & L2w6x6);
assign S9w6x6 = (Q2v6x6 | S2w6x6);
assign J8w6x6 = (Z9w6x6 & Gaw6x6);
assign Gaw6x6 = (M0v6x6 | N3w6x6);
assign Z9w6x6 = (A1v6x6 | U3w6x6);
assign V7w6x6 = (Naw6x6 ? I4w6x6 : B4w6x6);
assign H7w6x6 = (Byu6x6 | Naw6x6);
assign Naw6x6 = (P4w6x6 & Uaw6x6);
assign Uaw6x6 = (~(Bbw6x6 & Qgv6x6));
assign W4w6x6 = (~(Z04ov6 & Bl4jw6));
assign Bl4jw6 = (!Ej4jw6);
assign Ej4jw6 = (~(G4h6x6 & Ibw6x6));
assign Ibw6x6 = (~(Shv6x6 & R5w6x6));
assign Z04ov6 = (!Ci4jw6);
assign Ci4jw6 = (~(Pbw6x6 & Wbw6x6));
assign Wbw6x6 = (~(Dcw6x6 & Kcw6x6));
assign Kcw6x6 = (~(Rcw6x6 & Ycw6x6));
assign Ycw6x6 = (Fdw6x6 & Mdw6x6);
assign Mdw6x6 = (Q2v6x6 | L9w6x6);
assign Fdw6x6 = (Tdw6x6 & L2w6x6);
assign Tdw6x6 = (A1v6x6 | S2w6x6);
assign Rcw6x6 = (Aew6x6 & Hew6x6);
assign Hew6x6 = (C2v6x6 | Oew6x6);
assign Aew6x6 = (M0v6x6 | U3w6x6);
assign Dcw6x6 = (Vew6x6 ? I4w6x6 : B4w6x6);
assign Pbw6x6 = (Byu6x6 | Vew6x6);
assign Vew6x6 = (P4w6x6 & Cfw6x6);
assign Cfw6x6 = (~(Bbw6x6 & Sav6x6));
assign Dyv6x6 = (Jfw6x6 & Qfw6x6);
assign Qfw6x6 = (Xfw6x6 & Egw6x6);
assign Egw6x6 = (~(S04ov6 & Ohbjw6));
assign Ohbjw6 = (!Rfbjw6);
assign Rfbjw6 = (~(G4h6x6 & Lgw6x6));
assign Lgw6x6 = (~(Sgw6x6 & Shv6x6));
assign Sgw6x6 = (R5w6x6 & M0ziw6);
assign S04ov6 = (!Pebjw6);
assign Pebjw6 = (~(Zgw6x6 & Ghw6x6));
assign Ghw6x6 = (~(Nhw6x6 & Uhw6x6));
assign Uhw6x6 = (~(Biw6x6 & Iiw6x6));
assign Iiw6x6 = (Piw6x6 & Wiw6x6);
assign Wiw6x6 = (A1v6x6 | L9w6x6);
assign Piw6x6 = (Djw6x6 & L2w6x6);
assign Djw6x6 = (M0v6x6 | S2w6x6);
assign S2w6x6 = (Kjw6x6 & Rjw6x6);
assign Rjw6x6 = (Yjw6x6 & Fkw6x6);
assign Fkw6x6 = (Mkw6x6 | Tkw6x6);
assign Yjw6x6 = (Lvv6x6 | Alw6x6);
assign Kjw6x6 = (Hlw6x6 & Olw6x6);
assign Olw6x6 = (~(Vlw6x6 & Cmw6x6));
assign Hlw6x6 = (~(Zvv6x6 & Jmw6x6));
assign Biw6x6 = (Qmw6x6 & Xmw6x6);
assign Xmw6x6 = (Q2v6x6 | Oew6x6);
assign Qmw6x6 = (C2v6x6 | Enw6x6);
assign Nhw6x6 = (Lnw6x6 ? I4w6x6 : B4w6x6);
assign Zgw6x6 = (Byu6x6 | Lnw6x6);
assign Lnw6x6 = (P4w6x6 & Snw6x6);
assign Snw6x6 = (~(Bbw6x6 & Jnv6x6));
assign Xfw6x6 = (~(N14ov6 & G4h6x6));
assign G4h6x6 = (~(Mv3jw6 & Znw6x6));
assign Znw6x6 = (~(M6w6x6 & Iv8jw6));
assign Mv3jw6 = (~(Gow6x6 & Iv8jw6));
assign Gow6x6 = (~(R5w6x6 & Lvziw6));
assign N14ov6 = (!X2h6x6);
assign X2h6x6 = (~(Now6x6 & Uow6x6));
assign Uow6x6 = (~(Bpw6x6 & Ipw6x6));
assign Ipw6x6 = (~(Ppw6x6 & Wpw6x6));
assign Wpw6x6 = (Dqw6x6 & Kqw6x6);
assign Kqw6x6 = (A1v6x6 | Oew6x6);
assign Dqw6x6 = (Rqw6x6 & L2w6x6);
assign Rqw6x6 = (M0v6x6 | L9w6x6);
assign L9w6x6 = (Yqw6x6 & Frw6x6);
assign Frw6x6 = (Mrw6x6 & Trw6x6);
assign Trw6x6 = (Mkw6x6 | Asw6x6);
assign Mrw6x6 = (Lvv6x6 | Hsw6x6);
assign Yqw6x6 = (Osw6x6 & Vsw6x6);
assign Vsw6x6 = (~(Vlw6x6 & Ctw6x6));
assign Osw6x6 = (~(Zvv6x6 & Jtw6x6));
assign Ppw6x6 = (Qtw6x6 & Xtw6x6);
assign Xtw6x6 = (Q2v6x6 | Enw6x6);
assign Qtw6x6 = (C2v6x6 | Euw6x6);
assign Bpw6x6 = (Luw6x6 ? I4w6x6 : B4w6x6);
assign Now6x6 = (Byu6x6 | Luw6x6);
assign Luw6x6 = (P4w6x6 & Suw6x6);
assign Suw6x6 = (~(Bbw6x6 & Zuw6x6));
assign Jfw6x6 = (Gvw6x6 & Nvw6x6);
assign Nvw6x6 = (~(G14ov6 & Jrk6x6));
assign Jrk6x6 = (!Fpk6x6);
assign Fpk6x6 = (~(Ffn6x6 & Uvw6x6));
assign Uvw6x6 = (~(Bww6x6 & Pxv6x6));
assign Bww6x6 = (R5w6x6 & Lvziw6);
assign G14ov6 = (!Dok6x6);
assign Dok6x6 = (~(Iww6x6 & Pww6x6));
assign Pww6x6 = (~(Www6x6 & Dxw6x6));
assign Dxw6x6 = (~(Kxw6x6 & Rxw6x6));
assign Rxw6x6 = (Yxw6x6 & Fyw6x6);
assign Fyw6x6 = (A1v6x6 | Enw6x6);
assign Yxw6x6 = (Myw6x6 & L2w6x6);
assign Myw6x6 = (M0v6x6 | Oew6x6);
assign Oew6x6 = (Tyw6x6 & Azw6x6);
assign Azw6x6 = (Hzw6x6 & Ozw6x6);
assign Ozw6x6 = (Mkw6x6 | Vzw6x6);
assign Hzw6x6 = (Lvv6x6 | C0x6x6);
assign Tyw6x6 = (J0x6x6 & Q0x6x6);
assign Q0x6x6 = (~(Vlw6x6 & X0x6x6));
assign J0x6x6 = (E1x6x6 | L1x6x6);
assign Kxw6x6 = (S1x6x6 & Z1x6x6);
assign Z1x6x6 = (Q2v6x6 | Euw6x6);
assign S1x6x6 = (C2v6x6 | G2x6x6);
assign Www6x6 = (N2x6x6 ? I4w6x6 : B4w6x6);
assign Iww6x6 = (Byu6x6 | N2x6x6);
assign N2x6x6 = (P4w6x6 & U2x6x6);
assign U2x6x6 = (~(Bbw6x6 & B3x6x6));
assign Gvw6x6 = (~(P24ov6 & Ffn6x6));
assign Ffn6x6 = (!Bdn6x6);
assign Bdn6x6 = (~(Iv8jw6 & I3x6x6));
assign I3x6x6 = (~(P3x6x6 & Shv6x6));
assign P3x6x6 = (R5w6x6 & Drv6x6);
assign P24ov6 = (!Zbn6x6);
assign Zbn6x6 = (~(W3x6x6 & D4x6x6));
assign D4x6x6 = (~(K4x6x6 & R4x6x6));
assign R4x6x6 = (~(Y4x6x6 & F5x6x6));
assign F5x6x6 = (M5x6x6 & T5x6x6);
assign T5x6x6 = (A1v6x6 | Euw6x6);
assign M5x6x6 = (A6x6x6 & L2w6x6);
assign A6x6x6 = (M0v6x6 | Enw6x6);
assign Enw6x6 = (H6x6x6 & O6x6x6);
assign O6x6x6 = (V6x6x6 & C7x6x6);
assign C7x6x6 = (Mkw6x6 | J7x6x6);
assign V6x6x6 = (Lvv6x6 | Q7x6x6);
assign H6x6x6 = (X7x6x6 & E8x6x6);
assign E8x6x6 = (~(Vlw6x6 & L8x6x6));
assign X7x6x6 = (E1x6x6 | S8x6x6);
assign Y4x6x6 = (Z8x6x6 & G9x6x6);
assign G9x6x6 = (Q2v6x6 | G2x6x6);
assign Z8x6x6 = (C2v6x6 | N9x6x6);
assign K4x6x6 = (U9x6x6 ? I4w6x6 : B4w6x6);
assign W3x6x6 = (Byu6x6 | U9x6x6);
assign U9x6x6 = (P4w6x6 & Bax6x6);
assign Bax6x6 = (~(Bbw6x6 & Iax6x6));
assign Bbw6x6 = (Pax6x6 & Wax6x6);
assign Pax6x6 = (~(Dbx6x6 | Kbx6x6));
assign P4w6x6 = (Rbx6x6 | Ybx6x6);
assign E3v6x6 = (Fcx6x6 & Mcx6x6);
assign Mcx6x6 = (Tcx6x6 & Adx6x6);
assign Adx6x6 = (Hdx6x6 & Odx6x6);
assign Odx6x6 = (Vdx6x6 & Cex6x6);
assign Cex6x6 = (~(I24ov6 & Xa5jw6));
assign Xa5jw6 = (!O95jw6);
assign O95jw6 = (~(Iv8jw6 & Jex6x6));
assign Jex6x6 = (~(Qex6x6 & Pxv6x6));
assign Qex6x6 = (R5w6x6 & Shv6x6);
assign Shv6x6 = (Xex6x6 & Lvziw6);
assign Vdx6x6 = (~(D34ov6 & Imajw6));
assign Imajw6 = (!Qjajw6);
assign Qjajw6 = (~(Rz5jw6 & Efx6x6));
assign Efx6x6 = (~(Js8jw6 & M0ziw6));
assign D34ov6 = (!Oiajw6);
assign Oiajw6 = (~(Lfx6x6 & Sfx6x6));
assign Sfx6x6 = (~(Zfx6x6 & Ggx6x6));
assign Ggx6x6 = (~(Ngx6x6 & Ugx6x6));
assign Ugx6x6 = (Bhx6x6 & Ihx6x6);
assign Ihx6x6 = (C2v6x6 | Phx6x6);
assign Bhx6x6 = (Whx6x6 & L2w6x6);
assign Whx6x6 = (Q2v6x6 | Dix6x6);
assign Ngx6x6 = (Kix6x6 & Rix6x6);
assign Rix6x6 = (M0v6x6 | N9x6x6);
assign Kix6x6 = (A1v6x6 | Yix6x6);
assign Zfx6x6 = (Fjx6x6 ? I4w6x6 : B4w6x6);
assign Lfx6x6 = (Fjx6x6 | Byu6x6);
assign Fjx6x6 = (~(Mjx6x6 & Tjx6x6));
assign Mjx6x6 = (Akx6x6 & Hkx6x6);
assign Hkx6x6 = (Okx6x6 | Vkx6x6);
assign Akx6x6 = (~(Ybx6x6 & Iax6x6));
assign Hdx6x6 = (Clx6x6 & Jlx6x6);
assign Jlx6x6 = (~(W24ov6 & Rz5jw6));
assign Rz5jw6 = (!Gx5jw6);
assign Gx5jw6 = (~(G2q6x6 & Qlx6x6));
assign Qlx6x6 = (~(Js8jw6 & Xex6x6));
assign W24ov6 = (!Ew5jw6);
assign Ew5jw6 = (~(Xlx6x6 & Emx6x6));
assign Emx6x6 = (~(Lmx6x6 & Smx6x6));
assign Smx6x6 = (~(Zmx6x6 & Gnx6x6));
assign Gnx6x6 = (Nnx6x6 & Unx6x6);
assign Unx6x6 = (Q2v6x6 | Phx6x6);
assign Nnx6x6 = (Box6x6 & L2w6x6);
assign Box6x6 = (A1v6x6 | Dix6x6);
assign Zmx6x6 = (Iox6x6 & Pox6x6);
assign Pox6x6 = (C2v6x6 | Wox6x6);
assign Iox6x6 = (M0v6x6 | Yix6x6);
assign Lmx6x6 = (Dpx6x6 ? I4w6x6 : B4w6x6);
assign Xlx6x6 = (Dpx6x6 | Byu6x6);
assign Dpx6x6 = (~(Tjx6x6 & Kpx6x6));
assign Kpx6x6 = (~(Ybx6x6 & B3x6x6));
assign Tjx6x6 = (Jgv6x6 & Rpx6x6);
assign Rpx6x6 = (Okx6x6 | Sav6x6);
assign Clx6x6 = (~(T44ov6 & Bdcjw6));
assign Bdcjw6 = (!Qacjw6);
assign Qacjw6 = (~(G2q6x6 & Ypx6x6));
assign Ypx6x6 = (~(Fqx6x6 & Js8jw6));
assign T44ov6 = (!O9cjw6);
assign O9cjw6 = (~(Mqx6x6 & Tqx6x6));
assign Tqx6x6 = (~(Arx6x6 & Hrx6x6));
assign Hrx6x6 = (~(Orx6x6 & Vrx6x6));
assign Vrx6x6 = (Csx6x6 & Jsx6x6);
assign Jsx6x6 = (A1v6x6 | Phx6x6);
assign Csx6x6 = (Qsx6x6 & L2w6x6);
assign Qsx6x6 = (M0v6x6 | Dix6x6);
assign Orx6x6 = (Xsx6x6 & Etx6x6);
assign Etx6x6 = (Q2v6x6 | Wox6x6);
assign Xsx6x6 = (C2v6x6 | Ltx6x6);
assign Arx6x6 = (Stx6x6 ? I4w6x6 : B4w6x6);
assign Mqx6x6 = (Stx6x6 | Byu6x6);
assign Stx6x6 = (~(Ztx6x6 & Gux6x6));
assign Gux6x6 = (~(Ybx6x6 & Zuw6x6));
assign Ztx6x6 = (Nux6x6 & Jgv6x6);
assign Nux6x6 = (Okx6x6 | Jnv6x6);
assign Tcx6x6 = (Uux6x6 & Bvx6x6);
assign Bvx6x6 = (Ivx6x6 & Pvx6x6);
assign Pvx6x6 = (~(M44ov6 & G2q6x6));
assign G2q6x6 = (!Ozp6x6);
assign Ozp6x6 = (~(Az7jw6 & Wvx6x6));
assign Wvx6x6 = (~(Js8jw6 & Drv6x6));
assign M44ov6 = (!Myp6x6);
assign Myp6x6 = (~(Dwx6x6 & Kwx6x6));
assign Kwx6x6 = (~(Rwx6x6 & Ywx6x6));
assign Ywx6x6 = (~(Fxx6x6 & Mxx6x6));
assign Mxx6x6 = (Txx6x6 & Ayx6x6);
assign Ayx6x6 = (A1v6x6 | Wox6x6);
assign Txx6x6 = (Hyx6x6 & L2w6x6);
assign Hyx6x6 = (M0v6x6 | Phx6x6);
assign Phx6x6 = (Oyx6x6 & Vyx6x6);
assign Vyx6x6 = (Czx6x6 & Jzx6x6);
assign Jzx6x6 = (Mkw6x6 | Qzx6x6);
assign Czx6x6 = (~(Xzx6x6 & E0y6x6));
assign Oyx6x6 = (L0y6x6 & S0y6x6);
assign S0y6x6 = (Juv6x6 | Z0y6x6);
assign L0y6x6 = (~(Zvv6x6 & G1y6x6));
assign Fxx6x6 = (N1y6x6 & U1y6x6);
assign U1y6x6 = (Q2v6x6 | Ltx6x6);
assign N1y6x6 = (C2v6x6 | B2y6x6);
assign Rwx6x6 = (I2y6x6 ? I4w6x6 : B4w6x6);
assign Dwx6x6 = (I2y6x6 | Byu6x6);
assign I2y6x6 = (~(P2y6x6 & W2y6x6));
assign W2y6x6 = (Okx6x6 | Zuw6x6);
assign P2y6x6 = (D3y6x6 & Jgv6x6);
assign D3y6x6 = (~(Ybx6x6 & Jnv6x6));
assign Ivx6x6 = (~(H54ov6 & Pvj6x6));
assign Pvj6x6 = (!Etj6x6);
assign Etj6x6 = (~(Xim6x6 & K3y6x6));
assign K3y6x6 = (~(Pxv6x6 & Js8jw6));
assign H54ov6 = (!Csj6x6);
assign Csj6x6 = (~(R3y6x6 & Y3y6x6));
assign Y3y6x6 = (~(F4y6x6 & M4y6x6));
assign M4y6x6 = (~(T4y6x6 & A5y6x6));
assign A5y6x6 = (H5y6x6 & O5y6x6);
assign O5y6x6 = (A1v6x6 | Ltx6x6);
assign H5y6x6 = (V5y6x6 & L2w6x6);
assign V5y6x6 = (M0v6x6 | Wox6x6);
assign Wox6x6 = (C6y6x6 & J6y6x6);
assign J6y6x6 = (Q6y6x6 & X6y6x6);
assign X6y6x6 = (Mkw6x6 | E7y6x6);
assign Q6y6x6 = (Lvv6x6 | L7y6x6);
assign C6y6x6 = (S7y6x6 & Z7y6x6);
assign Z7y6x6 = (Juv6x6 | G8y6x6);
assign S7y6x6 = (~(Zvv6x6 & N8y6x6));
assign T4y6x6 = (U8y6x6 & B9y6x6);
assign B9y6x6 = (Q2v6x6 | B2y6x6);
assign U8y6x6 = (C2v6x6 | I9y6x6);
assign F4y6x6 = (P9y6x6 ? I4w6x6 : B4w6x6);
assign R3y6x6 = (P9y6x6 | Byu6x6);
assign P9y6x6 = (~(W9y6x6 & Day6x6));
assign Day6x6 = (~(Ybx6x6 & Sav6x6));
assign W9y6x6 = (Kay6x6 & Jgv6x6);
assign Kay6x6 = (Okx6x6 | B3x6x6);
assign B3x6x6 = (!Lav6x6);
assign Uux6x6 = (Ray6x6 & Yay6x6);
assign Yay6x6 = (~(A54ov6 & Xim6x6));
assign Xim6x6 = (!Ahm6x6);
assign Ahm6x6 = (~(Az7jw6 & Fby6x6));
assign Fby6x6 = (~(Mby6x6 & Js8jw6));
assign Mby6x6 = (Drv6x6 & Xex6x6);
assign A54ov6 = (!Yfm6x6);
assign Ray6x6 = (~(J64ov6 & Kcp6x6));
assign Kcp6x6 = (!Pbp6x6);
assign Pbp6x6 = (~(Az7jw6 & Tby6x6));
assign Tby6x6 = (~(Acy6x6 & Pxv6x6));
assign Pxv6x6 = (~(M6w6x6 | A7w6x6));
assign Acy6x6 = (Xex6x6 & Js8jw6);
assign J64ov6 = (!Nap6x6);
assign Nap6x6 = (~(Hcy6x6 & Ocy6x6));
assign Ocy6x6 = (~(Vcy6x6 & Cdy6x6));
assign Cdy6x6 = (~(Jdy6x6 & Qdy6x6));
assign Qdy6x6 = (Xdy6x6 & Eey6x6);
assign Eey6x6 = (C2v6x6 | Rdv6x6);
assign Xdy6x6 = (M0v6x6 | B2y6x6);
assign Jdy6x6 = (Ley6x6 & Sey6x6);
assign Sey6x6 = (A1v6x6 | I9y6x6);
assign Ley6x6 = (Q2v6x6 | Afv6x6);
assign Vcy6x6 = (~(Dzu6x6 ^ Zey6x6));
assign Hcy6x6 = (~(Xrbov6 & Gfy6x6));
assign Gfy6x6 = (Dzu6x6 | Zey6x6);
assign Zey6x6 = (Nfy6x6 & Ufy6x6);
assign Ufy6x6 = (Okx6x6 | Bgy6x6);
assign Fcx6x6 = (Igy6x6 & Pgy6x6);
assign Pgy6x6 = (Wgy6x6 & Dhy6x6);
assign Dhy6x6 = (Khy6x6 & Rhy6x6);
assign Rhy6x6 = (S6s6x6 | Qs3ov6);
assign Qs3ov6 = (Fiy6x6 ? Xrbov6 : Yhy6x6);
assign Fiy6x6 = (Pyu6x6 & Miy6x6);
assign Miy6x6 = (~(Tiy6x6 & Ajy6x6));
assign Tiy6x6 = (Sov6x6 & Hjy6x6);
assign Yhy6x6 = (~(Ojy6x6 & Vjy6x6));
assign Vjy6x6 = (Cky6x6 & Jky6x6);
assign Jky6x6 = (M0v6x6 | Rdv6x6);
assign Cky6x6 = (A1v6x6 | Ydv6x6);
assign Ojy6x6 = (Qky6x6 & Xky6x6);
assign Xky6x6 = (Q2v6x6 | Tev6x6);
assign Qky6x6 = (C2v6x6 | Ely6x6);
assign S6s6x6 = (~(Plt6x6 & Lly6x6));
assign Lly6x6 = (~(Pw7jw6 & Xex6x6));
assign Khy6x6 = (Cxs6x6 | St3ov6);
assign St3ov6 = (Zly6x6 ? Xrbov6 : Sly6x6);
assign Zly6x6 = (Pyu6x6 & Gmy6x6);
assign Gmy6x6 = (~(Nmy6x6 & Ajy6x6));
assign Nmy6x6 = (Umy6x6 & Sov6x6);
assign Umy6x6 = (!Jnv6x6);
assign Jnv6x6 = (~(Hjy6x6 & Bny6x6));
assign Bny6x6 = (~(Vkx6x6 & Zuw6x6));
assign Hjy6x6 = (!Sav6x6);
assign Sly6x6 = (~(Iny6x6 & Pny6x6));
assign Pny6x6 = (Wny6x6 & Doy6x6);
assign Doy6x6 = (M0v6x6 | Ydv6x6);
assign Wny6x6 = (A1v6x6 | Tev6x6);
assign Iny6x6 = (Koy6x6 & Roy6x6);
assign Roy6x6 = (Q2v6x6 | Ely6x6);
assign Koy6x6 = (C2v6x6 | Yoy6x6);
assign Cxs6x6 = (~(Plt6x6 & Fpy6x6));
assign Fpy6x6 = (~(Fqx6x6 & Pw7jw6));
assign Fqx6x6 = (Xex6x6 & M0ziw6);
assign Plt6x6 = (!Xit6x6);
assign Wgy6x6 = (Mpy6x6 & Tpy6x6);
assign Tpy6x6 = (Q71jw6 | Lt3ov6);
assign Lt3ov6 = (Hqy6x6 ? Xrbov6 : Aqy6x6);
assign Hqy6x6 = (Pyu6x6 & Oqy6x6);
assign Oqy6x6 = (~(Vqy6x6 & Ajy6x6));
assign Vqy6x6 = (Sov6x6 & Lav6x6);
assign Lav6x6 = (~(Cry6x6 & Iax6x6));
assign Cry6x6 = (~(Jry6x6 & Cnv6x6));
assign Aqy6x6 = (~(Qry6x6 & Xry6x6));
assign Xry6x6 = (Esy6x6 & Lsy6x6);
assign Lsy6x6 = (M0v6x6 | Ely6x6);
assign Esy6x6 = (A1v6x6 | Yoy6x6);
assign Qry6x6 = (Ssy6x6 & Zsy6x6);
assign Zsy6x6 = (Q2v6x6 | T0v6x6);
assign Ssy6x6 = (C2v6x6 | H1v6x6);
assign Q71jw6 = (~(Agu6x6 & Gty6x6));
assign Gty6x6 = (~(Xit6x6 & M0ziw6));
assign Agu6x6 = (!F0ziw6);
assign F0ziw6 = (Xit6x6 & Xex6x6);
assign Mpy6x6 = (~(C64ov6 & Bp0jw6));
assign Bp0jw6 = (!Lvziw6);
assign C64ov6 = (!Cuziw6);
assign Cuziw6 = (~(Nty6x6 & L2w6x6));
assign Nty6x6 = (~(Sov6x6 & Rvbov6));
assign Rvbov6 = (~(Uty6x6 & Buy6x6));
assign Buy6x6 = (Iuy6x6 & Puy6x6);
assign Puy6x6 = (Q2v6x6 | J2v6x6);
assign Iuy6x6 = (C2v6x6 | V8v6x6);
assign Uty6x6 = (Wuy6x6 & Dvy6x6);
assign Dvy6x6 = (A1v6x6 | X2v6x6);
assign Wuy6x6 = (M0v6x6 | H1v6x6);
assign Igy6x6 = (Kvy6x6 & Rvy6x6);
assign Rvy6x6 = (Uu3ov6 | Xit6x6);
assign Xit6x6 = (Pw7jw6 & Drv6x6);
assign Drv6x6 = (!M6w6x6);
assign M6w6x6 = (Yvy6x6 ^ Fwy6x6);
assign Yvy6x6 = (~(Mwy6x6 & M0ziw6));
assign Uu3ov6 = (Axy6x6 ? Xrbov6 : Twy6x6);
assign Axy6x6 = (Pyu6x6 & Hxy6x6);
assign Hxy6x6 = (~(Oxy6x6 & Ajy6x6));
assign Oxy6x6 = (Sov6x6 & Cnv6x6);
assign Twy6x6 = (~(Vxy6x6 & Cyy6x6));
assign Cyy6x6 = (Jyy6x6 & Qyy6x6);
assign Qyy6x6 = (M0v6x6 | Tev6x6);
assign Tev6x6 = (Xyy6x6 & Ezy6x6);
assign Ezy6x6 = (Lzy6x6 & Szy6x6);
assign Szy6x6 = (Mkw6x6 | Zzy6x6);
assign Lzy6x6 = (Lvv6x6 | G0z6x6);
assign Xyy6x6 = (N0z6x6 & U0z6x6);
assign U0z6x6 = (~(Vlw6x6 & B1z6x6));
assign N0z6x6 = (E1x6x6 | I1z6x6);
assign Jyy6x6 = (A1v6x6 | Ely6x6);
assign Ely6x6 = (P1z6x6 & W1z6x6);
assign W1z6x6 = (D2z6x6 & K2z6x6);
assign K2z6x6 = (Mkw6x6 | R2z6x6);
assign D2z6x6 = (Lvv6x6 | Y2z6x6);
assign P1z6x6 = (F3z6x6 & M3z6x6);
assign M3z6x6 = (~(Vlw6x6 & T3z6x6));
assign F3z6x6 = (E1x6x6 | A4z6x6);
assign Vxy6x6 = (H4z6x6 & O4z6x6);
assign O4z6x6 = (Q2v6x6 | Yoy6x6);
assign H4z6x6 = (C2v6x6 | T0v6x6);
assign Kvy6x6 = (V4z6x6 & C5z6x6);
assign C5z6x6 = (~(X64ov6 & Iv8jw6));
assign X64ov6 = (!Hr8jw6);
assign Hr8jw6 = (~(J5z6x6 & Q5z6x6));
assign Q5z6x6 = (~(X5z6x6 & E6z6x6));
assign E6z6x6 = (~(L6z6x6 & S6z6x6));
assign S6z6x6 = (Z6z6x6 & G7z6x6);
assign G7z6x6 = (C2v6x6 | Dix6x6);
assign Dix6x6 = (N7z6x6 & U7z6x6);
assign U7z6x6 = (B8z6x6 & I8z6x6);
assign I8z6x6 = (Mkw6x6 | P8z6x6);
assign B8z6x6 = (Lvv6x6 | W8z6x6);
assign N7z6x6 = (D9z6x6 & K9z6x6);
assign K9z6x6 = (Juv6x6 | R9z6x6);
assign D9z6x6 = (E1x6x6 | Y9z6x6);
assign Z6z6x6 = (M0v6x6 | G2x6x6);
assign L6z6x6 = (Faz6x6 & Maz6x6);
assign Maz6x6 = (A1v6x6 | N9x6x6);
assign Faz6x6 = (Q2v6x6 | Yix6x6);
assign X5z6x6 = (~(Dzu6x6 ^ Taz6x6));
assign J5z6x6 = (~(Xrbov6 & Abz6x6));
assign Abz6x6 = (Dzu6x6 | Taz6x6);
assign Taz6x6 = (Hbz6x6 & Nfy6x6);
assign Hbz6x6 = (Obz6x6 & Okx6x6);
assign Obz6x6 = (~(Ybx6x6 & Bgy6x6));
assign V4z6x6 = (~(Q64ov6 & Az7jw6));
assign Az7jw6 = (!Pw7jw6);
assign Pw7jw6 = (Js8jw6 & R5w6x6);
assign R5w6x6 = (Vbz6x6 ^ Ccz6x6);
assign Js8jw6 = (!Iv8jw6);
assign Iv8jw6 = (~(Jcz6x6 & Lvziw6));
assign Lvziw6 = (~(Qcz6x6 & Xcz6x6));
assign Xcz6x6 = (Edz6x6 & Ldz6x6);
assign Edz6x6 = (Xex6x6 & Sdz6x6);
assign Sdz6x6 = (Hfnnv6 | Zdz6x6);
assign Hfnnv6 = (~(Gez6x6 & V1c7z6[31]));
assign Gez6x6 = (~(Nez6x6 | Uez6x6));
assign Xex6x6 = (!T6w6x6);
assign T6w6x6 = (Mwy6x6 ^ M0ziw6);
assign M0ziw6 = (!A7w6x6);
assign Qcz6x6 = (~(Ccz6x6 | Bfz6x6));
assign Jcz6x6 = (~(Ifz6x6 ^ Bfz6x6));
assign Bfz6x6 = (~(Pfz6x6 & Wfz6x6));
assign Wfz6x6 = (~(Cgnnv6 & Swu6x6));
assign Cgnnv6 = (~(Dgz6x6 ^ V1c7z6[31]));
assign Dgz6x6 = (Nez6x6 | Uez6x6);
assign Pfz6x6 = (~(V1c7z6[12] & Uxyiw6));
assign Ifz6x6 = (~(Vbz6x6 & Kgz6x6));
assign Kgz6x6 = (!Ccz6x6);
assign Ccz6x6 = (~(Rgz6x6 & Ygz6x6));
assign Ygz6x6 = (~(Qgnnv6 & Swu6x6));
assign Qgnnv6 = (Uez6x6 ^ Nez6x6);
assign Nez6x6 = (!V1c7z6[30]);
assign Uez6x6 = (~(V1c7z6[29] & Fhz6x6));
assign Rgz6x6 = (~(Uxyiw6 & V1c7z6[11]));
assign Vbz6x6 = (Ldz6x6 & Mwy6x6);
assign Mwy6x6 = (Mhz6x6 & Thz6x6);
assign Thz6x6 = (~(Ehnnv6 & Swu6x6));
assign Ehnnv6 = (Aiz6x6 ^ V1c7z6[28]);
assign Mhz6x6 = (~(Uxyiw6 & V1c7z6[9]));
assign Ldz6x6 = (~(Fwy6x6 | A7w6x6));
assign A7w6x6 = (~(Hiz6x6 & Oiz6x6));
assign Oiz6x6 = (~(Lhnnv6 & Swu6x6));
assign Lhnnv6 = (Viz6x6 ^ V1c7z6[27]);
assign Hiz6x6 = (~(Uxyiw6 & V1c7z6[8]));
assign Fwy6x6 = (~(Cjz6x6 & Jjz6x6));
assign Jjz6x6 = (~(Xgnnv6 & Swu6x6));
assign Xgnnv6 = (Fhz6x6 ^ V1c7z6[29]);
assign Fhz6x6 = (Aiz6x6 & V1c7z6[28]);
assign Aiz6x6 = (V1c7z6[27] & Viz6x6);
assign Viz6x6 = (~(Ninnv6 & Evziw6));
assign Ninnv6 = (!Uxyiw6);
assign Cjz6x6 = (~(Uxyiw6 & V1c7z6[10]));
assign Uxyiw6 = (Dy1ov6 & Bqziw6);
assign Q64ov6 = (!T9kov6);
assign T9kov6 = (~(Qjz6x6 & Xjz6x6));
assign Xjz6x6 = (~(Ekz6x6 & Lkz6x6));
assign Lkz6x6 = (~(Skz6x6 & Zkz6x6));
assign Zkz6x6 = (Glz6x6 & Nlz6x6);
assign Nlz6x6 = (Q2v6x6 | Rdv6x6);
assign Rdv6x6 = (Ulz6x6 & Bmz6x6);
assign Bmz6x6 = (Imz6x6 & Pmz6x6);
assign Pmz6x6 = (Mkw6x6 | Wmz6x6);
assign Imz6x6 = (Lvv6x6 | Dnz6x6);
assign Ulz6x6 = (Knz6x6 & Rnz6x6);
assign Rnz6x6 = (~(Vlw6x6 & Ynz6x6));
assign Knz6x6 = (E1x6x6 | Foz6x6);
assign Glz6x6 = (C2v6x6 | Ydv6x6);
assign Ydv6x6 = (Moz6x6 & Toz6x6);
assign Toz6x6 = (Apz6x6 & Hpz6x6);
assign Hpz6x6 = (Mkw6x6 | Opz6x6);
assign Apz6x6 = (Lvv6x6 | Vpz6x6);
assign Moz6x6 = (Cqz6x6 & Jqz6x6);
assign Jqz6x6 = (~(Vlw6x6 & Qqz6x6));
assign Cqz6x6 = (E1x6x6 | Xqz6x6);
assign Skz6x6 = (Erz6x6 & Lrz6x6);
assign Lrz6x6 = (M0v6x6 | I9y6x6);
assign Erz6x6 = (A1v6x6 | Afv6x6);
assign Ekz6x6 = (~(Dzu6x6 ^ Nfy6x6));
assign Qjz6x6 = (~(Xrbov6 & Srz6x6));
assign Srz6x6 = (~(Ajy6x6 & Sov6x6));
assign Swu6x6 = (!Zdz6x6);
assign Zdz6x6 = (Evziw6 & Uinnv6);
assign Uinnv6 = (!Fzfov6);
assign Fzfov6 = (~(Rw3ov6 | Zao6x6));
assign Evziw6 = (!Ofnnv6);
assign Ofnnv6 = (Dy1ov6 & Zrz6x6);
assign Dy1ov6 = (!Rw3ov6);
assign Rw3ov6 = (~(Gsz6x6 & Dte7z6[15]));
assign Cau6x6 = (Nsz6x6 & Usz6x6);
assign Usz6x6 = (Btz6x6 & Itz6x6);
assign Itz6x6 = (~(J73ov6 & Ql3ov6));
assign Ql3ov6 = (Fvl6x6 ^ Dte7z6[1]);
assign Fvl6x6 = (T3cdt6 ? V1c7z6[6] : Nu3ov6);
assign Nu3ov6 = (Wtz6x6 ? Xrbov6 : Ptz6x6);
assign Wtz6x6 = (Eov6x6 & Duz6x6);
assign Duz6x6 = (~(Sov6x6 & Kuz6x6));
assign Eov6x6 = (~(Sov6x6 ^ Eav6x6));
assign Ptz6x6 = (~(Ruz6x6 & Yuz6x6));
assign Yuz6x6 = (Fvz6x6 & Mvz6x6);
assign Mvz6x6 = (M0v6x6 | Mlv6x6);
assign Mlv6x6 = (Tvz6x6 & Awz6x6);
assign Awz6x6 = (Juv6x6 | Hwz6x6);
assign Tvz6x6 = (Owz6x6 & Vwz6x6);
assign Vwz6x6 = (Lvv6x6 | Cxz6x6);
assign Owz6x6 = (~(Zvv6x6 & Jxz6x6));
assign Fvz6x6 = (A1v6x6 | Pqv6x6);
assign Ruz6x6 = (Qxz6x6 & Xxz6x6);
assign Xxz6x6 = (Q2v6x6 | Bxv6x6);
assign Qxz6x6 = (C2v6x6 | N3w6x6);
assign J73ov6 = (!Lf3ov6);
assign Lf3ov6 = (Ubo6x6 | Zho6x6);
assign Btz6x6 = (~(L0g7z6[30] & J2ziw6));
assign J2ziw6 = (~(Eyz6x6 & Lyz6x6));
assign Lyz6x6 = (Syz6x6 & Zgtiw6);
assign Syz6x6 = (~(Zyz6x6 & Gzz6x6));
assign Zyz6x6 = (E4lhw6 & Nzz6x6);
assign Eyz6x6 = (Dx0jw6 & Uzz6x6);
assign Uzz6x6 = (~(Uh2ov6 & Gvtiw6));
assign Nsz6x6 = (B007x6 & I007x6);
assign I007x6 = (~(R6ziw6 & Qe3ov6));
assign Qe3ov6 = (Eqm6x6 ^ Dte7z6[1]);
assign Eqm6x6 = (T3cdt6 ? V1c7z6[22] : Yfm6x6);
assign Yfm6x6 = (~(P007x6 & W007x6));
assign W007x6 = (~(D107x6 & K107x6));
assign K107x6 = (~(R107x6 & Y107x6));
assign Y107x6 = (F207x6 & M207x6);
assign M207x6 = (Q2v6x6 | I9y6x6);
assign I9y6x6 = (T207x6 & A307x6);
assign A307x6 = (H307x6 & O307x6);
assign O307x6 = (~(V307x6 & E0y6x6));
assign E0y6x6 = (~(C407x6 & J407x6));
assign H307x6 = (Lvv6x6 | Zzy6x6);
assign Zzy6x6 = (Q407x6 & X407x6);
assign T207x6 = (E507x6 & L507x6);
assign L507x6 = (~(Vlw6x6 & G1y6x6));
assign G1y6x6 = (~(S507x6 & Z507x6));
assign E507x6 = (~(Zvv6x6 & B1z6x6));
assign B1z6x6 = (~(G607x6 & N607x6));
assign F207x6 = (U607x6 & B707x6);
assign B707x6 = (M0v6x6 | Ltx6x6);
assign Ltx6x6 = (I707x6 & P707x6);
assign P707x6 = (W707x6 & D807x6);
assign D807x6 = (Mkw6x6 | K807x6);
assign W707x6 = (Lvv6x6 | Wmz6x6);
assign Wmz6x6 = (R807x6 & Y807x6);
assign I707x6 = (F907x6 & M907x6);
assign M907x6 = (Juv6x6 | T907x6);
assign F907x6 = (~(Zvv6x6 & Ynz6x6));
assign Ynz6x6 = (~(Aa07x6 & Ha07x6));
assign U607x6 = (A1v6x6 | B2y6x6);
assign B2y6x6 = (Oa07x6 & Va07x6);
assign Va07x6 = (Cb07x6 & Jb07x6);
assign Jb07x6 = (Mkw6x6 | W8z6x6);
assign W8z6x6 = (Qb07x6 & Xb07x6);
assign Qb07x6 = (Ec07x6 & Lc07x6);
assign Cb07x6 = (Lvv6x6 | Opz6x6);
assign Opz6x6 = (Sc07x6 & Zc07x6);
assign Oa07x6 = (Gd07x6 & Nd07x6);
assign Nd07x6 = (Juv6x6 | Y9z6x6);
assign Y9z6x6 = (Ud07x6 & Be07x6);
assign Ud07x6 = (Ie07x6 & Pe07x6);
assign Pe07x6 = (~(Cve7z6[15] & We07x6));
assign Ie07x6 = (~(Dbx6x6 & Neo7v6));
assign Gd07x6 = (~(Zvv6x6 & Qqz6x6));
assign Qqz6x6 = (~(Df07x6 & Kf07x6));
assign R107x6 = (L2w6x6 & Rf07x6);
assign Rf07x6 = (C2v6x6 | Afv6x6);
assign Afv6x6 = (Yf07x6 & Fg07x6);
assign Fg07x6 = (Mg07x6 & Tg07x6);
assign Tg07x6 = (Mkw6x6 | L7y6x6);
assign L7y6x6 = (Ah07x6 & Hh07x6);
assign Mg07x6 = (Lvv6x6 | R2z6x6);
assign R2z6x6 = (Oh07x6 & Vh07x6);
assign Yf07x6 = (Ci07x6 & Ji07x6);
assign Ji07x6 = (~(Vlw6x6 & N8y6x6));
assign N8y6x6 = (~(Qi07x6 & Xi07x6));
assign Ci07x6 = (~(Zvv6x6 & T3z6x6));
assign T3z6x6 = (~(Ej07x6 & Lj07x6));
assign D107x6 = (Sj07x6 ? I4w6x6 : B4w6x6);
assign I4w6x6 = (~(Zj07x6 & Dzu6x6));
assign B4w6x6 = (~(Zj07x6 & Gk07x6));
assign Zj07x6 = (L2w6x6 & Nk07x6);
assign L2w6x6 = (~(Xrbov6 & Dzu6x6));
assign P007x6 = (Sj07x6 | Byu6x6);
assign Sj07x6 = (~(Uk07x6 & Bl07x6));
assign Bl07x6 = (Okx6x6 | Iax6x6);
assign Iax6x6 = (!Kuz6x6);
assign Uk07x6 = (Il07x6 & Jgv6x6);
assign Il07x6 = (~(Ybx6x6 & Qgv6x6));
assign Ybx6x6 = (!Wax6x6);
assign R6ziw6 = (!Zf3ov6);
assign Zf3ov6 = (~(Pl07x6 & Zho6x6));
assign Pl07x6 = (~(Ubo6x6 | Mrbdt6));
assign B007x6 = (~(F7ziw6 & Je3ov6));
assign Je3ov6 = (Wl07x6 ^ Dte7z6[1]);
assign O9u6x6 = (Dm07x6 & Km07x6);
assign Km07x6 = (Rm07x6 & Ym07x6);
assign Ym07x6 = (Fn07x6 & Mn07x6);
assign Mn07x6 = (~(Cqf7z6[14] & Q2ziw6));
assign Q2ziw6 = (~(Tn07x6 & Ao07x6));
assign Ao07x6 = (~(Ho07x6 & Tdtiw6));
assign Ho07x6 = (Gzz6x6 & Nzz6x6);
assign Tn07x6 = (~(Dqtiw6 & Oo07x6));
assign Fn07x6 = (~(L0g7z6[14] & O1ziw6));
assign O1ziw6 = (~(Dqtiw6 | Vo07x6));
assign Rm07x6 = (Cp07x6 & Jp07x6);
assign Jp07x6 = (~(U4ziw6 & V1c7z6[30]));
assign U4ziw6 = (Qp07x6 & Xp07x6);
assign Cp07x6 = (~(B5ziw6 & D6gdt6));
assign B5ziw6 = (Kdo6x6 & Dte7z6[13]);
assign Kdo6x6 = (Eq07x6 & Dte7z6[17]);
assign Eq07x6 = (~(Dte7z6[15] | Dte7z6[16]));
assign Dm07x6 = (Lq07x6 & Sq07x6);
assign Sq07x6 = (Zq07x6 & Gr07x6);
assign Gr07x6 = (~(Z3ziw6 & E3c7z6[1]));
assign Z3ziw6 = (Qp07x6 & Zrz6x6);
assign Zq07x6 = (~(Pvkdt6 & Oztiw6));
assign Lq07x6 = (Kq2ov6 & T7ziw6);
assign T7ziw6 = (Nr07x6 & Ur07x6);
assign Ur07x6 = (~(H8ziw6 & Bs07x6));
assign Bs07x6 = (Is07x6 | Nll6x6);
assign Nll6x6 = (Ps07x6 & Mrbdt6);
assign Ps07x6 = (~(Zho6x6 | F7ziw6));
assign F7ziw6 = (Gg3ov6 & I0c7z6[1]);
assign Is07x6 = (~(Ubo6x6 | Bi2ov6));
assign Bi2ov6 = (!Mrbdt6);
assign H8ziw6 = (Gg3ov6 & Ws07x6);
assign Ws07x6 = (Dte7z6[1] ^ Soo6x6);
assign Soo6x6 = (T3cdt6 ? V1c7z6[7] : Bv3ov6);
assign Bv3ov6 = (Kt07x6 ? Dt07x6 : Xrbov6);
assign Kt07x6 = (~(Dzu6x6 ^ Rt07x6));
assign Rt07x6 = (Eav6x6 & Bgy6x6);
assign Bgy6x6 = (!Yt07x6);
assign Dt07x6 = (~(Fu07x6 & Mu07x6));
assign Mu07x6 = (Tu07x6 & Av07x6);
assign Av07x6 = (M0v6x6 | Pqv6x6);
assign Pqv6x6 = (Hv07x6 & Ov07x6);
assign Ov07x6 = (Vv07x6 & Cw07x6);
assign Cw07x6 = (~(V307x6 & Jw07x6));
assign Vv07x6 = (Lvv6x6 | Tkw6x6);
assign Hv07x6 = (Qw07x6 & Xw07x6);
assign Xw07x6 = (Juv6x6 | Ex07x6);
assign Qw07x6 = (~(Zvv6x6 & Cmw6x6));
assign Cmw6x6 = (~(Lx07x6 & Sx07x6));
assign Tu07x6 = (A1v6x6 | Bxv6x6);
assign Bxv6x6 = (Zx07x6 & Gy07x6);
assign Gy07x6 = (Ny07x6 & Uy07x6);
assign Uy07x6 = (Mkw6x6 | Bz07x6);
assign Ny07x6 = (Lvv6x6 | Asw6x6);
assign Zx07x6 = (Iz07x6 & Pz07x6);
assign Pz07x6 = (~(Vlw6x6 & Wz07x6));
assign Iz07x6 = (~(Zvv6x6 & Ctw6x6));
assign Ctw6x6 = (~(D017x6 & K017x6));
assign Fu07x6 = (R017x6 & Y017x6);
assign Y017x6 = (Q2v6x6 | N3w6x6);
assign N3w6x6 = (F117x6 & M117x6);
assign M117x6 = (T117x6 & A217x6);
assign A217x6 = (Mkw6x6 | Svv6x6);
assign T117x6 = (Lvv6x6 | Vzw6x6);
assign F117x6 = (H217x6 & O217x6);
assign O217x6 = (~(Vlw6x6 & Gwv6x6));
assign Gwv6x6 = (~(V217x6 & C317x6));
assign H217x6 = (~(Zvv6x6 & X0x6x6));
assign X0x6x6 = (~(J317x6 & Q317x6));
assign R017x6 = (C2v6x6 | U3w6x6);
assign U3w6x6 = (X317x6 & E417x6);
assign E417x6 = (L417x6 & S417x6);
assign S417x6 = (Mkw6x6 | Cxz6x6);
assign L417x6 = (Lvv6x6 | J7x6x6);
assign X317x6 = (Z417x6 & G517x6);
assign G517x6 = (~(Vlw6x6 & Jxz6x6));
assign Jxz6x6 = (~(N517x6 & U517x6));
assign Z417x6 = (~(Zvv6x6 & L8x6x6));
assign L8x6x6 = (~(B617x6 & I617x6));
assign Nr07x6 = (~(P617x6 & W617x6));
assign W617x6 = (Ok3ov6 & Ubo6x6);
assign Ubo6x6 = (~(Gg3ov6 & Bqziw6));
assign Ok3ov6 = (~(Pk5jw6 ^ Dte7z6[1]));
assign Pk5jw6 = (T3cdt6 ? S1ohw6 : I24ov6);
assign S1ohw6 = (!V1c7z6[15]);
assign I24ov6 = (!M85jw6);
assign M85jw6 = (~(D717x6 & K717x6));
assign K717x6 = (~(R717x6 & Y717x6));
assign Y717x6 = (~(F817x6 & M817x6));
assign M817x6 = (T817x6 & A917x6);
assign A917x6 = (M0v6x6 | Euw6x6);
assign Euw6x6 = (H917x6 & O917x6);
assign O917x6 = (V917x6 & Ca17x6);
assign Ca17x6 = (Mkw6x6 | Alw6x6);
assign Alw6x6 = (S507x6 & Ja17x6);
assign S507x6 = (Qa17x6 & Xa17x6);
assign Xa17x6 = (~(Cve7z6[16] & We07x6));
assign Qa17x6 = (~(Dbx6x6 & Cve7z6[0]));
assign V917x6 = (Lvv6x6 | P8z6x6);
assign P8z6x6 = (G607x6 & D017x6);
assign D017x6 = (Eb17x6 & Lb17x6);
assign Lb17x6 = (~(Cve7z6[28] & Sb17x6));
assign Eb17x6 = (~(Cve7z6[12] & Kbx6x6));
assign G607x6 = (Zb17x6 & Gc17x6);
assign Gc17x6 = (~(Cve7z6[20] & We07x6));
assign Zb17x6 = (~(Cve7z6[4] & Dbx6x6));
assign H917x6 = (Nc17x6 & Uc17x6);
assign Uc17x6 = (~(Vlw6x6 & Jmw6x6));
assign Jmw6x6 = (~(Bd17x6 & Id17x6));
assign Nc17x6 = (E1x6x6 | R9z6x6);
assign R9z6x6 = (Pd17x6 & R807x6);
assign R807x6 = (Wd17x6 & De17x6);
assign De17x6 = (~(Cve7z6[3] & Sb17x6));
assign Wd17x6 = (~(Cve7z6[19] & Kbx6x6));
assign Pd17x6 = (Ke17x6 & Re17x6);
assign Re17x6 = (~(Cve7z6[11] & We07x6));
assign Ke17x6 = (~(Cve7z6[27] & Dbx6x6));
assign T817x6 = (A1v6x6 | G2x6x6);
assign G2x6x6 = (Ye17x6 & Ff17x6);
assign Ff17x6 = (Mf17x6 & Tf17x6);
assign Tf17x6 = (Mkw6x6 | Hsw6x6);
assign Hsw6x6 = (Qi07x6 & V217x6);
assign V217x6 = (Ag17x6 & Hg17x6);
assign Hg17x6 = (~(Cve7z6[25] & Sb17x6));
assign Ag17x6 = (~(Cve7z6[9] & Kbx6x6));
assign Qi07x6 = (Og17x6 & Vg17x6);
assign Vg17x6 = (~(Cve7z6[17] & We07x6));
assign Og17x6 = (~(Cve7z6[1] & Dbx6x6));
assign Mf17x6 = (Lvv6x6 | Qzx6x6);
assign Qzx6x6 = (Ej07x6 & J317x6);
assign J317x6 = (Ch17x6 & Jh17x6);
assign Jh17x6 = (~(Cve7z6[29] & Sb17x6));
assign Ch17x6 = (~(Cve7z6[13] & Kbx6x6));
assign Ej07x6 = (Qh17x6 & Xh17x6);
assign Xh17x6 = (~(Cve7z6[21] & We07x6));
assign Qh17x6 = (~(Cve7z6[5] & Dbx6x6));
assign Ye17x6 = (Ei17x6 & Li17x6);
assign Li17x6 = (~(Vlw6x6 & Jtw6x6));
assign Jtw6x6 = (~(Si17x6 & Zi17x6));
assign Si17x6 = (Xb07x6 & Ec07x6);
assign Ec07x6 = (~(Cve7z6[16] & Kbx6x6));
assign Xb07x6 = (~(Sb17x6 & Cve7z6[0]));
assign Ei17x6 = (E1x6x6 | Z0y6x6);
assign Z0y6x6 = (Gj17x6 & Sc07x6);
assign Sc07x6 = (Nj17x6 & Uj17x6);
assign Uj17x6 = (~(Cve7z6[4] & Sb17x6));
assign Nj17x6 = (~(Cve7z6[20] & Kbx6x6));
assign Gj17x6 = (Bk17x6 & Ik17x6);
assign Ik17x6 = (~(Cve7z6[12] & We07x6));
assign Bk17x6 = (~(Cve7z6[28] & Dbx6x6));
assign F817x6 = (Pk17x6 & Wk17x6);
assign Wk17x6 = (Q2v6x6 | N9x6x6);
assign N9x6x6 = (Dl17x6 & Kl17x6);
assign Kl17x6 = (Rl17x6 & Yl17x6);
assign Yl17x6 = (Mkw6x6 | C0x6x6);
assign C0x6x6 = (Aa07x6 & N517x6);
assign N517x6 = (Fm17x6 & Mm17x6);
assign Mm17x6 = (~(Cve7z6[26] & Sb17x6));
assign Fm17x6 = (~(Cve7z6[10] & Kbx6x6));
assign Aa07x6 = (Tm17x6 & An17x6);
assign An17x6 = (~(Cve7z6[18] & We07x6));
assign Tm17x6 = (~(Cve7z6[2] & Dbx6x6));
assign Rl17x6 = (Lvv6x6 | E7y6x6);
assign E7y6x6 = (B617x6 & Hn17x6);
assign B617x6 = (On17x6 & Vn17x6);
assign Vn17x6 = (~(Cve7z6[30] & Sb17x6));
assign On17x6 = (~(Cve7z6[14] & Kbx6x6));
assign Dl17x6 = (Co17x6 & Jo17x6);
assign Jo17x6 = (Juv6x6 | L1x6x6);
assign L1x6x6 = (Qo17x6 & C407x6);
assign C407x6 = (Xo17x6 & Ep17x6);
assign Ep17x6 = (~(Cve7z6[1] & Sb17x6));
assign Xo17x6 = (~(Cve7z6[17] & Kbx6x6));
assign Qo17x6 = (Lp17x6 & Sp17x6);
assign Sp17x6 = (~(Cve7z6[9] & We07x6));
assign Lp17x6 = (~(Cve7z6[25] & Dbx6x6));
assign Co17x6 = (E1x6x6 | G8y6x6);
assign G8y6x6 = (Zp17x6 & Q407x6);
assign Q407x6 = (Gq17x6 & Nq17x6);
assign Nq17x6 = (~(Cve7z6[5] & Sb17x6));
assign Gq17x6 = (~(Cve7z6[21] & Kbx6x6));
assign Zp17x6 = (Uq17x6 & Br17x6);
assign Br17x6 = (~(Cve7z6[13] & We07x6));
assign Uq17x6 = (~(Cve7z6[29] & Dbx6x6));
assign Pk17x6 = (C2v6x6 | Yix6x6);
assign Yix6x6 = (Ir17x6 & Pr17x6);
assign Pr17x6 = (Wr17x6 & Ds17x6);
assign Ds17x6 = (Mkw6x6 | Q7x6x6);
assign Q7x6x6 = (Df07x6 & Lx07x6);
assign Lx07x6 = (Ks17x6 & Rs17x6);
assign Rs17x6 = (~(Cve7z6[27] & Sb17x6));
assign Ks17x6 = (~(Cve7z6[11] & Kbx6x6));
assign Df07x6 = (Ys17x6 & Ft17x6);
assign Ft17x6 = (~(Cve7z6[19] & We07x6));
assign Ys17x6 = (~(Cve7z6[3] & Dbx6x6));
assign Wr17x6 = (Lvv6x6 | K807x6);
assign K807x6 = (Bd17x6 & Mt17x6);
assign Bd17x6 = (Tt17x6 & Au17x6);
assign Au17x6 = (~(Sb17x6 & Neo7v6));
assign Tt17x6 = (~(Cve7z6[15] & Kbx6x6));
assign Ir17x6 = (Hu17x6 & Ou17x6);
assign Ou17x6 = (Juv6x6 | S8x6x6);
assign S8x6x6 = (Vu17x6 & Ah07x6);
assign Ah07x6 = (Cv17x6 & Jv17x6);
assign Jv17x6 = (~(Cve7z6[2] & Sb17x6));
assign Cv17x6 = (~(Cve7z6[18] & Kbx6x6));
assign Vu17x6 = (Qv17x6 & Xv17x6);
assign Xv17x6 = (~(Cve7z6[10] & We07x6));
assign Qv17x6 = (~(Cve7z6[26] & Dbx6x6));
assign Hu17x6 = (E1x6x6 | T907x6);
assign T907x6 = (Ew17x6 & Oh07x6);
assign Oh07x6 = (Lw17x6 & Sw17x6);
assign Sw17x6 = (~(Cve7z6[6] & Sb17x6));
assign Lw17x6 = (~(Cve7z6[22] & Kbx6x6));
assign Ew17x6 = (Zw17x6 & Gx17x6);
assign Gx17x6 = (~(Cve7z6[14] & We07x6));
assign Zw17x6 = (~(Cve7z6[30] & Dbx6x6));
assign R717x6 = (~(Dzu6x6 ^ Nx17x6));
assign D717x6 = (~(Xrbov6 & Ux17x6));
assign Ux17x6 = (Dzu6x6 | Nx17x6);
assign Nx17x6 = (By17x6 & Iy17x6);
assign Iy17x6 = (Wax6x6 & Okx6x6);
assign Wax6x6 = (Py17x6 | Dbx6x6);
assign By17x6 = (Nfy6x6 & Wy17x6);
assign Wy17x6 = (~(Sb17x6 & Yt07x6));
assign Nfy6x6 = (Vfv6x6 & Jgv6x6);
assign Jgv6x6 = (!Ajy6x6);
assign P617x6 = (Zho6x6 & Mrbdt6);
assign Zho6x6 = (Gg3ov6 & I0c7z6[0]);
assign Gg3ov6 = (Qp07x6 & Dz17x6);
assign Dz17x6 = (~(Bdu6x6 & Kz17x6));
assign Kq2ov6 = (Iymnv6 ? Yz17x6 : Rz17x6);
assign Iymnv6 = (F027x6 ^ Mennv6);
assign Mennv6 = (M027x6 & T027x6);
assign T027x6 = (A127x6 & Nu8jw6);
assign Nu8jw6 = (!Dte7z6[1]);
assign M027x6 = (H127x6 & O127x6);
assign O127x6 = (~(V127x6 & Nvtiw6));
assign V127x6 = (Gzz6x6 & Zrz6x6);
assign Gzz6x6 = (C227x6 & Dte7z6[15]);
assign C227x6 = (~(J227x6 | Djgdt6));
assign H127x6 = (Kxb7z6[31] ? X227x6 : Q227x6);
assign X227x6 = (~(E327x6 & L327x6));
assign L327x6 = (~(Z6jhw6 & S327x6));
assign S327x6 = (~(Z327x6 & G427x6));
assign Z327x6 = (Bdf7z6[3] & Nh2ov6);
assign Q227x6 = (~(N427x6 & Gvtiw6));
assign F027x6 = (~(U427x6 & B527x6));
assign B527x6 = (I527x6 & P527x6);
assign P527x6 = (W527x6 & D627x6);
assign D627x6 = (~(Su0jw6 & Yxf7z6[32]));
assign Su0jw6 = (K627x6 & Ijziw6);
assign Ijziw6 = (Pne7z6[1] & R627x6);
assign W527x6 = (Y627x6 & F727x6);
assign F727x6 = (~(Yxf7z6[30] & Nv0jw6));
assign Nv0jw6 = (K627x6 & Giziw6);
assign Giziw6 = (~(Pne7z6[0] | Pne7z6[1]));
assign Y627x6 = (~(Uv0jw6 & Yxf7z6[31]));
assign Uv0jw6 = (K627x6 & Niziw6);
assign Niziw6 = (~(R627x6 | Pne7z6[1]));
assign R627x6 = (!Pne7z6[0]);
assign I527x6 = (M727x6 & T727x6);
assign T727x6 = (~(Pw0jw6 & Yxf7z6[33]));
assign Pw0jw6 = (K627x6 & Pjziw6);
assign Pjziw6 = (Pne7z6[1] & Pne7z6[0]);
assign K627x6 = (Gvtiw6 & Ydziw6);
assign Gvtiw6 = (A827x6 & Bdf7z6[3]);
assign M727x6 = (~(Hz0jw6 & Kxb7z6[30]));
assign Hz0jw6 = (~(Z6jhw6 | H827x6));
assign U427x6 = (O827x6 & V827x6);
assign V827x6 = (C927x6 & J927x6);
assign J927x6 = (~(Alf7z6[14] & J01jw6));
assign J01jw6 = (Ydziw6 & Rkziw6);
assign Rkziw6 = (~(Q927x6 & X927x6));
assign Q927x6 = (Pbtiw6 & E4lhw6);
assign C927x6 = (Ea27x6 & La27x6);
assign La27x6 = (~(Oz0jw6 & Fhc7z6[30]));
assign Oz0jw6 = (Sa27x6 & Za27x6);
assign Sa27x6 = (Ydziw6 & Kxb7z6[31]);
assign Ea27x6 = (~(Onf7z6[30] & My0jw6));
assign My0jw6 = (Ydziw6 & Ofziw6);
assign O827x6 = (Gb27x6 & Nb27x6);
assign Nb27x6 = (~(Wl07x6 & Rdziw6));
assign Rdziw6 = (!Dx0jw6);
assign Wl07x6 = (T3cdt6 ? V1c7z6[30] : Iv3ov6);
assign Iv3ov6 = (Bc27x6 ? Xrbov6 : Ub27x6);
assign Bc27x6 = (Pyu6x6 & Ic27x6);
assign Ic27x6 = (~(Pc27x6 & Ajy6x6));
assign Pc27x6 = (Sov6x6 & Kuz6x6);
assign Sov6x6 = (!Dzu6x6);
assign Pyu6x6 = (Nk07x6 & Gk07x6);
assign Gk07x6 = (~(Vfv6x6 & Dzu6x6));
assign Nk07x6 = (Dzu6x6 | Vfv6x6);
assign Ub27x6 = (~(Wc27x6 & Dd27x6));
assign Dd27x6 = (Kd27x6 & Rd27x6);
assign Rd27x6 = (M0v6x6 | Yoy6x6);
assign Yoy6x6 = (Yd27x6 & Fe27x6);
assign Fe27x6 = (Me27x6 & Te27x6);
assign Te27x6 = (Mkw6x6 | Dnz6x6);
assign Dnz6x6 = (Be07x6 & Af27x6);
assign Be07x6 = (Hf27x6 & Of27x6);
assign Of27x6 = (~(Cve7z6[7] & Sb17x6));
assign Hf27x6 = (~(Cve7z6[23] & Kbx6x6));
assign Me27x6 = (Lvv6x6 | Vf27x6);
assign Yd27x6 = (Cg27x6 & Jg27x6);
assign Jg27x6 = (Juv6x6 | Foz6x6);
assign Foz6x6 = (Qg27x6 & Xg27x6);
assign Qg27x6 = (Hn17x6 & Eh27x6);
assign Eh27x6 = (~(Cve7z6[22] & We07x6));
assign Hn17x6 = (~(Cve7z6[6] & Dbx6x6));
assign Cg27x6 = (E1x6x6 | Lh27x6);
assign Kd27x6 = (A1v6x6 | T0v6x6);
assign T0v6x6 = (Sh27x6 & Zh27x6);
assign Zh27x6 = (Gi27x6 & Ni27x6);
assign Ni27x6 = (Mkw6x6 | Vpz6x6);
assign Vpz6x6 = (Ui27x6 & Z507x6);
assign Z507x6 = (Bj27x6 & Ij27x6);
assign Ij27x6 = (~(Cve7z6[8] & Sb17x6));
assign Bj27x6 = (~(Cve7z6[24] & Kbx6x6));
assign Gi27x6 = (Lvv6x6 | Pj27x6);
assign Sh27x6 = (Wj27x6 & Dk27x6);
assign Dk27x6 = (E1x6x6 | Kk27x6);
assign Wj27x6 = (Juv6x6 | Xqz6x6);
assign Xqz6x6 = (Rk27x6 & Yk27x6);
assign Rk27x6 = (Mt17x6 & Fl27x6);
assign Fl27x6 = (~(Cve7z6[23] & We07x6));
assign Mt17x6 = (~(Cve7z6[7] & Dbx6x6));
assign Wc27x6 = (Ml27x6 & Tl27x6);
assign Tl27x6 = (Q2v6x6 | H1v6x6);
assign H1v6x6 = (Am27x6 & Hm27x6);
assign Hm27x6 = (Om27x6 & Vm27x6);
assign Vm27x6 = (Mkw6x6 | G0z6x6);
assign G0z6x6 = (C317x6 & Xi07x6);
assign Xi07x6 = (Cn27x6 & Jn27x6);
assign Jn27x6 = (~(Cve7z6[9] & Sb17x6));
assign Cn27x6 = (~(Cve7z6[25] & Kbx6x6));
assign C317x6 = (Qn27x6 & Xn27x6);
assign Xn27x6 = (~(Cve7z6[1] & We07x6));
assign Qn27x6 = (~(Cve7z6[17] & Dbx6x6));
assign Om27x6 = (~(Xzx6x6 & Eo27x6));
assign Eo27x6 = (~(Q317x6 & Lj07x6));
assign Lj07x6 = (Lo27x6 & So27x6);
assign So27x6 = (~(Cve7z6[13] & Sb17x6));
assign Lo27x6 = (~(Cve7z6[29] & Kbx6x6));
assign Q317x6 = (Zo27x6 & Gp27x6);
assign Gp27x6 = (~(Cve7z6[5] & We07x6));
assign Zo27x6 = (~(Cve7z6[21] & Dbx6x6));
assign Am27x6 = (Np27x6 & Up27x6);
assign Up27x6 = (~(Zvv6x6 & Bq27x6));
assign Np27x6 = (Juv6x6 | I1z6x6);
assign I1z6x6 = (Iq27x6 & Pq27x6);
assign Iq27x6 = (Wq27x6 & Lc07x6);
assign Lc07x6 = (~(Cve7z6[8] & Dbx6x6));
assign Wq27x6 = (~(Cve7z6[24] & We07x6));
assign Ml27x6 = (C2v6x6 | X2v6x6);
assign Gb27x6 = (~(Alf7z6[30] & Q01jw6));
assign Q01jw6 = (~(H827x6 | Kkziw6));
assign Kkziw6 = (~(Frtiw6 | Wcnnv6));
assign Wcnnv6 = (!Uvtiw6);
assign Yz17x6 = (~(Bymnv6 & Ubziw6));
assign Ubziw6 = (!Bcziw6);
assign Rz17x6 = (Bymnv6 ? Icziw6 : Bcziw6);
assign Bymnv6 = (Dr27x6 ^ Dte7z6[0]);
assign Dr27x6 = (~(Kr27x6 & Rr27x6));
assign Rr27x6 = (~(Yxf7z6[14] & Laziw6));
assign Laziw6 = (~(H827x6 | T8riw6));
assign T8riw6 = (E4lhw6 & Mdtiw6);
assign Mdtiw6 = (!Dqtiw6);
assign Kr27x6 = (Yr27x6 & Fs27x6);
assign Fs27x6 = (~(Yxf7z6[30] & Gbziw6));
assign Gbziw6 = (Ydziw6 & Ms27x6);
assign Ms27x6 = (~(Ts27x6 & A127x6));
assign Yr27x6 = (~(Kxb7z6[30] & Nbziw6));
assign Nbziw6 = (~(Dx0jw6 & Zs2jw6));
assign Zs2jw6 = (H827x6 | At27x6);
assign At27x6 = (~(Ht27x6 | Ofziw6));
assign Ofziw6 = (~(Ot27x6 & Cmtiw6));
assign Ht27x6 = (~(Uvtiw6 & Qgziw6));
assign Qgziw6 = (~(Za27x6 & Fhc7z6[31]));
assign Za27x6 = (Vt27x6 & Hetiw6);
assign Vt27x6 = (Mrbdt6 & Cu27x6);
assign Uvtiw6 = (~(A827x6 & Ju27x6));
assign Dx0jw6 = (~(Fennv6 | Jm2ov6));
assign Jm2ov6 = (!Gw1ov6);
assign Gw1ov6 = (~(Dte7z6[3] & Qu27x6));
assign Qu27x6 = (~(Qp07x6 & J1gov6));
assign Fennv6 = (Xu27x6 & Bdu6x6);
assign Icziw6 = (Ev27x6 & Lv27x6);
assign Ev27x6 = (~(Zrz6x6 & Xu27x6));
assign Bcziw6 = (Sv27x6 & Lv27x6);
assign Lv27x6 = (~(Xu27x6 & Bqziw6));
assign Sv27x6 = (~(Xu27x6 & Xp07x6));
assign Gv9ov6 = (~(Zv27x6 | T1u6x6));
assign T1u6x6 = (~(Gw27x6 & Nw27x6));
assign Nw27x6 = (Uw27x6 & Bx27x6);
assign Bx27x6 = (Ylyiw6 ^ Ix27x6);
assign Ylyiw6 = (Px27x6 | D0u6x6);
assign Px27x6 = (~(Wx27x6 & Spyiw6));
assign Wx27x6 = (~(Dy27x6 & Ky27x6));
assign Ky27x6 = (Yy27x6 ? Ry27x6 : Qij7z6[1]);
assign Ry27x6 = (~(Fz27x6 & Mz27x6));
assign Fz27x6 = (~(M5e7z6[0] & Ldo7v6));
assign Dy27x6 = (Gt2jw6 & Tz27x6);
assign Tz27x6 = (~(A037x6 & M5e7z6[0]));
assign A037x6 = (~(F02nv6 | M5e7z6[1]));
assign Gt2jw6 = (H037x6 & O037x6);
assign Uw27x6 = (Liyiw6 & V037x6);
assign V037x6 = (Xgfhw6 ^ Bkyiw6);
assign Bkyiw6 = (!Siyiw6);
assign Liyiw6 = (Wzt6x6 & C137x6);
assign C137x6 = (~(J137x6 & H037x6));
assign H037x6 = (Q137x6 & X137x6);
assign Q137x6 = (~(E237x6 & L237x6));
assign E237x6 = (~(Gfihw6 | S237x6));
assign J137x6 = (Siyiw6 & D0u6x6);
assign D0u6x6 = (~(Z237x6 & G337x6));
assign Z237x6 = (N337x6 & U337x6);
assign U337x6 = (~(Vuyiw6 & B437x6));
assign N337x6 = (~(Ouyiw6 & X0oov6));
assign Siyiw6 = (O037x6 & Spyiw6);
assign O037x6 = (~(I437x6 & P437x6));
assign I437x6 = (W437x6 & D537x6);
assign D537x6 = (~(K537x6 & Vuyiw6));
assign W437x6 = (~(Ouyiw6 & R537x6));
assign Wzt6x6 = (~(Y537x6 & L237x6));
assign Y537x6 = (Z11jw6 & F637x6);
assign F637x6 = (!Vuyiw6);
assign Z11jw6 = (~(M637x6 & T637x6));
assign T637x6 = (Srknv6 | Gp1ov6);
assign Gp1ov6 = (A737x6 & H737x6);
assign A737x6 = (Dtadt6 & O737x6);
assign O737x6 = (!Kxb7z6[2]);
assign Gw27x6 = (V737x6 & C837x6);
assign C837x6 = (Mlziw6 ^ Uifhw6);
assign Mlziw6 = (!Ziyiw6);
assign Ziyiw6 = (~(J837x6 & Q837x6));
assign Q837x6 = (~(S237x6 | Gninv6));
assign S237x6 = (Vuyiw6 & X837x6);
assign J837x6 = (~(Ouyiw6 | Gfihw6));
assign V737x6 = (Coyiw6 ^ Bjfhw6);
assign Coyiw6 = (!Fmyiw6);
assign Fmyiw6 = (X137x6 | Gninv6);
assign Gninv6 = (!Spyiw6);
assign Spyiw6 = (~(K7e7z6[0] & Pxfov6));
assign X137x6 = (~(E937x6 & L237x6));
assign L237x6 = (!Ouyiw6);
assign E937x6 = (L937x6 & S937x6);
assign S937x6 = (~(Vuyiw6 & Z937x6));
assign Zv27x6 = (Pw9ov6 | R0u6x6);
assign Pw9ov6 = (!Y0u6x6);
assign Y0u6x6 = (~(Ga37x6 & Na37x6));
assign Na37x6 = (Ua37x6 & Bb37x6);
assign Bb37x6 = (Ypinv6 | Ib37x6);
assign Ua37x6 = (Pb37x6 & Wb37x6);
assign Pb37x6 = (~(Etq6x6 & Dc37x6));
assign Dc37x6 = (~(Kc37x6 & Rc37x6));
assign Rc37x6 = (Yc37x6 & Fd37x6);
assign Fd37x6 = (Md37x6 & Td37x6);
assign Td37x6 = (Bnviw6 & T6onv6);
assign Bnviw6 = (Dssov6 & Vnlhw6);
assign Yc37x6 = (Ae37x6 & He37x6);
assign He37x6 = (B5siw6 & Epsov6);
assign Ae37x6 = (Oe37x6 & I4ghw6);
assign Kc37x6 = (Ve37x6 & Cf37x6);
assign Cf37x6 = (Jf37x6 & Qf37x6);
assign Qf37x6 = (Ydsiw6 & Hulhw6);
assign Jf37x6 = (~(Zwlhw6 | Nxlhw6));
assign Zwlhw6 = (~(Bvohw6 & Hcviw6));
assign Bvohw6 = (Ddsiw6 & G3ghw6);
assign Ve37x6 = (Xf37x6 & Eg37x6);
assign Eg37x6 = (Bylhw6 & Iylhw6);
assign Iylhw6 = (Lg37x6 & Sg37x6);
assign Sg37x6 = (Iyriw6 & Nqehw6);
assign Iyriw6 = (Yzehw6 & T1riw6);
assign Lg37x6 = (Gqehw6 & Mefhw6);
assign Xf37x6 = (Liriw6 & Wrsov6);
assign Wrsov6 = (L4riw6 & D0riw6);
assign Liriw6 = (Vcviw6 & Zg37x6);
assign Zg37x6 = (~(Gh37x6 | Nh37x6));
assign Vcviw6 = (Rlriw6 & Uh37x6);
assign Etq6x6 = (~(Hs9ov6 & Bsrov6));
assign Hs9ov6 = (!Snvnv6);
assign Ga37x6 = (Bi37x6 & Ii37x6);
assign Ii37x6 = (~(Gr2et6 & Pi37x6));
assign Pi37x6 = (~(Wi37x6 & Dj37x6));
assign Tly7v6 = (Kj37x6 & Qf2ov6);
assign Kj37x6 = (~(Gepiw6 | Lg2ov6));
assign Gepiw6 = (~(Gh2ov6 & Fhc7z6[31]));
assign Gh2ov6 = (Rj37x6 & Yj37x6);
assign Yj37x6 = (Fk37x6 & Mk37x6);
assign Mk37x6 = (Tk37x6 & Al37x6);
assign Al37x6 = (~(Hl37x6 | Kxb7z6[28]));
assign Hl37x6 = (Kxb7z6[29] | Kxb7z6[30]);
assign Fk37x6 = (Ol37x6 & Vl37x6);
assign Rj37x6 = (Cm37x6 & Jm37x6);
assign Jm37x6 = (Qm37x6 & Xm37x6);
assign Xm37x6 = (~(En37x6 | Kxb7z6[19]));
assign En37x6 = (Kxb7z6[20] | Kxb7z6[21]);
assign Qm37x6 = (~(Kxb7z6[17] | Kxb7z6[18]));
assign Cm37x6 = (Ln37x6 & Sn37x6);
assign Sn37x6 = (~(Zn37x6 | Kxb7z6[16]));
assign Ln37x6 = (Go37x6 & E327x6);
assign Mly7v6 = (Lg2ov6 ? Elgdt6 : N427x6);
assign Lg2ov6 = (No37x6 & Uo37x6);
assign Uo37x6 = (~(Qf2ov6 & Qg2nv6));
assign No37x6 = (~(Fre7z6[0] | Fre7z6[1]));
assign Fly7v6 = (~(Bp37x6 & Ip37x6));
assign Ip37x6 = (~(Vi7et6 & Vrinv6));
assign Bp37x6 = (~(Pp37x6 & Wp37x6));
assign Pp37x6 = (Dq37x6 & Kq37x6);
assign Kq37x6 = (Ii9ov6 ? Yq37x6 : Rq37x6);
assign Yq37x6 = (Fr37x6 & Bi9ov6);
assign Fr37x6 = (Xvehw6 ? Tr37x6 : Mr37x6);
assign Tr37x6 = (As37x6 & Hs37x6);
assign Hs37x6 = (Os37x6 & Vs37x6);
assign Vs37x6 = (~(Lvg7z6[2] ^ S4lhw6));
assign Os37x6 = (~(Lvg7z6[1] ^ Xehov6));
assign As37x6 = (Ct37x6 & Jt37x6);
assign Jt37x6 = (~(Lvg7z6[0] ^ I6lhw6));
assign Ct37x6 = (~(Lvg7z6[3] ^ L4lhw6));
assign Mr37x6 = (Qt37x6 & Xt37x6);
assign Xt37x6 = (Eu37x6 & Lu37x6);
assign Lu37x6 = (~(Lvg7z6[3] ^ Nfihw6));
assign Eu37x6 = (~(Lvg7z6[2] ^ Xdihw6));
assign Qt37x6 = (Su37x6 & Zu37x6);
assign Zu37x6 = (Lvg7z6[0] ^ Mjq6x6);
assign Su37x6 = (Lvg7z6[1] ^ Ypq6x6);
assign Ypq6x6 = (!F4ihw6);
assign Rq37x6 = (Xvehw6 ? Nv37x6 : Gv37x6);
assign Nv37x6 = (Uv37x6 & Bw37x6);
assign Bw37x6 = (Iw37x6 & Pw37x6);
assign Pw37x6 = (Yelhw6 ^ S4lhw6);
assign S4lhw6 = (~(Ww37x6 & Dx37x6));
assign Dx37x6 = (Kx37x6 & Rx37x6);
assign Rx37x6 = (~(Zec7z6[30] & Yx37x6));
assign Kx37x6 = (Jlohw6 | Fy37x6);
assign Ww37x6 = (My37x6 & Ty37x6);
assign Iw37x6 = (~(Ntg7z6[1] ^ Xehov6));
assign Xehov6 = (~(Az37x6 & Hz37x6));
assign Hz37x6 = (Oz37x6 & Vz37x6);
assign Vz37x6 = (Buihw6 | Fy37x6);
assign Oz37x6 = (~(Yx37x6 & M6nhw6));
assign Az37x6 = (C047x6 & Jvlhw6);
assign Uv37x6 = (J047x6 & Q047x6);
assign Q047x6 = (~(Ntg7z6[0] ^ I6lhw6));
assign I6lhw6 = (~(X047x6 & E147x6));
assign E147x6 = (L147x6 & S147x6);
assign S147x6 = (~(Yx37x6 & Z9nhw6));
assign L147x6 = (Lofhw6 | Fy37x6);
assign X047x6 = (Z147x6 & Ty37x6);
assign J047x6 = (Oglhw6 ^ L4lhw6);
assign L4lhw6 = (~(G247x6 & N247x6));
assign N247x6 = (U247x6 & B347x6);
assign B347x6 = (Offhw6 | Fy37x6);
assign Fy37x6 = (I347x6 & P347x6);
assign P347x6 = (W347x6 & Onlhw6);
assign I347x6 = (D447x6 & Mquiw6);
assign U247x6 = (K447x6 & R447x6);
assign K447x6 = (~(Zec7z6[31] & Yx37x6));
assign Yx37x6 = (~(Y447x6 & F547x6));
assign G247x6 = (M547x6 & Ty37x6);
assign Ty37x6 = (Jvlhw6 & Hffhw6);
assign Gv37x6 = (T547x6 & A647x6);
assign A647x6 = (H647x6 & O647x6);
assign O647x6 = (Oglhw6 ^ Nfihw6);
assign H647x6 = (Yelhw6 ^ Xdihw6);
assign T547x6 = (V647x6 & C747x6);
assign C747x6 = (Gclhw6 ^ Zeihw6);
assign V647x6 = (Pdlhw6 ^ F4ihw6);
assign Dq37x6 = (Ypinv6 ? Atmov6 : Fsmov6);
assign Yky7v6 = (~(J747x6 & Q747x6));
assign Q747x6 = (X747x6 & E847x6);
assign E847x6 = (~(Ivwnv6 & E3c7z6[0]));
assign X747x6 = (L847x6 & S847x6);
assign S847x6 = (Z847x6 | G21jw6);
assign G21jw6 = (G947x6 & N947x6);
assign N947x6 = (U947x6 & Ba47x6);
assign Ba47x6 = (Ia47x6 & Pa47x6);
assign Pa47x6 = (~(Wa47x6 & Db47x6));
assign Db47x6 = (Kb47x6 & Ijmov6);
assign Wa47x6 = (R3h7z6[0] & Rb47x6);
assign Rb47x6 = (~(Yb47x6 & Fc47x6));
assign Fc47x6 = (~(EXRESPD & Mc47x6));
assign Yb47x6 = (~(Tc47x6 | R3h7z6[1]));
assign Tc47x6 = (EXRESPS & Ad47x6);
assign Ia47x6 = (~(Swlov6 & Rsyiw6));
assign U947x6 = (Hd47x6 & Od47x6);
assign Od47x6 = (~(Nqh7z6[0] & Ysyiw6));
assign Hd47x6 = (Vd47x6 | R3ihw6);
assign G947x6 = (Ce47x6 & Je47x6);
assign Ce47x6 = (Qe47x6 & Xe47x6);
assign Xe47x6 = (~(Fth7z6[0] & Ttyiw6));
assign Qe47x6 = (~(Uyb7z6[0] & Ef47x6));
assign L847x6 = (~(Lf47x6 & Sf47x6));
assign Sf47x6 = (~(Zf47x6 & Gg47x6));
assign Gg47x6 = (Ng47x6 & Ug47x6);
assign Ug47x6 = (~(Bh47x6 & Ve9ov6));
assign Ng47x6 = (Ih47x6 & Ph47x6);
assign Ph47x6 = (~(Wh47x6 & Zfhov6));
assign Ih47x6 = (~(Di47x6 & Et9iw6));
assign Zf47x6 = (Ki47x6 & Ri47x6);
assign Ri47x6 = (~(Yi47x6 & Td9ov6));
assign Ki47x6 = (Fj47x6 & Mj47x6);
assign Mj47x6 = (~(Tj47x6 & Jf9ov6));
assign Fj47x6 = (~(Ak47x6 & Fd9ov6));
assign J747x6 = (Hk47x6 & Ok47x6);
assign Ok47x6 = (~(Kwwnv6 & Fth7z6[0]));
assign Hk47x6 = (Vk47x6 & Cl47x6);
assign Cl47x6 = (~(Ztwnv6 & Kxb7z6[0]));
assign Vk47x6 = (~(Nqh7z6[0] & Dwwnv6));
assign Rky7v6 = (~(Jl47x6 & Ql47x6));
assign Ql47x6 = (Xl47x6 & Em47x6);
assign Em47x6 = (~(Ztwnv6 & Kxb7z6[30]));
assign Xl47x6 = (Lm47x6 & Sm47x6);
assign Sm47x6 = (~(Uuwnv6 & Acxnv6));
assign Acxnv6 = (~(Zm47x6 & Gn47x6));
assign Gn47x6 = (Nn47x6 & Un47x6);
assign Un47x6 = (~(Wryiw6 & Xkjnv6));
assign Nn47x6 = (Bo47x6 & Io47x6);
assign Io47x6 = (~(Tk2ov6 & Rsyiw6));
assign Bo47x6 = (~(Nqh7z6[30] & Ysyiw6));
assign Zm47x6 = (Ftyiw6 & Po47x6);
assign Po47x6 = (~(Fth7z6[30] & Ttyiw6));
assign Lm47x6 = (~(Ivwnv6 & Fhc7z6[30]));
assign Jl47x6 = (Wo47x6 & Dp47x6);
assign Dp47x6 = (~(Dwwnv6 & Nqh7z6[30]));
assign Wo47x6 = (~(Kwwnv6 & Fth7z6[30]));
assign Kky7v6 = (~(Kp47x6 & Rp47x6));
assign Rp47x6 = (Yp47x6 & Fq47x6);
assign Fq47x6 = (~(Ztwnv6 & Kxb7z6[29]));
assign Yp47x6 = (Mq47x6 & Tq47x6);
assign Tq47x6 = (~(Uuwnv6 & Pgxnv6));
assign Pgxnv6 = (~(Ar47x6 & Hr47x6));
assign Hr47x6 = (Or47x6 & Vr47x6);
assign Vr47x6 = (~(Wryiw6 & Dojnv6));
assign Or47x6 = (Cs47x6 & Js47x6);
assign Js47x6 = (~(Bnbov6 & Rsyiw6));
assign Cs47x6 = (~(Nqh7z6[29] & Ysyiw6));
assign Ar47x6 = (Ftyiw6 & Qs47x6);
assign Qs47x6 = (~(Fth7z6[29] & Ttyiw6));
assign Mq47x6 = (~(Ivwnv6 & Fhc7z6[29]));
assign Kp47x6 = (Xs47x6 & Et47x6);
assign Et47x6 = (~(Dwwnv6 & Nqh7z6[29]));
assign Xs47x6 = (~(Kwwnv6 & Fth7z6[29]));
assign Dky7v6 = (~(Lt47x6 & St47x6));
assign St47x6 = (Zt47x6 & Gu47x6);
assign Gu47x6 = (~(Ztwnv6 & Kxb7z6[28]));
assign Zt47x6 = (Nu47x6 & Uu47x6);
assign Uu47x6 = (~(Uuwnv6 & Elxnv6));
assign Elxnv6 = (~(Bv47x6 & Iv47x6));
assign Iv47x6 = (Pv47x6 & Wv47x6);
assign Wv47x6 = (~(Wryiw6 & Tpjnv6));
assign Pv47x6 = (Dw47x6 & Kw47x6);
assign Kw47x6 = (~(My9ov6 & Rsyiw6));
assign Dw47x6 = (~(Nqh7z6[28] & Ysyiw6));
assign Bv47x6 = (Ftyiw6 & Rw47x6);
assign Rw47x6 = (~(Fth7z6[28] & Ttyiw6));
assign Nu47x6 = (~(Ivwnv6 & Fhc7z6[28]));
assign Lt47x6 = (Yw47x6 & Fx47x6);
assign Fx47x6 = (~(Dwwnv6 & Nqh7z6[28]));
assign Yw47x6 = (~(Kwwnv6 & Fth7z6[28]));
assign Wjy7v6 = (~(Mx47x6 & Tx47x6));
assign Tx47x6 = (Ay47x6 & Hy47x6);
assign Hy47x6 = (~(Ztwnv6 & Kxb7z6[27]));
assign Ay47x6 = (Oy47x6 & Vy47x6);
assign Vy47x6 = (~(Uuwnv6 & Tpxnv6));
assign Tpxnv6 = (~(Cz47x6 & Jz47x6));
assign Jz47x6 = (Qz47x6 & Xz47x6);
assign Xz47x6 = (~(Wryiw6 & Jrjnv6));
assign Qz47x6 = (E057x6 & L057x6);
assign L057x6 = (~(Htfov6 & Rsyiw6));
assign E057x6 = (~(Nqh7z6[27] & Ysyiw6));
assign Cz47x6 = (Ftyiw6 & S057x6);
assign S057x6 = (~(Fth7z6[27] & Ttyiw6));
assign Oy47x6 = (~(Ivwnv6 & Fhc7z6[27]));
assign Mx47x6 = (Z057x6 & G157x6);
assign G157x6 = (~(Dwwnv6 & Nqh7z6[27]));
assign Z057x6 = (~(Kwwnv6 & Fth7z6[27]));
assign Pjy7v6 = (~(N157x6 & U157x6));
assign U157x6 = (B257x6 & I257x6);
assign I257x6 = (~(Ztwnv6 & Kxb7z6[26]));
assign B257x6 = (P257x6 & W257x6);
assign W257x6 = (~(Uuwnv6 & Iuxnv6));
assign Iuxnv6 = (~(D357x6 & K357x6));
assign K357x6 = (R357x6 & Y357x6);
assign Y357x6 = (~(Wryiw6 & Zsjnv6));
assign R357x6 = (F457x6 & M457x6);
assign M457x6 = (~(Q2mov6 & Rsyiw6));
assign F457x6 = (~(Nqh7z6[26] & Ysyiw6));
assign D357x6 = (Ftyiw6 & T457x6);
assign T457x6 = (~(Fth7z6[26] & Ttyiw6));
assign P257x6 = (~(Ivwnv6 & Fhc7z6[26]));
assign N157x6 = (A557x6 & H557x6);
assign H557x6 = (~(Dwwnv6 & Nqh7z6[26]));
assign A557x6 = (~(Kwwnv6 & Fth7z6[26]));
assign Ijy7v6 = (~(O557x6 & V557x6));
assign V557x6 = (C657x6 & J657x6);
assign J657x6 = (~(Ztwnv6 & Kxb7z6[25]));
assign C657x6 = (Q657x6 & X657x6);
assign X657x6 = (~(Uuwnv6 & Xyxnv6));
assign Xyxnv6 = (~(E757x6 & L757x6));
assign L757x6 = (S757x6 & Z757x6);
assign Z757x6 = (~(Od9iw6 & Rsyiw6));
assign S757x6 = (G857x6 & N857x6);
assign N857x6 = (~(Nqh7z6[25] & Ysyiw6));
assign G857x6 = (~(Wryiw6 & Pujnv6));
assign E757x6 = (Ftyiw6 & U857x6);
assign U857x6 = (~(Fth7z6[25] & Ttyiw6));
assign Q657x6 = (~(Ivwnv6 & Fhc7z6[25]));
assign O557x6 = (B957x6 & I957x6);
assign I957x6 = (~(Dwwnv6 & Nqh7z6[25]));
assign B957x6 = (~(Kwwnv6 & Fth7z6[25]));
assign Bjy7v6 = (~(P957x6 & W957x6));
assign W957x6 = (Da57x6 & Ka57x6);
assign Ka57x6 = (~(Ztwnv6 & Kxb7z6[24]));
assign Da57x6 = (Ra57x6 & Ya57x6);
assign Ya57x6 = (~(Uuwnv6 & M3ynv6));
assign M3ynv6 = (~(Fb57x6 & Mb57x6));
assign Mb57x6 = (Tb57x6 & Ac57x6);
assign Ac57x6 = (~(Wryiw6 & Fwjnv6));
assign Tb57x6 = (Hc57x6 & Oc57x6);
assign Oc57x6 = (~(Zfhov6 & Rsyiw6));
assign Zfhov6 = (Xgmov6 ? Fd9ov6 : Td9ov6);
assign Hc57x6 = (~(Nqh7z6[24] & Ysyiw6));
assign Fb57x6 = (Ftyiw6 & Vc57x6);
assign Vc57x6 = (~(Fth7z6[24] & Ttyiw6));
assign Ra57x6 = (~(Ivwnv6 & Fhc7z6[24]));
assign P957x6 = (Cd57x6 & Jd57x6);
assign Jd57x6 = (~(Dwwnv6 & Nqh7z6[24]));
assign Cd57x6 = (~(Kwwnv6 & Fth7z6[24]));
assign Uiy7v6 = (~(Qd57x6 & Xd57x6));
assign Xd57x6 = (Ee57x6 & Le57x6);
assign Le57x6 = (~(Ztwnv6 & Kxb7z6[23]));
assign Ee57x6 = (Se57x6 & Ze57x6);
assign Ze57x6 = (~(Uuwnv6 & N7ynv6));
assign N7ynv6 = (~(Gf57x6 & Nf57x6));
assign Nf57x6 = (Uf57x6 & Bg57x6);
assign Bg57x6 = (~(Nqh7z6[23] & Ysyiw6));
assign Uf57x6 = (Ig57x6 & Pg57x6);
assign Pg57x6 = (~(Wg57x6 & Dh57x6));
assign Ig57x6 = (~(Kh57x6 & Rh57x6));
assign Gf57x6 = (Yh57x6 & Ftyiw6);
assign Yh57x6 = (Fi57x6 & Mi57x6);
assign Mi57x6 = (~(Wryiw6 & Vxjnv6));
assign Fi57x6 = (~(Fth7z6[23] & Ttyiw6));
assign Se57x6 = (~(Ivwnv6 & Fhc7z6[23]));
assign Qd57x6 = (Ti57x6 & Aj57x6);
assign Aj57x6 = (~(Dwwnv6 & Nqh7z6[23]));
assign Ti57x6 = (~(Kwwnv6 & Fth7z6[23]));
assign Niy7v6 = (~(Hj57x6 & Oj57x6));
assign Oj57x6 = (Vj57x6 & Ck57x6);
assign Ck57x6 = (~(Ztwnv6 & Kxb7z6[22]));
assign Vj57x6 = (Jk57x6 & Qk57x6);
assign Qk57x6 = (~(Uuwnv6 & Ccynv6));
assign Ccynv6 = (~(Xk57x6 & El57x6));
assign El57x6 = (Ll57x6 & Sl57x6);
assign Sl57x6 = (~(Nqh7z6[22] & Ysyiw6));
assign Ll57x6 = (Zl57x6 & Gm57x6);
assign Gm57x6 = (~(Wg57x6 & Nm57x6));
assign Zl57x6 = (~(Kh57x6 & Um57x6));
assign Xk57x6 = (Bn57x6 & Ftyiw6);
assign Bn57x6 = (In57x6 & Pn57x6);
assign Pn57x6 = (~(Wryiw6 & Lzjnv6));
assign In57x6 = (~(Fth7z6[22] & Ttyiw6));
assign Jk57x6 = (~(Ivwnv6 & Fhc7z6[22]));
assign Hj57x6 = (Wn57x6 & Do57x6);
assign Do57x6 = (~(Dwwnv6 & Nqh7z6[22]));
assign Wn57x6 = (~(Kwwnv6 & Fth7z6[22]));
assign Giy7v6 = (~(Ko57x6 & Ro57x6));
assign Ro57x6 = (Yo57x6 & Fp57x6);
assign Fp57x6 = (~(Ztwnv6 & Kxb7z6[21]));
assign Yo57x6 = (Mp57x6 & Tp57x6);
assign Tp57x6 = (~(Uuwnv6 & Rgynv6));
assign Rgynv6 = (~(Aq57x6 & Hq57x6));
assign Hq57x6 = (Oq57x6 & Vq57x6);
assign Vq57x6 = (~(Nqh7z6[21] & Ysyiw6));
assign Oq57x6 = (Cr57x6 & Jr57x6);
assign Jr57x6 = (~(Wg57x6 & Qr57x6));
assign Cr57x6 = (~(Kh57x6 & Xr57x6));
assign Aq57x6 = (Es57x6 & Ftyiw6);
assign Es57x6 = (Ls57x6 & Ss57x6);
assign Ss57x6 = (~(Wryiw6 & B1knv6));
assign Ls57x6 = (~(Fth7z6[21] & Ttyiw6));
assign Mp57x6 = (~(Ivwnv6 & Fhc7z6[21]));
assign Ko57x6 = (Zs57x6 & Gt57x6);
assign Gt57x6 = (~(Dwwnv6 & Nqh7z6[21]));
assign Zs57x6 = (~(Kwwnv6 & Fth7z6[21]));
assign Zhy7v6 = (~(Nt57x6 & Ut57x6));
assign Ut57x6 = (Bu57x6 & Iu57x6);
assign Iu57x6 = (~(Ztwnv6 & Kxb7z6[20]));
assign Bu57x6 = (Pu57x6 & Wu57x6);
assign Wu57x6 = (~(Uuwnv6 & Glynv6));
assign Glynv6 = (~(Dv57x6 & Kv57x6));
assign Kv57x6 = (Rv57x6 & Yv57x6);
assign Yv57x6 = (~(Nqh7z6[20] & Ysyiw6));
assign Rv57x6 = (Fw57x6 & Mw57x6);
assign Mw57x6 = (~(Wg57x6 & Tw57x6));
assign Fw57x6 = (~(Kh57x6 & Ax57x6));
assign Dv57x6 = (Hx57x6 & Ftyiw6);
assign Hx57x6 = (Ox57x6 & Vx57x6);
assign Vx57x6 = (~(Wryiw6 & R2knv6));
assign Ox57x6 = (~(Fth7z6[20] & Ttyiw6));
assign Pu57x6 = (~(Ivwnv6 & Fhc7z6[20]));
assign Nt57x6 = (Cy57x6 & Jy57x6);
assign Jy57x6 = (~(Dwwnv6 & Nqh7z6[20]));
assign Cy57x6 = (~(Kwwnv6 & Fth7z6[20]));
assign Shy7v6 = (~(Qy57x6 & Xy57x6));
assign Xy57x6 = (Ez57x6 & Lz57x6);
assign Lz57x6 = (~(Ztwnv6 & Kxb7z6[19]));
assign Ez57x6 = (Sz57x6 & Zz57x6);
assign Zz57x6 = (~(Uuwnv6 & Vpynv6));
assign Vpynv6 = (~(G067x6 & N067x6));
assign N067x6 = (U067x6 & B167x6);
assign B167x6 = (~(Nqh7z6[19] & Ysyiw6));
assign U067x6 = (I167x6 & P167x6);
assign P167x6 = (~(Wg57x6 & Onlov6));
assign I167x6 = (~(Kh57x6 & Hnlov6));
assign G067x6 = (W167x6 & Ftyiw6);
assign W167x6 = (D267x6 & K267x6);
assign K267x6 = (~(Wryiw6 & L6knv6));
assign D267x6 = (~(Fth7z6[19] & Ttyiw6));
assign Sz57x6 = (~(Ivwnv6 & Fhc7z6[19]));
assign Qy57x6 = (R267x6 & Y267x6);
assign Y267x6 = (~(Dwwnv6 & Nqh7z6[19]));
assign R267x6 = (~(Kwwnv6 & Fth7z6[19]));
assign Lhy7v6 = (~(F367x6 & M367x6));
assign M367x6 = (T367x6 & A467x6);
assign A467x6 = (~(Ztwnv6 & Kxb7z6[18]));
assign T367x6 = (H467x6 & O467x6);
assign O467x6 = (~(Uuwnv6 & Kuynv6));
assign Kuynv6 = (~(V467x6 & C567x6));
assign C567x6 = (J567x6 & Q567x6);
assign Q567x6 = (~(Nqh7z6[18] & Ysyiw6));
assign J567x6 = (X567x6 & E667x6);
assign E667x6 = (~(Wg57x6 & Kdfov6));
assign X567x6 = (~(Kh57x6 & Ddfov6));
assign V467x6 = (L667x6 & Ftyiw6);
assign L667x6 = (S667x6 & Z667x6);
assign Z667x6 = (~(Wryiw6 & B8knv6));
assign S667x6 = (~(Fth7z6[18] & Ttyiw6));
assign H467x6 = (~(Ivwnv6 & Fhc7z6[18]));
assign F367x6 = (G767x6 & N767x6);
assign N767x6 = (~(Dwwnv6 & Nqh7z6[18]));
assign G767x6 = (~(Kwwnv6 & Fth7z6[18]));
assign Ehy7v6 = (~(U767x6 & B867x6));
assign B867x6 = (I867x6 & P867x6);
assign P867x6 = (~(Ztwnv6 & Kxb7z6[17]));
assign I867x6 = (W867x6 & D967x6);
assign D967x6 = (~(Uuwnv6 & Zyynv6));
assign Zyynv6 = (~(K967x6 & R967x6));
assign R967x6 = (Y967x6 & Fa67x6);
assign Fa67x6 = (~(Nqh7z6[17] & Ysyiw6));
assign Y967x6 = (Ma67x6 & Ta67x6);
assign Ta67x6 = (~(Wg57x6 & Ab67x6));
assign Wg57x6 = (~(Xgmov6 | Hb67x6));
assign Ma67x6 = (~(Kh57x6 & Ob67x6));
assign Kh57x6 = (~(Hb67x6 | No7et6));
assign Hb67x6 = (!Rsyiw6);
assign K967x6 = (Vb67x6 & Ftyiw6);
assign Vb67x6 = (Cc67x6 & Jc67x6);
assign Jc67x6 = (~(Wryiw6 & R9knv6));
assign Cc67x6 = (~(Fth7z6[17] & Ttyiw6));
assign W867x6 = (~(Ivwnv6 & Fhc7z6[17]));
assign U767x6 = (Qc67x6 & Xc67x6);
assign Xc67x6 = (~(Dwwnv6 & Nqh7z6[17]));
assign Qc67x6 = (~(Kwwnv6 & Fth7z6[17]));
assign Xgy7v6 = (~(Ed67x6 & Ld67x6));
assign Ld67x6 = (Sd67x6 & Zd67x6);
assign Zd67x6 = (~(Ztwnv6 & Kxb7z6[16]));
assign Sd67x6 = (Ge67x6 & Ne67x6);
assign Ne67x6 = (~(Uuwnv6 & O3znv6));
assign O3znv6 = (~(Ue67x6 & Bf67x6));
assign Bf67x6 = (If67x6 & Pf67x6);
assign Pf67x6 = (~(Wryiw6 & Hbknv6));
assign If67x6 = (Wf67x6 & Dg67x6);
assign Dg67x6 = (~(Ykfov6 & Rsyiw6));
assign Wf67x6 = (~(Nqh7z6[16] & Ysyiw6));
assign Ue67x6 = (Ftyiw6 & Kg67x6);
assign Kg67x6 = (~(Fth7z6[16] & Ttyiw6));
assign Ge67x6 = (~(Ivwnv6 & Fhc7z6[16]));
assign Ed67x6 = (Rg67x6 & Yg67x6);
assign Yg67x6 = (~(Dwwnv6 & Nqh7z6[16]));
assign Rg67x6 = (~(Kwwnv6 & Fth7z6[16]));
assign Qgy7v6 = (Mh67x6 ? Fh67x6 : Fth7z6[15]);
assign Fh67x6 = (~(Th67x6 & Ai67x6));
assign Ai67x6 = (Hi67x6 & Oi67x6);
assign Oi67x6 = (Vi67x6 & Cj67x6);
assign Cj67x6 = (~(Jj67x6 & Dh57x6));
assign Vi67x6 = (Qj67x6 & Xj67x6);
assign Xj67x6 = (~(Ek67x6 & D8znv6));
assign D8znv6 = (~(Lk67x6 & Sk67x6));
assign Sk67x6 = (Zk67x6 & Gl67x6);
assign Gl67x6 = (~(Wryiw6 & Xcknv6));
assign Zk67x6 = (Nl67x6 & Ul67x6);
assign Ul67x6 = (~(Fzmov6 & Rsyiw6));
assign Nl67x6 = (~(Nqh7z6[15] & Ysyiw6));
assign Lk67x6 = (Ftyiw6 & Bm67x6);
assign Bm67x6 = (~(Fth7z6[15] & Ttyiw6));
assign Qj67x6 = (~(Im67x6 & Rh57x6));
assign Hi67x6 = (Pm67x6 & Wm67x6);
assign Wm67x6 = (~(Dn67x6 & Kn67x6));
assign Pm67x6 = (~(Rn67x6 & Zwlov6));
assign Th67x6 = (Yn67x6 & Fo67x6);
assign Fo67x6 = (Mo67x6 & To67x6);
assign To67x6 = (~(Ap67x6 & Hp67x6));
assign Mo67x6 = (~(Op67x6 & Fhc7z6[15]));
assign Yn67x6 = (Vp67x6 & Cq67x6);
assign Cq67x6 = (~(Kxb7z6[15] & Jq67x6));
assign Vp67x6 = (~(Qq67x6 & Nqh7z6[15]));
assign Jgy7v6 = (Mh67x6 ? Xq67x6 : Fth7z6[14]);
assign Xq67x6 = (~(Er67x6 & Lr67x6));
assign Lr67x6 = (Sr67x6 & Zr67x6);
assign Zr67x6 = (Gs67x6 & Ns67x6);
assign Ns67x6 = (~(Jj67x6 & Nm57x6));
assign Gs67x6 = (Us67x6 & Bt67x6);
assign Bt67x6 = (~(Ek67x6 & Ecznv6));
assign Ecznv6 = (~(It67x6 & Pt67x6));
assign Pt67x6 = (Wt67x6 & Du67x6);
assign Du67x6 = (~(Wryiw6 & Neknv6));
assign Wt67x6 = (Ku67x6 & Ru67x6);
assign Ru67x6 = (~(E2nov6 & Rsyiw6));
assign Ku67x6 = (~(Nqh7z6[14] & Ysyiw6));
assign It67x6 = (Ftyiw6 & Yu67x6);
assign Yu67x6 = (~(Fth7z6[14] & Ttyiw6));
assign Us67x6 = (~(Im67x6 & Um57x6));
assign Sr67x6 = (Fv67x6 & Mv67x6);
assign Mv67x6 = (~(Dn67x6 & Tv67x6));
assign Fv67x6 = (~(Rn67x6 & Xs9iw6));
assign Er67x6 = (Aw67x6 & Hw67x6);
assign Hw67x6 = (Ow67x6 & Vw67x6);
assign Vw67x6 = (~(Ap67x6 & Cx67x6));
assign Ow67x6 = (~(Op67x6 & Fhc7z6[14]));
assign Aw67x6 = (Jx67x6 & Qx67x6);
assign Qx67x6 = (~(Kxb7z6[14] & Jq67x6));
assign Jx67x6 = (~(Qq67x6 & Nqh7z6[14]));
assign Cgy7v6 = (Mh67x6 ? Xx67x6 : Fth7z6[13]);
assign Xx67x6 = (~(Ey67x6 & Ly67x6));
assign Ly67x6 = (Sy67x6 & Zy67x6);
assign Zy67x6 = (Gz67x6 & Nz67x6);
assign Nz67x6 = (~(Jj67x6 & Qr57x6));
assign Gz67x6 = (Uz67x6 & B077x6);
assign B077x6 = (~(Ek67x6 & Fgznv6));
assign Fgznv6 = (~(I077x6 & P077x6));
assign P077x6 = (W077x6 & D177x6);
assign D177x6 = (~(Wryiw6 & Dgknv6));
assign W077x6 = (K177x6 & R177x6);
assign R177x6 = (~(Ng9iw6 & Rsyiw6));
assign K177x6 = (~(Nqh7z6[13] & Ysyiw6));
assign I077x6 = (Ftyiw6 & Y177x6);
assign Y177x6 = (~(Fth7z6[13] & Ttyiw6));
assign Uz67x6 = (~(Im67x6 & Xr57x6));
assign Sy67x6 = (F277x6 & M277x6);
assign M277x6 = (~(Dn67x6 & T277x6));
assign F277x6 = (~(Rn67x6 & Qs9iw6));
assign Ey67x6 = (A377x6 & H377x6);
assign H377x6 = (O377x6 & V377x6);
assign V377x6 = (~(Ap67x6 & C477x6));
assign O377x6 = (~(Op67x6 & Fhc7z6[13]));
assign A377x6 = (J477x6 & Q477x6);
assign Q477x6 = (~(Kxb7z6[13] & Jq67x6));
assign J477x6 = (~(Qq67x6 & Nqh7z6[13]));
assign Vfy7v6 = (Mh67x6 ? X477x6 : Fth7z6[12]);
assign X477x6 = (~(E577x6 & L577x6));
assign L577x6 = (S577x6 & Z577x6);
assign Z577x6 = (G677x6 & N677x6);
assign N677x6 = (~(Jj67x6 & Tw57x6));
assign G677x6 = (U677x6 & B777x6);
assign B777x6 = (~(Ek67x6 & Gkznv6));
assign Gkznv6 = (~(I777x6 & P777x6));
assign P777x6 = (W777x6 & D877x6);
assign D877x6 = (~(Wryiw6 & Thknv6));
assign W777x6 = (K877x6 & R877x6);
assign R877x6 = (~(Tj9iw6 & Rsyiw6));
assign K877x6 = (~(Nqh7z6[12] & Ysyiw6));
assign I777x6 = (Ftyiw6 & Y877x6);
assign Y877x6 = (~(Fth7z6[12] & Ttyiw6));
assign U677x6 = (~(Im67x6 & Ax57x6));
assign S577x6 = (F977x6 & M977x6);
assign M977x6 = (~(Dn67x6 & T977x6));
assign F977x6 = (~(Rn67x6 & Js9iw6));
assign E577x6 = (Aa77x6 & Ha77x6);
assign Ha77x6 = (Oa77x6 & Va77x6);
assign Va77x6 = (~(Ap67x6 & Cb77x6));
assign Oa77x6 = (~(Op67x6 & Fhc7z6[12]));
assign Aa77x6 = (Jb77x6 & Qb77x6);
assign Qb77x6 = (~(Kxb7z6[12] & Jq67x6));
assign Jb77x6 = (~(Qq67x6 & Nqh7z6[12]));
assign Ofy7v6 = (Mh67x6 ? Xb77x6 : Fth7z6[11]);
assign Xb77x6 = (~(Ec77x6 & Lc77x6));
assign Lc77x6 = (Sc77x6 & Zc77x6);
assign Zc77x6 = (Gd77x6 & Nd77x6);
assign Nd77x6 = (~(Jj67x6 & Onlov6));
assign Gd77x6 = (Ud77x6 & Be77x6);
assign Be77x6 = (~(Ek67x6 & Hoznv6));
assign Hoznv6 = (~(Ie77x6 & Pe77x6));
assign Pe77x6 = (We77x6 & Df77x6);
assign Df77x6 = (~(Wryiw6 & Jjknv6));
assign We77x6 = (Kf77x6 & Rf77x6);
assign Rf77x6 = (~(Ph9iw6 & Rsyiw6));
assign Kf77x6 = (~(Nqh7z6[11] & Ysyiw6));
assign Ie77x6 = (Ftyiw6 & Yf77x6);
assign Yf77x6 = (~(Fth7z6[11] & Ttyiw6));
assign Ud77x6 = (~(Im67x6 & Hnlov6));
assign Sc77x6 = (Fg77x6 & Mg77x6);
assign Mg77x6 = (~(Dn67x6 & Fmlov6));
assign Fg77x6 = (~(Rn67x6 & Cs9iw6));
assign Ec77x6 = (Tg77x6 & Ah77x6);
assign Ah77x6 = (Hh77x6 & Oh77x6);
assign Oh77x6 = (~(Ap67x6 & Mmlov6));
assign Hh77x6 = (~(Op67x6 & Fhc7z6[11]));
assign Tg77x6 = (Vh77x6 & Ci77x6);
assign Ci77x6 = (~(Kxb7z6[11] & Jq67x6));
assign Vh77x6 = (~(Qq67x6 & Nqh7z6[11]));
assign Hfy7v6 = (Mh67x6 ? Ji77x6 : Fth7z6[10]);
assign Ji77x6 = (~(Qi77x6 & Xi77x6));
assign Xi77x6 = (Ej77x6 & Lj77x6);
assign Lj77x6 = (Sj77x6 & Zj77x6);
assign Zj77x6 = (~(Jj67x6 & Kdfov6));
assign Sj77x6 = (Gk77x6 & Nk77x6);
assign Nk77x6 = (~(Ek67x6 & Isznv6));
assign Isznv6 = (~(Uk77x6 & Bl77x6));
assign Bl77x6 = (Il77x6 & Pl77x6);
assign Pl77x6 = (~(Wryiw6 & Glknv6));
assign Il77x6 = (Wl77x6 & Dm77x6);
assign Dm77x6 = (~(Uanov6 & Rsyiw6));
assign Wl77x6 = (~(Nqh7z6[10] & Ysyiw6));
assign Uk77x6 = (Ftyiw6 & Km77x6);
assign Km77x6 = (~(Fth7z6[10] & Ttyiw6));
assign Gk77x6 = (~(Im67x6 & Ddfov6));
assign Ej77x6 = (Rm77x6 & Ym77x6);
assign Ym77x6 = (~(Dn67x6 & Bcfov6));
assign Rm77x6 = (~(Rn67x6 & Vr9iw6));
assign Qi77x6 = (Fn77x6 & Mn77x6);
assign Mn77x6 = (Tn77x6 & Ao77x6);
assign Ao77x6 = (~(Ap67x6 & Icfov6));
assign Tn77x6 = (~(Op67x6 & Fhc7z6[10]));
assign Fn77x6 = (Ho77x6 & Oo77x6);
assign Oo77x6 = (~(Kxb7z6[10] & Jq67x6));
assign Ho77x6 = (~(Qq67x6 & Nqh7z6[10]));
assign Afy7v6 = (Mh67x6 ? Vo77x6 : Fth7z6[9]);
assign Vo77x6 = (~(Cp77x6 & Jp77x6));
assign Jp77x6 = (Qp77x6 & Xp77x6);
assign Xp77x6 = (Eq77x6 & Lq77x6);
assign Lq77x6 = (~(Ek67x6 & Jwznv6));
assign Jwznv6 = (~(Sq77x6 & Zq77x6));
assign Zq77x6 = (Gr77x6 & Nr77x6);
assign Nr77x6 = (~(H737x6 & Rsyiw6));
assign Gr77x6 = (Ur77x6 & Bs77x6);
assign Bs77x6 = (~(Nqh7z6[9] & Ysyiw6));
assign Ur77x6 = (~(Wryiw6 & L7jnv6));
assign Sq77x6 = (Ftyiw6 & Is77x6);
assign Is77x6 = (~(Fth7z6[9] & Ttyiw6));
assign Eq77x6 = (Ps77x6 & Ws77x6);
assign Ws77x6 = (~(Im67x6 & Ob67x6));
assign Im67x6 = (Nvvnv6 & Dt77x6);
assign Dt77x6 = (~(Kt77x6 & Rt77x6));
assign Rt77x6 = (~(Di47x6 & Xgmov6));
assign Ps77x6 = (~(Jj67x6 & Ab67x6));
assign Jj67x6 = (~(Yt77x6 & Fu77x6));
assign Fu77x6 = (~(Mu77x6 & Di47x6));
assign Mu77x6 = (No7et6 & Nvvnv6);
assign Yt77x6 = (~(Tu77x6 & Av77x6));
assign Qp77x6 = (Hv77x6 & Ov77x6);
assign Ov77x6 = (~(Dn67x6 & Vv77x6));
assign Hv77x6 = (~(Rn67x6 & Or9iw6));
assign Cp77x6 = (Cw77x6 & Jw77x6);
assign Jw77x6 = (Qw77x6 & Xw77x6);
assign Xw77x6 = (~(Ap67x6 & Ex77x6));
assign Qw77x6 = (~(Op67x6 & Fhc7z6[9]));
assign Cw77x6 = (Lx77x6 & Sx77x6);
assign Sx77x6 = (~(Kxb7z6[9] & Jq67x6));
assign Lx77x6 = (~(Qq67x6 & Nqh7z6[9]));
assign Tey7v6 = (Mh67x6 ? Zx77x6 : Fth7z6[8]);
assign Zx77x6 = (~(Gy77x6 & Ny77x6));
assign Ny77x6 = (Uy77x6 & Bz77x6);
assign Bz77x6 = (Iz77x6 & Pz77x6);
assign Pz77x6 = (~(Nvvnv6 & Wz77x6));
assign Wz77x6 = (~(D087x6 & K087x6));
assign K087x6 = (~(Di47x6 & Ykfov6));
assign Ykfov6 = (Xgmov6 ? Ve9ov6 : Jf9ov6);
assign D087x6 = (R087x6 & Y087x6);
assign Y087x6 = (~(F187x6 & M187x6));
assign M187x6 = (Jf9ov6 & Xgmov6);
assign F187x6 = (I0c7z6[0] & Av77x6);
assign R087x6 = (~(T187x6 & A287x6));
assign T187x6 = (H287x6 & Ve9ov6);
assign Iz77x6 = (~(Dn67x6 & Fd9ov6));
assign Dn67x6 = (Tu77x6 & H287x6);
assign Tu77x6 = (O287x6 & I0c7z6[0]);
assign O287x6 = (Nvvnv6 & Xgmov6);
assign Uy77x6 = (V287x6 & C387x6);
assign C387x6 = (~(Ek67x6 & K00ov6));
assign K00ov6 = (~(J387x6 & Q387x6));
assign Q387x6 = (X387x6 & E487x6);
assign E487x6 = (~(Wryiw6 & P9jnv6));
assign X387x6 = (L487x6 & S487x6);
assign S487x6 = (~(Et9iw6 & Rsyiw6));
assign Et9iw6 = (!Pylov6);
assign Pylov6 = (No7et6 ? G587x6 : Z487x6);
assign L487x6 = (~(Nqh7z6[8] & Ysyiw6));
assign J387x6 = (Ftyiw6 & N587x6);
assign N587x6 = (~(Fth7z6[8] & Ttyiw6));
assign V287x6 = (~(Rn67x6 & Swlov6));
assign Swlov6 = (Xgmov6 ? Td9ov6 : Fd9ov6);
assign Rn67x6 = (Wh47x6 & Nvvnv6);
assign Gy77x6 = (U587x6 & B687x6);
assign B687x6 = (I687x6 & P687x6);
assign P687x6 = (~(Ap67x6 & Td9ov6));
assign Ap67x6 = (W687x6 & A287x6);
assign W687x6 = (Av77x6 & Nvvnv6);
assign I687x6 = (~(Op67x6 & Fhc7z6[8]));
assign U587x6 = (D787x6 & K787x6);
assign K787x6 = (~(Kxb7z6[8] & Jq67x6));
assign D787x6 = (~(Qq67x6 & Nqh7z6[8]));
assign Mey7v6 = (~(R787x6 & Y787x6));
assign Y787x6 = (F887x6 & M887x6);
assign M887x6 = (~(Ivwnv6 & Fhc7z6[7]));
assign F887x6 = (T887x6 & A987x6);
assign A987x6 = (~(Lf47x6 & H987x6));
assign H987x6 = (~(O987x6 & V987x6));
assign V987x6 = (Ca87x6 & Ja87x6);
assign Ja87x6 = (~(Bh47x6 & Rh57x6));
assign Ca87x6 = (Qa87x6 & Xa87x6);
assign Xa87x6 = (~(Wh47x6 & Ju1ov6));
assign Ju1ov6 = (Xgmov6 ? Kn67x6 : Hp67x6);
assign Qa87x6 = (~(Di47x6 & Fzmov6));
assign Fzmov6 = (No7et6 ? Rh57x6 : Dh57x6);
assign O987x6 = (Eb87x6 & Lb87x6);
assign Lb87x6 = (~(Yi47x6 & Hp67x6));
assign Eb87x6 = (Sb87x6 & Zb87x6);
assign Zb87x6 = (~(Tj47x6 & Dh57x6));
assign Sb87x6 = (~(Ak47x6 & Kn67x6));
assign T887x6 = (~(Uuwnv6 & L40ov6));
assign L40ov6 = (~(Gc87x6 & Nc87x6));
assign Nc87x6 = (Uc87x6 & Bd87x6);
assign Bd87x6 = (~(Wryiw6 & Fbjnv6));
assign Uc87x6 = (Id87x6 & Pd87x6);
assign Pd87x6 = (~(Zwlov6 & Rsyiw6));
assign Zwlov6 = (No7et6 ? Kn67x6 : Hp67x6);
assign Id87x6 = (~(Nqh7z6[7] & Ysyiw6));
assign Gc87x6 = (Ftyiw6 & Wd87x6);
assign Wd87x6 = (~(Fth7z6[7] & Ttyiw6));
assign R787x6 = (De87x6 & Ke87x6);
assign Ke87x6 = (~(Kwwnv6 & Fth7z6[7]));
assign De87x6 = (Re87x6 & Ye87x6);
assign Ye87x6 = (~(Ztwnv6 & Kxb7z6[7]));
assign Re87x6 = (~(Dwwnv6 & Nqh7z6[7]));
assign Fey7v6 = (~(Ff87x6 & Mf87x6));
assign Mf87x6 = (Tf87x6 & Ag87x6);
assign Ag87x6 = (~(Ivwnv6 & Fhc7z6[6]));
assign Tf87x6 = (Hg87x6 & Og87x6);
assign Og87x6 = (~(Lf47x6 & Vg87x6));
assign Vg87x6 = (~(Ch87x6 & Jh87x6));
assign Jh87x6 = (Qh87x6 & Xh87x6);
assign Xh87x6 = (~(Bh47x6 & Um57x6));
assign Qh87x6 = (Ei87x6 & Li87x6);
assign Li87x6 = (~(Wh47x6 & Tk2ov6));
assign Tk2ov6 = (Xgmov6 ? Tv67x6 : Cx67x6);
assign Ei87x6 = (~(Di47x6 & E2nov6));
assign E2nov6 = (No7et6 ? Um57x6 : Nm57x6);
assign Ch87x6 = (Si87x6 & Zi87x6);
assign Zi87x6 = (~(Yi47x6 & Cx67x6));
assign Si87x6 = (Gj87x6 & Nj87x6);
assign Nj87x6 = (~(Tj47x6 & Nm57x6));
assign Gj87x6 = (~(Ak47x6 & Tv67x6));
assign Hg87x6 = (~(Uuwnv6 & M80ov6));
assign M80ov6 = (~(Uj87x6 & Bk87x6));
assign Bk87x6 = (Ik87x6 & Pk87x6);
assign Pk87x6 = (~(Wryiw6 & Vcjnv6));
assign Ik87x6 = (Wk87x6 & Dl87x6);
assign Dl87x6 = (~(Xs9iw6 & Rsyiw6));
assign Xs9iw6 = (!Nxlov6);
assign Nxlov6 = (No7et6 ? Rl87x6 : Kl87x6);
assign Wk87x6 = (~(Nqh7z6[6] & Ysyiw6));
assign Uj87x6 = (Ftyiw6 & Yl87x6);
assign Yl87x6 = (~(Fth7z6[6] & Ttyiw6));
assign Ff87x6 = (Fm87x6 & Mm87x6);
assign Mm87x6 = (~(Kwwnv6 & Fth7z6[6]));
assign Fm87x6 = (Tm87x6 & An87x6);
assign An87x6 = (~(Ztwnv6 & Kxb7z6[6]));
assign Tm87x6 = (~(Dwwnv6 & Nqh7z6[6]));
assign Ydy7v6 = (~(Hn87x6 & On87x6));
assign On87x6 = (Vn87x6 & Co87x6);
assign Co87x6 = (~(Ivwnv6 & Fhc7z6[5]));
assign Vn87x6 = (Jo87x6 & Qo87x6);
assign Qo87x6 = (~(Lf47x6 & Xo87x6));
assign Xo87x6 = (~(Ep87x6 & Lp87x6));
assign Lp87x6 = (Sp87x6 & Zp87x6);
assign Zp87x6 = (~(Bh47x6 & Xr57x6));
assign Sp87x6 = (Gq87x6 & Nq87x6);
assign Nq87x6 = (~(Wh47x6 & Bnbov6));
assign Bnbov6 = (Xgmov6 ? T277x6 : C477x6);
assign Gq87x6 = (~(Di47x6 & Ng9iw6));
assign Ng9iw6 = (No7et6 ? Xr57x6 : Qr57x6);
assign Ep87x6 = (Uq87x6 & Br87x6);
assign Br87x6 = (~(Yi47x6 & C477x6));
assign Uq87x6 = (Ir87x6 & Pr87x6);
assign Pr87x6 = (~(Tj47x6 & Qr57x6));
assign Ir87x6 = (~(Ak47x6 & T277x6));
assign Jo87x6 = (~(Uuwnv6 & Nc0ov6));
assign Nc0ov6 = (~(Wr87x6 & Ds87x6));
assign Ds87x6 = (Ks87x6 & Rs87x6);
assign Rs87x6 = (~(Wryiw6 & Lejnv6));
assign Ks87x6 = (Ys87x6 & Ft87x6);
assign Ft87x6 = (~(Qs9iw6 & Rsyiw6));
assign Qs9iw6 = (!Gxlov6);
assign Gxlov6 = (No7et6 ? Tt87x6 : Mt87x6);
assign Ys87x6 = (~(Nqh7z6[5] & Ysyiw6));
assign Wr87x6 = (Ftyiw6 & Au87x6);
assign Au87x6 = (~(Fth7z6[5] & Ttyiw6));
assign Ftyiw6 = (Je47x6 & Elphw6);
assign Hn87x6 = (Hu87x6 & Ou87x6);
assign Ou87x6 = (~(Kwwnv6 & Fth7z6[5]));
assign Hu87x6 = (Vu87x6 & Cv87x6);
assign Cv87x6 = (~(Ztwnv6 & Kxb7z6[5]));
assign Vu87x6 = (~(Dwwnv6 & Nqh7z6[5]));
assign Rdy7v6 = (~(Jv87x6 & Qv87x6));
assign Qv87x6 = (Xv87x6 & Ew87x6);
assign Ew87x6 = (~(Ivwnv6 & E3c7z6[4]));
assign Xv87x6 = (Lw87x6 & Sw87x6);
assign Sw87x6 = (~(Lf47x6 & Zw87x6));
assign Zw87x6 = (~(Gx87x6 & Nx87x6));
assign Nx87x6 = (Ux87x6 & By87x6);
assign By87x6 = (~(Bh47x6 & Ax57x6));
assign Ux87x6 = (Iy87x6 & Py87x6);
assign Py87x6 = (~(Wh47x6 & My9ov6));
assign My9ov6 = (Xgmov6 ? T977x6 : Cb77x6);
assign Iy87x6 = (~(Di47x6 & Tj9iw6));
assign Tj9iw6 = (No7et6 ? Ax57x6 : Tw57x6);
assign Gx87x6 = (Wy87x6 & Dz87x6);
assign Dz87x6 = (~(Yi47x6 & Cb77x6));
assign Wy87x6 = (Kz87x6 & Rz87x6);
assign Rz87x6 = (~(Tj47x6 & Tw57x6));
assign Kz87x6 = (~(Ak47x6 & T977x6));
assign Lw87x6 = (~(Uuwnv6 & Og0ov6));
assign Og0ov6 = (~(Yz87x6 & F097x6));
assign F097x6 = (M097x6 & T097x6);
assign T097x6 = (~(Wryiw6 & Bgjnv6));
assign M097x6 = (A197x6 & H197x6);
assign H197x6 = (~(Js9iw6 & Rsyiw6));
assign Js9iw6 = (!Iylov6);
assign Iylov6 = (No7et6 ? V197x6 : O197x6);
assign A197x6 = (~(Nqh7z6[4] & Ysyiw6));
assign Yz87x6 = (C297x6 & Je47x6);
assign C297x6 = (J297x6 & Q297x6);
assign Q297x6 = (~(Fth7z6[4] & Ttyiw6));
assign J297x6 = (~(Uyb7z6[4] & Ef47x6));
assign Jv87x6 = (X297x6 & E397x6);
assign E397x6 = (~(Kwwnv6 & Fth7z6[4]));
assign X297x6 = (L397x6 & S397x6);
assign S397x6 = (~(Ztwnv6 & Kxb7z6[4]));
assign L397x6 = (~(Dwwnv6 & Nqh7z6[4]));
assign Kdy7v6 = (~(Z397x6 & G497x6));
assign G497x6 = (N497x6 & U497x6);
assign U497x6 = (~(Ivwnv6 & E3c7z6[3]));
assign N497x6 = (B597x6 & I597x6);
assign I597x6 = (~(Lf47x6 & P597x6));
assign P597x6 = (~(W597x6 & D697x6));
assign D697x6 = (K697x6 & R697x6);
assign R697x6 = (~(Bh47x6 & Hnlov6));
assign K697x6 = (Y697x6 & F797x6);
assign F797x6 = (~(Wh47x6 & Htfov6));
assign Htfov6 = (Xgmov6 ? Fmlov6 : Mmlov6);
assign Y697x6 = (~(Di47x6 & Ph9iw6));
assign Ph9iw6 = (!Cl9iw6);
assign Cl9iw6 = (No7et6 ? T797x6 : M797x6);
assign W597x6 = (A897x6 & H897x6);
assign H897x6 = (~(Yi47x6 & Mmlov6));
assign A897x6 = (O897x6 & V897x6);
assign V897x6 = (~(Tj47x6 & Onlov6));
assign O897x6 = (~(Ak47x6 & Fmlov6));
assign B597x6 = (~(Uuwnv6 & Pk0ov6));
assign Pk0ov6 = (~(C997x6 & J997x6));
assign J997x6 = (Q997x6 & X997x6);
assign X997x6 = (~(Wryiw6 & Rhjnv6));
assign Q997x6 = (Ea97x6 & La97x6);
assign La97x6 = (~(Cs9iw6 & Rsyiw6));
assign Cs9iw6 = (!Lwlov6);
assign Lwlov6 = (No7et6 ? Za97x6 : Sa97x6);
assign Ea97x6 = (~(Nqh7z6[3] & Ysyiw6));
assign C997x6 = (Gb97x6 & Je47x6);
assign Gb97x6 = (Nb97x6 & Ub97x6);
assign Ub97x6 = (~(Fth7z6[3] & Ttyiw6));
assign Nb97x6 = (~(Uyb7z6[3] & Ef47x6));
assign Z397x6 = (Bc97x6 & Ic97x6);
assign Ic97x6 = (~(Kwwnv6 & Fth7z6[3]));
assign Bc97x6 = (Pc97x6 & Wc97x6);
assign Wc97x6 = (~(Ztwnv6 & Kxb7z6[3]));
assign Pc97x6 = (~(Dwwnv6 & Nqh7z6[3]));
assign Ddy7v6 = (~(Dd97x6 & Kd97x6));
assign Kd97x6 = (Rd97x6 & Yd97x6);
assign Yd97x6 = (~(Ivwnv6 & E3c7z6[2]));
assign Rd97x6 = (Fe97x6 & Me97x6);
assign Me97x6 = (~(Lf47x6 & Te97x6));
assign Te97x6 = (~(Af97x6 & Hf97x6));
assign Hf97x6 = (Of97x6 & Vf97x6);
assign Vf97x6 = (~(Bh47x6 & Ddfov6));
assign Of97x6 = (Cg97x6 & Jg97x6);
assign Jg97x6 = (~(Wh47x6 & Q2mov6));
assign Q2mov6 = (!Xl9iw6);
assign Xl9iw6 = (No7et6 ? Xg97x6 : Qg97x6);
assign Cg97x6 = (~(Di47x6 & Uanov6));
assign Uanov6 = (!Ql9iw6);
assign Ql9iw6 = (No7et6 ? Lh97x6 : Eh97x6);
assign Af97x6 = (Sh97x6 & Zh97x6);
assign Zh97x6 = (~(Yi47x6 & Icfov6));
assign Sh97x6 = (Gi97x6 & Ni97x6);
assign Ni97x6 = (~(Tj47x6 & Kdfov6));
assign Gi97x6 = (~(Ak47x6 & Bcfov6));
assign Fe97x6 = (~(Uuwnv6 & Qo0ov6));
assign Qo0ov6 = (~(Ui97x6 & Bj97x6));
assign Bj97x6 = (Ij97x6 & Pj97x6);
assign Pj97x6 = (~(Wryiw6 & Nmjnv6));
assign Ij97x6 = (Wj97x6 & Dk97x6);
assign Dk97x6 = (~(Nqh7z6[2] & Kk97x6));
assign Kk97x6 = (~(Rk97x6 & Yk97x6));
assign Yk97x6 = (Fl97x6 | Hfliw6);
assign Fl97x6 = (Ml97x6 | Ir7et6);
assign Wj97x6 = (~(Vr9iw6 & Rsyiw6));
assign Vr9iw6 = (!Wylov6);
assign Wylov6 = (No7et6 ? Qg97x6 : Xg97x6);
assign Ui97x6 = (Tl97x6 & Je47x6);
assign Tl97x6 = (Am97x6 & Hm97x6);
assign Hm97x6 = (~(Fth7z6[2] & Ttyiw6));
assign Am97x6 = (~(Uyb7z6[2] & Ef47x6));
assign Dd97x6 = (Om97x6 & Vm97x6);
assign Vm97x6 = (~(Kwwnv6 & Fth7z6[2]));
assign Om97x6 = (Cn97x6 & Jn97x6);
assign Jn97x6 = (~(Ztwnv6 & Kxb7z6[2]));
assign Cn97x6 = (~(Dwwnv6 & Nqh7z6[2]));
assign Wcy7v6 = (~(Qn97x6 & Xn97x6));
assign Xn97x6 = (Eo97x6 & Lo97x6);
assign Lo97x6 = (~(Ivwnv6 & E3c7z6[1]));
assign Ivwnv6 = (Op67x6 & Mh67x6);
assign Op67x6 = (~(So97x6 | Zo97x6));
assign So97x6 = (~(Gp97x6 & Np97x6));
assign Eo97x6 = (Up97x6 & Bq97x6);
assign Bq97x6 = (Z847x6 | Kdmhw6);
assign Kdmhw6 = (Iq97x6 & Pq97x6);
assign Pq97x6 = (Wq97x6 & Dr97x6);
assign Dr97x6 = (~(Or9iw6 & Rsyiw6));
assign Rsyiw6 = (~(Kr97x6 & Rr97x6));
assign Rr97x6 = (Yr97x6 & Fs97x6);
assign Fs97x6 = (~(Ms97x6 & Clhhw6));
assign Yr97x6 = (~(Ts97x6 | Ztaov6));
assign Kr97x6 = (At97x6 & Ht97x6);
assign Ht97x6 = (~(Ot97x6 & Vt97x6));
assign Or9iw6 = (!Dzlov6);
assign Dzlov6 = (No7et6 ? Ju97x6 : Cu97x6);
assign Wq97x6 = (Qu97x6 & Xu97x6);
assign Xu97x6 = (~(Nqh7z6[1] & Ysyiw6));
assign Ysyiw6 = (~(Rk97x6 & Ml97x6));
assign Ml97x6 = (~(Puphw6 | Lyknv6));
assign Puphw6 = (!Eminv6);
assign Rk97x6 = (Ev97x6 & Lv97x6);
assign Lv97x6 = (~(Sv97x6 & Vxihw6));
assign Qu97x6 = (Vd47x6 | J5knv6);
assign Vd47x6 = (!Wryiw6);
assign Wryiw6 = (Zv97x6 & Kb47x6);
assign Zv97x6 = (~(Uebdt6 | R3h7z6[0]));
assign Iq97x6 = (Gw97x6 & Je47x6);
assign Je47x6 = (Nw97x6 & Uw97x6);
assign Nw97x6 = (Bx97x6 & Ix97x6);
assign Bx97x6 = (~(Px97x6 & Dwb7z6[5]));
assign Gw97x6 = (Wx97x6 & Dy97x6);
assign Dy97x6 = (~(Fth7z6[1] & Ttyiw6));
assign Ttyiw6 = (Ky97x6 | Ry97x6);
assign Ky97x6 = (~(Yy97x6 & Fz97x6));
assign Fz97x6 = (~(Uebdt6 & Kb47x6));
assign Kb47x6 = (~(Mz97x6 & Tz97x6));
assign Tz97x6 = (~(A0a7x6 & Ev97x6));
assign Ev97x6 = (H0a7x6 & O0a7x6);
assign O0a7x6 = (V0a7x6 & C1a7x6);
assign C1a7x6 = (J1a7x6 & Xxknv6);
assign V0a7x6 = (Q1a7x6 & X1a7x6);
assign H0a7x6 = (E2a7x6 & L2a7x6);
assign L2a7x6 = (~(S2a7x6 & Dwb7z6[3]));
assign E2a7x6 = (Z2a7x6 & G3a7x6);
assign A0a7x6 = (Ywaov6 & Bwvnv6);
assign Mz97x6 = (N3a7x6 & U3a7x6);
assign Yy97x6 = (Twphw6 | Ms97x6);
assign Ms97x6 = (B4a7x6 & I4a7x6);
assign I4a7x6 = (~(P4a7x6 & W4a7x6));
assign P4a7x6 = (Tnzdt6 & Vxihw6);
assign B4a7x6 = (~(D5a7x6 & K5a7x6));
assign K5a7x6 = (~(R5a7x6 & Bfo7v6));
assign R5a7x6 = (~(E9nov6 & Y5a7x6));
assign Y5a7x6 = (~(F6a7x6 & M6a7x6));
assign Wx97x6 = (~(Uyb7z6[1] & Ef47x6));
assign Z847x6 = (~(T6a7x6 & Uuwnv6));
assign Uuwnv6 = (Ek67x6 & Mh67x6);
assign Ek67x6 = (~(Np97x6 | A7a7x6));
assign T6a7x6 = (T3cdt6 ? O7a7x6 : H7a7x6);
assign O7a7x6 = (~(V7a7x6 & C8a7x6));
assign H7a7x6 = (~(J8a7x6 & Pdlhw6));
assign Up97x6 = (~(Lf47x6 & Q8a7x6));
assign Q8a7x6 = (~(X8a7x6 & E9a7x6));
assign E9a7x6 = (L9a7x6 & S9a7x6);
assign S9a7x6 = (~(Ak47x6 & Vv77x6));
assign Ak47x6 = (~(Z9a7x6 & Kt77x6));
assign Kt77x6 = (~(A287x6 & H287x6));
assign Z9a7x6 = (~(Gaa7x6 & Naa7x6));
assign L9a7x6 = (Uaa7x6 & Bba7x6);
assign Bba7x6 = (~(Bh47x6 & Ob67x6));
assign Bh47x6 = (~(Iba7x6 | A287x6));
assign Uaa7x6 = (~(Tj47x6 & Ab67x6));
assign Tj47x6 = (~(Pba7x6 & Wba7x6));
assign Wba7x6 = (~(A287x6 & Av77x6));
assign Pba7x6 = (~(Dca7x6 & Naa7x6));
assign X8a7x6 = (Kca7x6 & Rca7x6);
assign Rca7x6 = (~(Yi47x6 & Ex77x6));
assign Yi47x6 = (~(Yca7x6 | A287x6));
assign A287x6 = (I0c7z6[0] & No7et6);
assign Kca7x6 = (Fda7x6 & Mda7x6);
assign Mda7x6 = (~(Wh47x6 & Od9iw6));
assign Od9iw6 = (!Jl9iw6);
assign Jl9iw6 = (No7et6 ? Cu97x6 : Ju97x6);
assign Wh47x6 = (~(Naa7x6 | Tda7x6));
assign Fda7x6 = (~(Di47x6 & H737x6));
assign H737x6 = (Xgmov6 ? Ab67x6 : Ob67x6);
assign Di47x6 = (~(Naa7x6 | Aea7x6));
assign Naa7x6 = (!I0c7z6[0]);
assign Lf47x6 = (Nvvnv6 & Mh67x6);
assign Qn97x6 = (Hea7x6 & Oea7x6);
assign Oea7x6 = (~(Kwwnv6 & Fth7z6[1]));
assign Kwwnv6 = (!Mh67x6);
assign Hea7x6 = (Vea7x6 & Cfa7x6);
assign Cfa7x6 = (~(Ztwnv6 & Kxb7z6[1]));
assign Ztwnv6 = (Jq67x6 & Mh67x6);
assign Jq67x6 = (~(Jfa7x6 & Qfa7x6));
assign Qfa7x6 = (~(Xfa7x6 & Ega7x6));
assign Jfa7x6 = (Lga7x6 & Sga7x6);
assign Lga7x6 = (~(Zga7x6 & Gp97x6));
assign Gp97x6 = (!A7a7x6);
assign A7a7x6 = (Gha7x6 & Mulnv6);
assign Zga7x6 = (Zo97x6 & Np97x6);
assign Np97x6 = (~(Nha7x6 & Uha7x6));
assign Nha7x6 = (Vi7et6 & P2jnv6);
assign Zo97x6 = (~(Bia7x6 & Uha7x6));
assign Bia7x6 = (T3cdt6 & P2jnv6);
assign Vea7x6 = (~(Dwwnv6 & Nqh7z6[1]));
assign Dwwnv6 = (Qq67x6 & Mh67x6);
assign Mh67x6 = (~(Iia7x6 & Pia7x6));
assign Pia7x6 = (Wia7x6 & Dja7x6);
assign Dja7x6 = (~(Gr2et6 & Kja7x6));
assign Kja7x6 = (~(Rja7x6 & Yja7x6));
assign Yja7x6 = (~(Fka7x6 & Vxihw6));
assign Fka7x6 = (Mka7x6 & Tka7x6);
assign Mka7x6 = (~(Wbxdt6 & B2jnv6));
assign Wia7x6 = (~(Ala7x6 & Hla7x6));
assign Hla7x6 = (Ola7x6 & Tka7x6);
assign Ola7x6 = (~(Vla7x6 & Vi7et6));
assign Vla7x6 = (Wbxdt6 & Ii9ov6);
assign Ala7x6 = (T3cdt6 & O5a7z6);
assign Iia7x6 = (Cma7x6 & Jma7x6);
assign Jma7x6 = (Qma7x6 | Xma7x6);
assign Qma7x6 = (~(O5a7z6 & Qg2nv6));
assign Cma7x6 = (~(Ena7x6 & Lna7x6));
assign Ena7x6 = (Nhonv6 & Sna7x6);
assign Qq67x6 = (~(Ega7x6 | Zna7x6));
assign Ega7x6 = (~(Goa7x6 & Noa7x6));
assign Goa7x6 = (Uoa7x6 & Yioov6);
assign Uoa7x6 = (~(Ecc7z6[11] & X4xiw6));
assign Pcy7v6 = (Bpa7x6 | Ipa7x6);
assign Ipa7x6 = (Ppa7x6 & Wpa7x6);
assign Wpa7x6 = (Dqa7x6 & Lidiw6);
assign Dqa7x6 = (~(O5a7z6 & Kqa7x6));
assign Kqa7x6 = (~(Fsmov6 & Rqa7x6));
assign Rqa7x6 = (~(Uha7x6 & Qodiw6));
assign Uha7x6 = (~(Zzihw6 | Nhonv6));
assign Ppa7x6 = (X4xiw6 & Vxihw6);
assign Bpa7x6 = (Lidiw6 ? Yqa7x6 : U6i7z6[1]);
assign Lidiw6 = (!Sidiw6);
assign Sidiw6 = (Fra7x6 & Xnmov6);
assign Xnmov6 = (~(Atmov6 & Nhonv6));
assign Fra7x6 = (~(Gr2et6 & Mra7x6));
assign Mra7x6 = (~(B3wnv6 & Rja7x6));
assign B3wnv6 = (!Fsmov6);
assign Yqa7x6 = (Tra7x6 & Asa7x6);
assign Asa7x6 = (~(Hsa7x6 | Ecc7z6[10]));
assign Tra7x6 = (G6xiw6 & X4xiw6);
assign Icy7v6 = (Osa7x6 & Vsa7x6);
assign Vsa7x6 = (~(Cta7x6 | Jta7x6));
assign Bcy7v6 = (~(Qta7x6 & Xta7x6));
assign Xta7x6 = (~(Eua7x6 & Zamov6));
assign Eua7x6 = (Ldo7v6 & Lua7x6);
assign Qta7x6 = (~(Sua7x6 & Xsinv6));
assign Sua7x6 = (~(Zua7x6 & Gva7x6));
assign Gva7x6 = (Nva7x6 & Uva7x6);
assign Nva7x6 = (Bwa7x6 & Iwa7x6);
assign Bwa7x6 = (~(Pwa7x6 & Mlmov6));
assign Pwa7x6 = (~(Wwa7x6 & Dxa7x6));
assign Dxa7x6 = (Losiw6 | Sfoov6);
assign Zua7x6 = (Kxa7x6 & Wwgov6);
assign Kxa7x6 = (Vmsiw6 & Rxa7x6);
assign Rxa7x6 = (Sfoov6 | Gd77z6);
assign Uby7v6 = (Yxa7x6 & Fya7x6);
assign Fya7x6 = (~(Kihov6 & Mya7x6));
assign Mya7x6 = (~(Teliw6 & Tya7x6));
assign Tya7x6 = (~(Aza7x6 & Hza7x6));
assign Hza7x6 = (~(Oza7x6 & Vza7x6));
assign Vza7x6 = (~(X0wnv6 & Wqsiw6));
assign Wqsiw6 = (~(Gpmov6 & C0b7x6));
assign Oza7x6 = (Qv0ov6 & J0b7x6);
assign Aza7x6 = (~(Q0b7x6 & Tnzdt6));
assign Q0b7x6 = (X0b7x6 & Lua7x6);
assign Kihov6 = (~(Phhov6 & Mlfov6));
assign Yxa7x6 = (~(E1b7x6 & Nrsnv6));
assign Nrsnv6 = (!Ac77z6);
assign Nby7v6 = (Wkb7z6[0] | L1b7x6);
assign L1b7x6 = (Bzi7z6[0] & S1b7x6);
assign S1b7x6 = (~(Z1b7x6 & U42nv6));
assign Gby7v6 = (~(Jm8iw6 & G2b7x6));
assign G2b7x6 = (~(Bzi7z6[25] & N2b7x6));
assign N2b7x6 = (~(U2b7x6 & Iklov6));
assign Zay7v6 = (Zjb7z6[8] | B3b7x6);
assign B3b7x6 = (Bzi7z6[24] & I3b7x6);
assign I3b7x6 = (~(U2b7x6 & Wf4iw6));
assign U2b7x6 = (P3b7x6 & Bqi7z6[3]);
assign Say7v6 = (~(W3b7x6 & D4b7x6));
assign D4b7x6 = (~(Bzi7z6[19] & K4b7x6));
assign K4b7x6 = (~(R4b7x6 & Mn5iw6));
assign Lay7v6 = (~(Y4b7x6 & Qc77z6));
assign Y4b7x6 = (Wwgov6 & F5b7x6);
assign F5b7x6 = (~(Bzi7z6[18] & M5b7x6));
assign M5b7x6 = (~(R4b7x6 & Jp5iw6));
assign Eay7v6 = (~(T5b7x6 & A6b7x6));
assign A6b7x6 = (~(Bzi7z6[17] & H6b7x6));
assign H6b7x6 = (~(R4b7x6 & Gr5iw6));
assign X9y7v6 = (~(O6b7x6 & V6b7x6));
assign V6b7x6 = (~(Bzi7z6[16] & C7b7x6));
assign C7b7x6 = (~(R4b7x6 & Is5iw6));
assign R4b7x6 = (P3b7x6 & Bqi7z6[2]);
assign J9y7v6 = (~(Losiw6 & Q7b7x6));
assign Q7b7x6 = (~(Bzi7z6[12] & X7b7x6));
assign X7b7x6 = (~(J7b7x6 & Emhov6));
assign C9y7v6 = (~(Zosiw6 & E8b7x6));
assign E8b7x6 = (~(Bzi7z6[11] & L8b7x6));
assign L8b7x6 = (~(J7b7x6 & Dz6iw6));
assign Zosiw6 = (!Tlb7z6[3]);
assign V8y7v6 = (~(S8b7x6 & Z8b7x6));
assign Z8b7x6 = (~(Bzi7z6[10] & G9b7x6));
assign G9b7x6 = (~(J7b7x6 & H17iw6));
assign O8y7v6 = (~(N9b7x6 & U9b7x6));
assign U9b7x6 = (~(Bzi7z6[9] & Bab7x6));
assign Bab7x6 = (~(J7b7x6 & J27iw6));
assign H8y7v6 = (Tlb7z6[0] | Iab7x6);
assign Iab7x6 = (Bzi7z6[8] & Pab7x6);
assign Pab7x6 = (~(J7b7x6 & U47iw6));
assign J7b7x6 = (P3b7x6 & Bqi7z6[1]);
assign T7y7v6 = (~(Wab7x6 & Dbb7x6));
assign Dbb7x6 = (~(Kbb7x6 & R62nv6));
assign Wab7x6 = (Rbb7x6 & Ybb7x6);
assign Ybb7x6 = (~(Fcb7x6 & Cmm7z6[7]));
assign Rbb7x6 = (~(Mcb7x6 & Wui7z6[7]));
assign M7y7v6 = (~(Tcb7x6 & Adb7x6));
assign Adb7x6 = (~(Kbb7x6 & B52nv6));
assign Tcb7x6 = (Hdb7x6 & Odb7x6);
assign Odb7x6 = (~(Fcb7x6 & Cmm7z6[1]));
assign Hdb7x6 = (~(Mcb7x6 & Wui7z6[1]));
assign F7y7v6 = (~(Vdb7x6 & Ceb7x6));
assign Ceb7x6 = (~(Kbb7x6 & I52nv6));
assign Vdb7x6 = (Jeb7x6 & Qeb7x6);
assign Qeb7x6 = (~(Fcb7x6 & Yefnv6));
assign Jeb7x6 = (~(Mcb7x6 & Wui7z6[2]));
assign Y6y7v6 = (~(Xeb7x6 & Efb7x6));
assign Efb7x6 = (~(Kbb7x6 & P52nv6));
assign Xeb7x6 = (Lfb7x6 & Sfb7x6);
assign Sfb7x6 = (~(Fcb7x6 & Cmm7z6[3]));
assign Lfb7x6 = (~(Mcb7x6 & Wui7z6[3]));
assign R6y7v6 = (~(Zfb7x6 & Ggb7x6));
assign Ggb7x6 = (~(Kbb7x6 & W52nv6));
assign Zfb7x6 = (Ngb7x6 & Ugb7x6);
assign Ugb7x6 = (~(Fcb7x6 & Cmm7z6[4]));
assign Ngb7x6 = (~(Mcb7x6 & Wui7z6[4]));
assign K6y7v6 = (~(Bhb7x6 & Ihb7x6));
assign Ihb7x6 = (~(Kbb7x6 & D62nv6));
assign Bhb7x6 = (Phb7x6 & Whb7x6);
assign Whb7x6 = (~(Fcb7x6 & Cmm7z6[5]));
assign Phb7x6 = (~(Mcb7x6 & Wui7z6[5]));
assign D6y7v6 = (~(Dib7x6 & Kib7x6));
assign Kib7x6 = (~(Kbb7x6 & K62nv6));
assign Dib7x6 = (Rib7x6 & Yib7x6);
assign Yib7x6 = (~(Fcb7x6 & Cmm7z6[6]));
assign Rib7x6 = (~(Mcb7x6 & Wui7z6[6]));
assign W5y7v6 = (~(Fjb7x6 & Mjb7x6));
assign Mjb7x6 = (~(Kbb7x6 & U42nv6));
assign Fjb7x6 = (Tjb7x6 & Akb7x6);
assign Akb7x6 = (~(Fcb7x6 & Cmm7z6[0]));
assign Fcb7x6 = (~(Mcb7x6 | Kbb7x6));
assign Tjb7x6 = (~(Mcb7x6 & Wui7z6[0]));
assign Mcb7x6 = (~(Kbb7x6 | Hkb7x6));
assign Kbb7x6 = (~(Okb7x6 | Twaiw6));
assign P5y7v6 = (~(Vkb7x6 & Clb7x6));
assign Clb7x6 = (~(Jlb7x6 & Z0iov6));
assign Vkb7x6 = (Qlb7x6 & Xlb7x6);
assign Xlb7x6 = (~(Emb7x6 & Cmm7z6[15]));
assign Qlb7x6 = (~(Lmb7x6 & Wui7z6[15]));
assign I5y7v6 = (~(Smb7x6 & Zmb7x6));
assign Zmb7x6 = (~(Jlb7x6 & U47iw6));
assign Smb7x6 = (Gnb7x6 & Nnb7x6);
assign Nnb7x6 = (~(Emb7x6 & Cmm7z6[8]));
assign Gnb7x6 = (~(Lmb7x6 & Wui7z6[8]));
assign B5y7v6 = (~(Unb7x6 & Bob7x6));
assign Bob7x6 = (~(Jlb7x6 & J27iw6));
assign Unb7x6 = (Iob7x6 & Pob7x6);
assign Pob7x6 = (~(Emb7x6 & Cmm7z6[9]));
assign Iob7x6 = (~(Lmb7x6 & Wui7z6[9]));
assign U4y7v6 = (~(Wob7x6 & Dpb7x6));
assign Dpb7x6 = (~(Jlb7x6 & H17iw6));
assign Wob7x6 = (Kpb7x6 & Rpb7x6);
assign Rpb7x6 = (~(Emb7x6 & Cmm7z6[10]));
assign Kpb7x6 = (~(Lmb7x6 & Wui7z6[10]));
assign N4y7v6 = (~(Ypb7x6 & Fqb7x6));
assign Fqb7x6 = (~(Jlb7x6 & Dz6iw6));
assign Ypb7x6 = (Mqb7x6 & Tqb7x6);
assign Tqb7x6 = (~(Emb7x6 & Cmm7z6[11]));
assign Mqb7x6 = (~(Lmb7x6 & Wui7z6[11]));
assign G4y7v6 = (~(Arb7x6 & Hrb7x6));
assign Hrb7x6 = (~(Jlb7x6 & Emhov6));
assign Arb7x6 = (Orb7x6 & Vrb7x6);
assign Vrb7x6 = (~(Emb7x6 & Cmm7z6[12]));
assign Orb7x6 = (~(Lmb7x6 & Wui7z6[12]));
assign Z3y7v6 = (~(Csb7x6 & Jsb7x6));
assign Jsb7x6 = (~(Jlb7x6 & Guhov6));
assign Csb7x6 = (Qsb7x6 & Xsb7x6);
assign Xsb7x6 = (~(Emb7x6 & Cmm7z6[13]));
assign Qsb7x6 = (~(Lmb7x6 & Wui7z6[13]));
assign S3y7v6 = (~(Etb7x6 & Ltb7x6));
assign Ltb7x6 = (~(Jlb7x6 & Bk6iw6));
assign Etb7x6 = (Stb7x6 & Ztb7x6);
assign Ztb7x6 = (~(Emb7x6 & Cmm7z6[14]));
assign Emb7x6 = (~(Lmb7x6 | Jlb7x6));
assign Stb7x6 = (~(Lmb7x6 & Wui7z6[14]));
assign Lmb7x6 = (~(Jlb7x6 | Hkb7x6));
assign Jlb7x6 = (~(Okb7x6 | Nq6iw6));
assign L3y7v6 = (~(Gub7x6 & Nub7x6));
assign Nub7x6 = (~(Uub7x6 & Cx4iw6));
assign Gub7x6 = (Bvb7x6 & Ivb7x6);
assign Ivb7x6 = (~(Pvb7x6 & Cmm7z6[23]));
assign Bvb7x6 = (~(Wvb7x6 & Wui7z6[23]));
assign E3y7v6 = (~(Dwb7x6 & Kwb7x6));
assign Kwb7x6 = (~(Uub7x6 & Is5iw6));
assign Dwb7x6 = (Rwb7x6 & Ywb7x6);
assign Ywb7x6 = (~(Pvb7x6 & Cmm7z6[16]));
assign Rwb7x6 = (~(Wvb7x6 & Wui7z6[16]));
assign X2y7v6 = (~(Fxb7x6 & Mxb7x6));
assign Mxb7x6 = (~(Uub7x6 & Gr5iw6));
assign Fxb7x6 = (Txb7x6 & Ayb7x6);
assign Ayb7x6 = (~(Pvb7x6 & Cmm7z6[17]));
assign Txb7x6 = (~(Wvb7x6 & Wui7z6[17]));
assign Q2y7v6 = (~(Hyb7x6 & Oyb7x6));
assign Oyb7x6 = (~(Uub7x6 & Jp5iw6));
assign Hyb7x6 = (Vyb7x6 & Czb7x6);
assign Czb7x6 = (~(Pvb7x6 & Cmm7z6[18]));
assign Vyb7x6 = (~(Wvb7x6 & Wui7z6[18]));
assign J2y7v6 = (~(Jzb7x6 & Qzb7x6));
assign Qzb7x6 = (~(Uub7x6 & Mn5iw6));
assign Jzb7x6 = (Xzb7x6 & E0c7x6);
assign E0c7x6 = (~(Pvb7x6 & Cmm7z6[19]));
assign Xzb7x6 = (~(Wvb7x6 & Wui7z6[19]));
assign C2y7v6 = (~(L0c7x6 & S0c7x6));
assign S0c7x6 = (~(Uub7x6 & Bl5iw6));
assign L0c7x6 = (Z0c7x6 & G1c7x6);
assign G1c7x6 = (~(Pvb7x6 & Cmm7z6[20]));
assign Z0c7x6 = (~(Wvb7x6 & Wui7z6[20]));
assign V1y7v6 = (~(N1c7x6 & U1c7x6));
assign U1c7x6 = (~(Uub7x6 & Ej5iw6));
assign N1c7x6 = (B2c7x6 & I2c7x6);
assign I2c7x6 = (~(Pvb7x6 & Cmm7z6[21]));
assign B2c7x6 = (~(Wvb7x6 & Wui7z6[21]));
assign O1y7v6 = (~(P2c7x6 & W2c7x6));
assign W2c7x6 = (~(Uub7x6 & D85iw6));
assign P2c7x6 = (D3c7x6 & K3c7x6);
assign K3c7x6 = (~(Pvb7x6 & Cmm7z6[22]));
assign Pvb7x6 = (~(Wvb7x6 | Uub7x6));
assign D3c7x6 = (~(Wvb7x6 & Wui7z6[22]));
assign Wvb7x6 = (~(Uub7x6 | Hkb7x6));
assign Uub7x6 = (R3c7x6 & Bqi7z6[2]);
assign R3c7x6 = (!Okb7x6);
assign H1y7v6 = (~(Y3c7x6 & F4c7x6));
assign F4c7x6 = (~(M4c7x6 & X0hov6));
assign Y3c7x6 = (T4c7x6 & A5c7x6);
assign A5c7x6 = (~(H5c7x6 & Cmm7z6[31]));
assign T4c7x6 = (~(O5c7x6 & Wui7z6[31]));
assign A1y7v6 = (~(V5c7x6 & C6c7x6));
assign C6c7x6 = (~(M4c7x6 & Wf4iw6));
assign V5c7x6 = (J6c7x6 & Q6c7x6);
assign Q6c7x6 = (~(H5c7x6 & Cmm7z6[24]));
assign J6c7x6 = (~(O5c7x6 & Wui7z6[24]));
assign T0y7v6 = (~(X6c7x6 & E7c7x6));
assign E7c7x6 = (~(M4c7x6 & Iklov6));
assign X6c7x6 = (L7c7x6 & S7c7x6);
assign S7c7x6 = (~(H5c7x6 & Cmm7z6[25]));
assign L7c7x6 = (~(O5c7x6 & Wui7z6[25]));
assign M0y7v6 = (~(Z7c7x6 & G8c7x6));
assign G8c7x6 = (~(M4c7x6 & E64iw6));
assign Z7c7x6 = (N8c7x6 & U8c7x6);
assign U8c7x6 = (~(H5c7x6 & Cmm7z6[26]));
assign N8c7x6 = (~(O5c7x6 & Wui7z6[26]));
assign F0y7v6 = (~(B9c7x6 & I9c7x6));
assign I9c7x6 = (~(M4c7x6 & H44iw6));
assign B9c7x6 = (P9c7x6 & W9c7x6);
assign W9c7x6 = (~(H5c7x6 & Cmm7z6[27]));
assign P9c7x6 = (~(O5c7x6 & Wui7z6[27]));
assign Yzx7v6 = (~(Dac7x6 & Kac7x6));
assign Kac7x6 = (~(M4c7x6 & W14iw6));
assign Dac7x6 = (Rac7x6 & Yac7x6);
assign Yac7x6 = (~(H5c7x6 & Cmm7z6[28]));
assign Rac7x6 = (~(O5c7x6 & Wui7z6[28]));
assign Rzx7v6 = (~(Fbc7x6 & Mbc7x6));
assign Mbc7x6 = (~(M4c7x6 & Zz3iw6));
assign Fbc7x6 = (Tbc7x6 & Acc7x6);
assign Acc7x6 = (~(H5c7x6 & Cmm7z6[29]));
assign Tbc7x6 = (~(O5c7x6 & Wui7z6[29]));
assign Kzx7v6 = (~(Hcc7x6 & Occ7x6));
assign Occ7x6 = (~(M4c7x6 & Ro3iw6));
assign Hcc7x6 = (Vcc7x6 & Cdc7x6);
assign Cdc7x6 = (~(H5c7x6 & Cmm7z6[30]));
assign H5c7x6 = (~(O5c7x6 | M4c7x6));
assign Vcc7x6 = (~(O5c7x6 & Wui7z6[30]));
assign O5c7x6 = (~(Hkb7x6 | M4c7x6));
assign M4c7x6 = (~(Okb7x6 | Dv3iw6));
assign Okb7x6 = (~(Jdc7x6 & Qdc7x6));
assign Qdc7x6 = (Xdc7x6 & G92iw6);
assign Xdc7x6 = (~(Toi7z6[3] & Toi7z6[2]));
assign Jdc7x6 = (Eec7x6 & Toi7z6[4]);
assign Hkb7x6 = (Lec7x6 & Sec7x6);
assign Sec7x6 = (~(Zec7x6 | A8y7v6));
assign A8y7v6 = (~(M697z6 & Gfc7x6));
assign Gfc7x6 = (~(Bzi7z6[7] & Nfc7x6));
assign Nfc7x6 = (~(P3b7x6 & O87iw6));
assign Zec7x6 = (Q9y7v6 | Ihnet6);
assign Q9y7v6 = (~(N9b7x6 & Ufc7x6));
assign Ufc7x6 = (~(Bzi7z6[15] & Bgc7x6));
assign Bgc7x6 = (~(P3b7x6 & Hv5iw6));
assign N9b7x6 = (!Tlb7z6[1]);
assign Lec7x6 = (Vfmov6 & Qvkiw6);
assign Dzx7v6 = (~(Gd77z6 & Igc7x6));
assign Igc7x6 = (~(Bzi7z6[4] & Pgc7x6));
assign Pgc7x6 = (~(Z1b7x6 & W52nv6));
assign Wyx7v6 = (~(Sosiw6 & Wgc7x6));
assign Wgc7x6 = (~(Bzi7z6[3] & Dhc7x6));
assign Dhc7x6 = (~(Z1b7x6 & P52nv6));
assign Pyx7v6 = (~(M697z6 & Khc7x6));
assign Khc7x6 = (~(Bzi7z6[1] & Rhc7x6));
assign Rhc7x6 = (~(Z1b7x6 & B52nv6));
assign Z1b7x6 = (P3b7x6 & Bqi7z6[0]);
assign P3b7x6 = (Yhc7x6 & T68iw6);
assign Iyx7v6 = (~(Fic7x6 & Mic7x6));
assign Mic7x6 = (~(Tic7x6 & Snvnv6));
assign Snvnv6 = (B8cdt6 & N3onv6);
assign Tic7x6 = (Ajc7x6 & Hjc7x6);
assign Hjc7x6 = (~(Tltov6 & Ojc7x6));
assign Ojc7x6 = (~(G5sov6 & Xeinv6));
assign Tltov6 = (Vjc7x6 & Ckc7x6);
assign Ckc7x6 = (~(Auehw6 & Q8onv6));
assign Vjc7x6 = (Jkc7x6 & Yvihw6);
assign Yvihw6 = (!Qkc7x6);
assign Ajc7x6 = (~(J2cdt6 & Ga3nv6));
assign Fic7x6 = (~(Bqbdt6 & Dcnov6));
assign Byx7v6 = (Pb9ov6 ? D6c7z6[4] : Xkc7x6);
assign Xkc7x6 = (~(Elc7x6 & Llc7x6));
assign Llc7x6 = (Slc7x6 & Zlc7x6);
assign Zlc7x6 = (~(Yc9ov6 & T977x6));
assign Slc7x6 = (~(Md9ov6 & Cb77x6));
assign Elc7x6 = (Gmc7x6 & Nmc7x6);
assign Nmc7x6 = (~(Oe9ov6 & Ax57x6));
assign Gmc7x6 = (~(Cf9ov6 & Tw57x6));
assign Uxx7v6 = (Pb9ov6 ? D6c7z6[1] : Umc7x6);
assign Pb9ov6 = (~(J7l8v6 | Cubdt6));
assign J7l8v6 = (Bnc7x6 & Inc7x6);
assign Inc7x6 = (Pnc7x6 & Wnc7x6);
assign Wnc7x6 = (Doc7x6 & Koc7x6);
assign Koc7x6 = (Hp67x6 & Bfo7v6);
assign Doc7x6 = (Nm57x6 & Dh57x6);
assign Pnc7x6 = (Roc7x6 & C477x6);
assign Roc7x6 = (Qr57x6 & Cx67x6);
assign Bnc7x6 = (Yoc7x6 & Fpc7x6);
assign Fpc7x6 = (Mpc7x6 & Tpc7x6);
assign Tpc7x6 = (~(Aqc7x6 & Hqc7x6));
assign Hqc7x6 = (~(Oqc7x6 & Vqc7x6));
assign Vqc7x6 = (Crc7x6 & Hnlov6);
assign Crc7x6 = (Ob67x6 & Ve9ov6);
assign Oqc7x6 = (Jrc7x6 & Ddfov6);
assign Jrc7x6 = (~(Qrc7x6 & Xrc7x6));
assign Xrc7x6 = (~(Esc7x6 & Lsc7x6));
assign Lsc7x6 = (Yc9ov6 & Ssc7x6);
assign Esc7x6 = (Zsc7x6 & Gtc7x6);
assign Qrc7x6 = (~(Ntc7x6 & Utc7x6));
assign Utc7x6 = (~(Buc7x6 & Iuc7x6));
assign Iuc7x6 = (~(Ssc7x6 & Cf9ov6));
assign Buc7x6 = (~(Gtc7x6 & Md9ov6));
assign Aqc7x6 = (~(Puc7x6 & Wuc7x6));
assign Wuc7x6 = (Oe9ov6 & Ssc7x6);
assign Ssc7x6 = (Dvc7x6 & Kvc7x6);
assign Kvc7x6 = (Td9ov6 & Icfov6);
assign Dvc7x6 = (Mmlov6 & Ex77x6);
assign Puc7x6 = (Ntc7x6 & Gtc7x6);
assign Gtc7x6 = (Rvc7x6 & Yvc7x6);
assign Yvc7x6 = (Ab67x6 & Jf9ov6);
assign Rvc7x6 = (Kdfov6 & Onlov6);
assign Ntc7x6 = (Fwc7x6 & Mwc7x6);
assign Mwc7x6 = (Twc7x6 & Vv77x6);
assign Twc7x6 = (Fd9ov6 & Bcfov6);
assign Fwc7x6 = (Zsc7x6 & Fmlov6);
assign Zsc7x6 = (Axc7x6 & Hxc7x6);
assign Hxc7x6 = (Oxc7x6 & Vxc7x6);
assign Vxc7x6 = (Kn67x6 & Rh57x6);
assign Oxc7x6 = (Um57x6 & Tv67x6);
assign Axc7x6 = (Cyc7x6 & Jyc7x6);
assign Jyc7x6 = (Xr57x6 & T277x6);
assign Cyc7x6 = (Ax57x6 & T977x6);
assign Mpc7x6 = (Cb77x6 & Tw57x6);
assign Yoc7x6 = (Qyc7x6 & Bqbdt6);
assign Qyc7x6 = (O5a7z6 & Xyc7x6);
assign Xyc7x6 = (~(Ezc7x6 & Lzc7x6));
assign Lzc7x6 = (Szc7x6 | Twphw6);
assign Ezc7x6 = (Zzc7x6 & G0d7x6);
assign G0d7x6 = (~(N0d7x6 & J8a7x6));
assign N0d7x6 = (Ntg7z6[1] & U0d7x6);
assign U0d7x6 = (~(B1d7x6 & I1d7x6));
assign B1d7x6 = (~(P1d7x6 & W1d7x6));
assign W1d7x6 = (~(I0c7z6[0] | Zdxdt6));
assign P1d7x6 = (I0c7z6[1] & D2d7x6);
assign D2d7x6 = (~(K2d7x6 & I3wnv6));
assign Zzc7x6 = (~(R2d7x6 & V7a7x6));
assign V7a7x6 = (Y2d7x6 & Pxg7z6[3]);
assign Y2d7x6 = (Pxg7z6[2] & Pxg7z6[0]);
assign R2d7x6 = (Ot97x6 & Pxg7z6[1]);
assign Umc7x6 = (~(F3d7x6 & M3d7x6));
assign M3d7x6 = (T3d7x6 & A4d7x6);
assign A4d7x6 = (~(Yc9ov6 & Vv77x6));
assign T3d7x6 = (~(Md9ov6 & Ex77x6));
assign F3d7x6 = (H4d7x6 & O4d7x6);
assign O4d7x6 = (~(Oe9ov6 & Ob67x6));
assign H4d7x6 = (~(Cf9ov6 & Ab67x6));
assign Nxx7v6 = (V4d7x6 | C5d7x6);
assign V4d7x6 = (J5d7x6 | Q5d7x6);
assign J5d7x6 = (X5d7x6 & Uyb7z6[0]);
assign Gxx7v6 = (~(E6d7x6 & L6d7x6));
assign L6d7x6 = (~(X5d7x6 & Uyb7z6[1]));
assign Zwx7v6 = (~(S6d7x6 & Ad9iw6));
assign S6d7x6 = (Z6d7x6 & G7d7x6);
assign G7d7x6 = (~(N7d7x6 & Q5d7x6));
assign N7d7x6 = (J2cdt6 & Jjbdt6);
assign Z6d7x6 = (~(X5d7x6 & Uyb7z6[2]));
assign Swx7v6 = (~(U7d7x6 & Qolov6));
assign U7d7x6 = (B8d7x6 & I8d7x6);
assign I8d7x6 = (~(Q5d7x6 & J2cdt6));
assign B8d7x6 = (~(X5d7x6 & Uyb7z6[3]));
assign Lwx7v6 = (~(P8d7x6 & W8d7x6));
assign W8d7x6 = (~(Q5d7x6 | D9d7x6));
assign Q5d7x6 = (~(K9d7x6 | X5d7x6));
assign P8d7x6 = (R9d7x6 & Y9d7x6);
assign Y9d7x6 = (~(X5d7x6 & Uyb7z6[4]));
assign X5d7x6 = (Q0wnv6 & Kkmhw6);
assign R9d7x6 = (~(D6c7z6[4] & Cubdt6));
assign Xvx7v6 = (Ad2iw6 & Bu4ov6);
assign Qvx7v6 = (Ut4ov6 ? Fad7x6 : Zas7z6[0]);
assign Jvx7v6 = (Ut4ov6 ? A62iw6 : Zfs7z6[11]);
assign Cvx7v6 = (Ut4ov6 ? O62iw6 : Zfs7z6[10]);
assign Vux7v6 = (Ut4ov6 ? V62iw6 : Zfs7z6[9]);
assign Oux7v6 = (Ut4ov6 ? C72iw6 : Zfs7z6[8]);
assign Hux7v6 = (Ut4ov6 ? J72iw6 : Zfs7z6[7]);
assign Aux7v6 = (Ut4ov6 ? Q72iw6 : Mm27v6);
assign Q72iw6 = (~(Mad7x6 & Tad7x6));
assign Tad7x6 = (~(Fvb7z6[6] & M52iw6));
assign Mad7x6 = (~(Se3iw6 & Cmm7z6[6]));
assign Ttx7v6 = (Ut4ov6 ? X72iw6 : Tn27v6);
assign Ut4ov6 = (!Abd7x6);
assign X72iw6 = (~(Hbd7x6 & Obd7x6));
assign Obd7x6 = (~(Fvb7z6[5] & M52iw6));
assign Hbd7x6 = (~(Se3iw6 & Cmm7z6[5]));
assign Mtx7v6 = (Abd7x6 ? Ap27v6 : E82iw6);
assign E82iw6 = (~(Vbd7x6 & Ccd7x6));
assign Ccd7x6 = (~(Fvb7z6[4] & M52iw6));
assign Vbd7x6 = (~(Se3iw6 & Cmm7z6[4]));
assign Ftx7v6 = (Abd7x6 ? Hq27v6 : L82iw6);
assign L82iw6 = (~(Jcd7x6 & Qcd7x6));
assign Qcd7x6 = (~(Fvb7z6[3] & M52iw6));
assign Jcd7x6 = (~(Se3iw6 & Cmm7z6[3]));
assign Ysx7v6 = (Abd7x6 ? Or27v6 : S82iw6);
assign S82iw6 = (~(Xcd7x6 & Edd7x6));
assign Edd7x6 = (~(Se3iw6 & Yefnv6));
assign Xcd7x6 = (~(Fvb7z6[2] & M52iw6));
assign Wrx7v6 = (~(Ldd7x6 & Sdd7x6));
assign Sdd7x6 = (~(Iqeiw6 & Zdd7x6));
assign Zdd7x6 = (~(Ged7x6 & Ned7x6));
assign Ned7x6 = (~(Rsx7v6 | Ewx7v6));
assign Ewx7v6 = (Ued7x6 & Ujlov6);
assign Ujlov6 = (~(Bfd7x6 & Ifd7x6));
assign Ifd7x6 = (Pfd7x6 | Wfd7x6);
assign Rsx7v6 = (Ued7x6 & Pa2iw6);
assign Pa2iw6 = (~(Bfd7x6 & Dgd7x6));
assign Dgd7x6 = (Kgd7x6 | G83iw6);
assign Ged7x6 = (~(Dsx7v6 | Ksx7v6));
assign Ksx7v6 = (Ued7x6 & Kb2iw6);
assign Kb2iw6 = (~(Bfd7x6 & Rgd7x6));
assign Rgd7x6 = (Wfd7x6 | G83iw6);
assign G83iw6 = (!Pfd7x6);
assign Wfd7x6 = (Ygd7x6 & Fhd7x6);
assign Fhd7x6 = (~(N83iw6 & Fad7x6));
assign Dsx7v6 = (Ued7x6 & Fc2iw6);
assign Fc2iw6 = (~(Bfd7x6 & Mhd7x6));
assign Mhd7x6 = (Pfd7x6 | Kgd7x6);
assign Kgd7x6 = (Ygd7x6 & Thd7x6);
assign Thd7x6 = (Aid7x6 | N83iw6);
assign N83iw6 = (Hid7x6 & Oid7x6);
assign Oid7x6 = (~(M52iw6 & Mbqnv6));
assign Hid7x6 = (~(Se3iw6 & Cmm7z6[0]));
assign Pfd7x6 = (~(Vid7x6 & Cjd7x6));
assign Cjd7x6 = (~(M52iw6 & Stpnv6));
assign Vid7x6 = (~(Se3iw6 & Cmm7z6[1]));
assign Ued7x6 = (~(Jjd7x6 | Ad2iw6));
assign Ad2iw6 = (!D42iw6);
assign D42iw6 = (~(Qjd7x6 & Xjd7x6));
assign Xjd7x6 = (~(Se3iw6 & Lhmov6));
assign Qjd7x6 = (~(L3bdt6 & M52iw6));
assign Iqeiw6 = (Ekd7x6 & Lkd7x6);
assign Lkd7x6 = (~(Skd7x6 | C72iw6));
assign C72iw6 = (~(Zkd7x6 & Gld7x6));
assign Gld7x6 = (~(Fvb7z6[8] & M52iw6));
assign Zkd7x6 = (~(Se3iw6 & Cmm7z6[8]));
assign Skd7x6 = (J72iw6 | V62iw6);
assign V62iw6 = (~(Nld7x6 & Uld7x6));
assign Uld7x6 = (~(Fvb7z6[9] & M52iw6));
assign Nld7x6 = (~(Se3iw6 & Cmm7z6[9]));
assign J72iw6 = (~(Bmd7x6 & Imd7x6));
assign Imd7x6 = (~(Fvb7z6[7] & M52iw6));
assign Bmd7x6 = (~(Se3iw6 & Cmm7z6[7]));
assign Ekd7x6 = (~(O62iw6 | A62iw6));
assign A62iw6 = (~(Pmd7x6 & Wmd7x6));
assign Wmd7x6 = (~(Fvb7z6[11] & M52iw6));
assign Pmd7x6 = (~(Se3iw6 & Cmm7z6[11]));
assign O62iw6 = (~(Dnd7x6 & Knd7x6));
assign Knd7x6 = (~(Fvb7z6[10] & M52iw6));
assign Dnd7x6 = (~(Se3iw6 & Cmm7z6[10]));
assign Ldd7x6 = (~(Ci27v6 & Abd7x6));
assign Prx7v6 = (Abd7x6 ? Zas7z6[1] : Rnd7x6);
assign Abd7x6 = (Ynd7x6 & Fod7x6);
assign Fod7x6 = (~(Mod7x6 | Ihs7z6[1]));
assign Mod7x6 = (Ihs7z6[2] | Ihs7z6[3]);
assign Ynd7x6 = (Tod7x6 & Jjd7x6);
assign Jjd7x6 = (!Bu4ov6);
assign Bu4ov6 = (Apd7x6 & Ofeiw6);
assign Ofeiw6 = (Hpd7x6 & Opd7x6);
assign Hpd7x6 = (Rkeiw6 & Oteiw6);
assign Rkeiw6 = (!Jrhiw6);
assign Apd7x6 = (~(C63iw6 | Kygnv6));
assign Tod7x6 = (Cch7v6 & Vpd7x6);
assign Rnd7x6 = (~(Bfd7x6 & Ygd7x6));
assign Ygd7x6 = (~(Cqd7x6 & Jqd7x6));
assign Cqd7x6 = (Qqd7x6 & Aid7x6);
assign Bfd7x6 = (Aid7x6 | Xqd7x6);
assign Xqd7x6 = (Jqd7x6 & Qqd7x6);
assign Qqd7x6 = (~(Se3iw6 & Anehw6));
assign Jqd7x6 = (~(M52iw6 & Hub7z6[1]));
assign Aid7x6 = (!Fad7x6);
assign Fad7x6 = (Erd7x6 & Lrd7x6);
assign Lrd7x6 = (~(M52iw6 & Hub7z6[0]));
assign Erd7x6 = (~(Se3iw6 & Wbhnv6));
assign Irx7v6 = (~(Srd7x6 & Zrd7x6));
assign Zrd7x6 = (~(Dpwnv6 & Itb7z6[1]));
assign Srd7x6 = (Gsd7x6 & Nsd7x6);
assign Nsd7x6 = (~(Usd7x6 & Fqwnv6));
assign Usd7x6 = (~(Btd7x6 & Itd7x6));
assign Itd7x6 = (Ptd7x6 & Wtd7x6);
assign Wtd7x6 = (Wawnv6 | Dud7x6);
assign Ptd7x6 = (~(Dtm7z6[3] & Kud7x6));
assign Btd7x6 = (Rud7x6 & Yud7x6);
assign Yud7x6 = (~(Dtm7z6[0] & HRDATAD[1]));
assign Rud7x6 = (~(Dtm7z6[1] & HRDATAS[1]));
assign Gsd7x6 = (~(Qvzhw6 & Fvd7x6));
assign Qvzhw6 = (!Jvzhw6);
assign Jvzhw6 = (~(Dbymz6[0] & Cbyhw6));
assign Cbyhw6 = (JTAGNSW ? Aixmz6[1] : Ulxmz6[1]);
assign Brx7v6 = (~(Mvd7x6 & Tvd7x6));
assign Tvd7x6 = (~(Dpwnv6 & Itb7z6[2]));
assign Mvd7x6 = (Awd7x6 & Hwd7x6);
assign Hwd7x6 = (~(Owd7x6 & Fqwnv6));
assign Owd7x6 = (~(Vwd7x6 & Cxd7x6));
assign Cxd7x6 = (Jxd7x6 & Qxd7x6);
assign Qxd7x6 = (Wawnv6 | Xxd7x6);
assign Jxd7x6 = (~(Dtm7z6[3] & Eyd7x6));
assign Vwd7x6 = (Lyd7x6 & Syd7x6);
assign Syd7x6 = (~(Dtm7z6[0] & HRDATAD[2]));
assign Lyd7x6 = (~(Dtm7z6[1] & HRDATAS[2]));
assign Awd7x6 = (~(Fcwnv6 & P7yhw6));
assign P7yhw6 = (Dz1nv6 ? Ulxmz6[2] : Aixmz6[2]);
assign Uqx7v6 = (~(Zyd7x6 & Gzd7x6));
assign Gzd7x6 = (~(Dpwnv6 & Itb7z6[3]));
assign Zyd7x6 = (Nzd7x6 & Uzd7x6);
assign Uzd7x6 = (~(B0e7x6 & Fqwnv6));
assign B0e7x6 = (~(I0e7x6 & P0e7x6));
assign P0e7x6 = (W0e7x6 & D1e7x6);
assign D1e7x6 = (Wawnv6 | K1e7x6);
assign W0e7x6 = (~(Dtm7z6[3] & R1e7x6));
assign I0e7x6 = (Y1e7x6 & F2e7x6);
assign F2e7x6 = (~(Dtm7z6[0] & HRDATAD[3]));
assign Y1e7x6 = (~(Dtm7z6[1] & HRDATAS[3]));
assign Nzd7x6 = (~(Fcwnv6 & Z5yhw6));
assign Z5yhw6 = (Dz1nv6 ? Ulxmz6[3] : Aixmz6[3]);
assign Nqx7v6 = (~(M2e7x6 & T2e7x6));
assign T2e7x6 = (~(Dpwnv6 & Itb7z6[4]));
assign M2e7x6 = (A3e7x6 & H3e7x6);
assign H3e7x6 = (~(O3e7x6 & Fqwnv6));
assign O3e7x6 = (~(V3e7x6 & C4e7x6));
assign C4e7x6 = (J4e7x6 & Q4e7x6);
assign Q4e7x6 = (Wawnv6 | X4e7x6);
assign J4e7x6 = (~(Dtm7z6[3] & E5e7x6));
assign V3e7x6 = (L5e7x6 & S5e7x6);
assign S5e7x6 = (~(Dtm7z6[0] & HRDATAD[4]));
assign L5e7x6 = (~(Dtm7z6[1] & HRDATAS[4]));
assign A3e7x6 = (~(Fcwnv6 & Q20iw6));
assign Q20iw6 = (JTAGNSW ? Aixmz6[4] : Ulxmz6[4]);
assign Gqx7v6 = (~(Z5e7x6 & G6e7x6));
assign G6e7x6 = (~(Dpwnv6 & Itb7z6[5]));
assign Z5e7x6 = (N6e7x6 & U6e7x6);
assign U6e7x6 = (~(B7e7x6 & Fqwnv6));
assign B7e7x6 = (~(I7e7x6 & P7e7x6));
assign P7e7x6 = (W7e7x6 & D8e7x6);
assign D8e7x6 = (Wawnv6 | K8e7x6);
assign W7e7x6 = (~(Dtm7z6[3] & R8e7x6));
assign I7e7x6 = (Y8e7x6 & F9e7x6);
assign F9e7x6 = (~(Dtm7z6[0] & HRDATAD[5]));
assign Y8e7x6 = (~(Dtm7z6[1] & HRDATAS[5]));
assign N6e7x6 = (~(Rszhw6 & Fvd7x6));
assign Rszhw6 = (Dbymz6[0] & L5yhw6);
assign L5yhw6 = (JTAGNSW ? Aixmz6[5] : Ulxmz6[5]);
assign Zpx7v6 = (~(M9e7x6 & T9e7x6));
assign T9e7x6 = (~(Dpwnv6 & Itb7z6[6]));
assign M9e7x6 = (Aae7x6 & Hae7x6);
assign Hae7x6 = (~(Oae7x6 & Fqwnv6));
assign Oae7x6 = (~(Vae7x6 & Cbe7x6));
assign Cbe7x6 = (Jbe7x6 & Qbe7x6);
assign Qbe7x6 = (Wawnv6 | Xbe7x6);
assign Jbe7x6 = (~(Dtm7z6[3] & Ece7x6));
assign Vae7x6 = (Lce7x6 & Sce7x6);
assign Sce7x6 = (~(Dtm7z6[0] & HRDATAD[6]));
assign Lce7x6 = (~(Dtm7z6[1] & HRDATAS[6]));
assign Aae7x6 = (~(Fcwnv6 & F9yhw6));
assign F9yhw6 = (Dz1nv6 ? Ulxmz6[6] : Aixmz6[6]);
assign Spx7v6 = (~(Zce7x6 & Gde7x6));
assign Gde7x6 = (~(Fcwnv6 & B7yhw6));
assign B7yhw6 = (Dz1nv6 ? Ulxmz6[7] : Aixmz6[7]);
assign Zce7x6 = (Nde7x6 & Ude7x6);
assign Ude7x6 = (~(Bee7x6 & Fqwnv6));
assign Bee7x6 = (~(Iee7x6 & Pee7x6));
assign Pee7x6 = (Wee7x6 & Dfe7x6);
assign Dfe7x6 = (Wawnv6 | Kfe7x6);
assign Wee7x6 = (~(Dtm7z6[3] & Rfe7x6));
assign Iee7x6 = (Yfe7x6 & Fge7x6);
assign Fge7x6 = (~(Dtm7z6[0] & HRDATAD[7]));
assign Yfe7x6 = (~(Dtm7z6[1] & HRDATAS[7]));
assign Nde7x6 = (~(Dpwnv6 & Itb7z6[7]));
assign Dpwnv6 = (~(Fqwnv6 | Fvd7x6));
assign Fqwnv6 = (~(Mge7x6 & Tge7x6));
assign Tge7x6 = (~(Ahe7x6 & Hhe7x6));
assign Hhe7x6 = (~(Ohe7x6 & Vhe7x6));
assign Vhe7x6 = (~(Cie7x6 & Jie7x6));
assign Cie7x6 = (Qie7x6 & Xie7x6);
assign Mge7x6 = (Eje7x6 | Xie7x6);
assign Lpx7v6 = (~(Lje7x6 & Sje7x6));
assign Sje7x6 = (~(Zje7x6 & Itb7z6[9]));
assign Lje7x6 = (Gke7x6 & Nke7x6);
assign Nke7x6 = (~(Uke7x6 & Ble7x6));
assign Ble7x6 = (~(Ile7x6 & Ple7x6));
assign Ple7x6 = (Wle7x6 & Dme7x6);
assign Dme7x6 = (Wawnv6 | Kme7x6);
assign Wle7x6 = (~(Dtm7z6[3] & Rme7x6));
assign Ile7x6 = (Yme7x6 & Fne7x6);
assign Fne7x6 = (~(Dtm7z6[0] & HRDATAD[9]));
assign Yme7x6 = (~(Dtm7z6[1] & HRDATAS[9]));
assign Gke7x6 = (~(Fcwnv6 & R0zhw6));
assign R0zhw6 = (Dz1nv6 ? Ulxmz6[9] : Aixmz6[9]);
assign Epx7v6 = (~(Mne7x6 & Tne7x6));
assign Tne7x6 = (~(Zje7x6 & Itb7z6[10]));
assign Mne7x6 = (Aoe7x6 & Hoe7x6);
assign Hoe7x6 = (~(Uke7x6 & Ooe7x6));
assign Ooe7x6 = (~(Voe7x6 & Cpe7x6));
assign Cpe7x6 = (Jpe7x6 & Qpe7x6);
assign Qpe7x6 = (Wawnv6 | Xpe7x6);
assign Jpe7x6 = (~(Dtm7z6[3] & Eqe7x6));
assign Voe7x6 = (Lqe7x6 & Sqe7x6);
assign Sqe7x6 = (~(Dtm7z6[0] & HRDATAD[10]));
assign Lqe7x6 = (~(Dtm7z6[1] & HRDATAS[10]));
assign Aoe7x6 = (~(Fcwnv6 & Lxyhw6));
assign Lxyhw6 = (Dz1nv6 ? Ulxmz6[10] : Aixmz6[10]);
assign Xox7v6 = (~(Zqe7x6 & Gre7x6));
assign Gre7x6 = (~(Zje7x6 & Itb7z6[11]));
assign Zqe7x6 = (Nre7x6 & Ure7x6);
assign Ure7x6 = (~(Uke7x6 & Bse7x6));
assign Bse7x6 = (~(Ise7x6 & Pse7x6));
assign Pse7x6 = (Wse7x6 & Dte7x6);
assign Dte7x6 = (Wawnv6 | Kte7x6);
assign Wse7x6 = (~(Dtm7z6[3] & Rte7x6));
assign Ise7x6 = (Yte7x6 & Fue7x6);
assign Fue7x6 = (~(Dtm7z6[0] & HRDATAD[11]));
assign Yte7x6 = (~(Dtm7z6[1] & HRDATAS[11]));
assign Nre7x6 = (~(Fcwnv6 & Vvyhw6));
assign Vvyhw6 = (Dz1nv6 ? Ulxmz6[11] : Aixmz6[11]);
assign Qox7v6 = (~(Mue7x6 & Tue7x6));
assign Tue7x6 = (~(Zje7x6 & Itb7z6[12]));
assign Mue7x6 = (Ave7x6 & Hve7x6);
assign Hve7x6 = (~(Uke7x6 & Ove7x6));
assign Ove7x6 = (~(Vve7x6 & Cwe7x6));
assign Cwe7x6 = (Jwe7x6 & Qwe7x6);
assign Qwe7x6 = (Wawnv6 | Xwe7x6);
assign Jwe7x6 = (~(Dtm7z6[3] & Exe7x6));
assign Vve7x6 = (Lxe7x6 & Sxe7x6);
assign Sxe7x6 = (~(Dtm7z6[0] & HRDATAD[12]));
assign Lxe7x6 = (~(Dtm7z6[1] & HRDATAS[12]));
assign Ave7x6 = (~(Fcwnv6 & Bzyhw6));
assign Bzyhw6 = (JTAGNSW ? Aixmz6[12] : Ulxmz6[12]);
assign Jox7v6 = (~(Zxe7x6 & Gye7x6));
assign Gye7x6 = (~(Zje7x6 & Itb7z6[13]));
assign Zxe7x6 = (Nye7x6 & Uye7x6);
assign Uye7x6 = (~(Uke7x6 & Bze7x6));
assign Bze7x6 = (~(Ize7x6 & Pze7x6));
assign Pze7x6 = (Wze7x6 & D0f7x6);
assign D0f7x6 = (Wawnv6 | K0f7x6);
assign Wze7x6 = (~(Dtm7z6[3] & R0f7x6));
assign Ize7x6 = (Y0f7x6 & F1f7x6);
assign F1f7x6 = (~(Dtm7z6[0] & HRDATAD[13]));
assign Y0f7x6 = (~(Dtm7z6[1] & HRDATAS[13]));
assign Nye7x6 = (~(Fcwnv6 & Hvyhw6));
assign Hvyhw6 = (JTAGNSW ? Aixmz6[13] : Ulxmz6[13]);
assign Cox7v6 = (~(M1f7x6 & T1f7x6));
assign T1f7x6 = (~(Zje7x6 & Itb7z6[14]));
assign M1f7x6 = (A2f7x6 & H2f7x6);
assign H2f7x6 = (~(Uke7x6 & O2f7x6));
assign O2f7x6 = (~(V2f7x6 & C3f7x6));
assign C3f7x6 = (J3f7x6 & Q3f7x6);
assign Q3f7x6 = (Wawnv6 | X3f7x6);
assign J3f7x6 = (~(Dtm7z6[3] & E4f7x6));
assign V2f7x6 = (L4f7x6 & S4f7x6);
assign S4f7x6 = (~(Dtm7z6[0] & HRDATAD[14]));
assign L4f7x6 = (~(Dtm7z6[1] & HRDATAS[14]));
assign A2f7x6 = (~(Fcwnv6 & Pzyhw6));
assign Pzyhw6 = (JTAGNSW ? Aixmz6[14] : Ulxmz6[14]);
assign Vnx7v6 = (~(Z4f7x6 & G5f7x6));
assign G5f7x6 = (~(Zje7x6 & Itb7z6[15]));
assign Z4f7x6 = (N5f7x6 & U5f7x6);
assign U5f7x6 = (~(Uke7x6 & B6f7x6));
assign B6f7x6 = (~(I6f7x6 & P6f7x6));
assign P6f7x6 = (W6f7x6 & D7f7x6);
assign D7f7x6 = (Wawnv6 | K7f7x6);
assign W6f7x6 = (~(Dtm7z6[3] & R7f7x6));
assign I6f7x6 = (Y7f7x6 & F8f7x6);
assign F8f7x6 = (~(Dtm7z6[0] & HRDATAD[15]));
assign Y7f7x6 = (~(Dtm7z6[1] & HRDATAS[15]));
assign N5f7x6 = (~(Fcwnv6 & Xwyhw6));
assign Xwyhw6 = (JTAGNSW ? Aixmz6[15] : Ulxmz6[15]);
assign Onx7v6 = (~(M8f7x6 & T8f7x6));
assign T8f7x6 = (~(Fcwnv6 & F1zhw6));
assign F1zhw6 = (Dz1nv6 ? Ulxmz6[8] : Aixmz6[8]);
assign M8f7x6 = (A9f7x6 & H9f7x6);
assign H9f7x6 = (~(Uke7x6 & O9f7x6));
assign O9f7x6 = (~(V9f7x6 & Caf7x6));
assign Caf7x6 = (Jaf7x6 & Qaf7x6);
assign Qaf7x6 = (Wawnv6 | Xaf7x6);
assign Jaf7x6 = (~(Dtm7z6[3] & Ebf7x6));
assign V9f7x6 = (Lbf7x6 & Sbf7x6);
assign Sbf7x6 = (~(Dtm7z6[0] & HRDATAD[8]));
assign Lbf7x6 = (~(Dtm7z6[1] & HRDATAS[8]));
assign A9f7x6 = (~(Zje7x6 & Itb7z6[8]));
assign Zje7x6 = (~(Fvd7x6 | Uke7x6));
assign Uke7x6 = (Ahe7x6 & Zbf7x6);
assign Zbf7x6 = (~(Ohe7x6 & Gcf7x6));
assign Gcf7x6 = (~(Ncf7x6 & Xie7x6));
assign Hnx7v6 = (~(Ucf7x6 & Bdf7x6));
assign Bdf7x6 = (~(Idf7x6 & Itb7z6[17]));
assign Ucf7x6 = (Pdf7x6 & Wdf7x6);
assign Wdf7x6 = (~(Def7x6 & Kef7x6));
assign Def7x6 = (~(Ref7x6 & Yef7x6));
assign Yef7x6 = (Fff7x6 & Mff7x6);
assign Mff7x6 = (Wawnv6 | Tff7x6);
assign Fff7x6 = (~(Dtm7z6[3] & Agf7x6));
assign Ref7x6 = (Hgf7x6 & Ogf7x6);
assign Ogf7x6 = (~(Dtm7z6[0] & HRDATAD[17]));
assign Hgf7x6 = (~(Dtm7z6[1] & HRDATAS[17]));
assign Pdf7x6 = (~(Fcwnv6 & Ejyhw6));
assign Ejyhw6 = (JTAGNSW ? Aixmz6[17] : Ulxmz6[17]);
assign Anx7v6 = (~(Vgf7x6 & Chf7x6));
assign Chf7x6 = (~(Idf7x6 & Itb7z6[18]));
assign Vgf7x6 = (Jhf7x6 & Qhf7x6);
assign Qhf7x6 = (~(Xhf7x6 & Kef7x6));
assign Xhf7x6 = (~(Eif7x6 & Lif7x6));
assign Lif7x6 = (Sif7x6 & Zif7x6);
assign Zif7x6 = (Wawnv6 | Gjf7x6);
assign Sif7x6 = (~(Dtm7z6[3] & Njf7x6));
assign Eif7x6 = (Ujf7x6 & Bkf7x6);
assign Bkf7x6 = (~(Dtm7z6[0] & HRDATAD[18]));
assign Ujf7x6 = (~(Dtm7z6[1] & HRDATAS[18]));
assign Jhf7x6 = (~(Fcwnv6 & Yfyhw6));
assign Yfyhw6 = (JTAGNSW ? Aixmz6[18] : Ulxmz6[18]);
assign Tmx7v6 = (~(Ikf7x6 & Pkf7x6));
assign Pkf7x6 = (~(Idf7x6 & Itb7z6[19]));
assign Ikf7x6 = (Wkf7x6 & Dlf7x6);
assign Dlf7x6 = (~(Klf7x6 & Kef7x6));
assign Klf7x6 = (~(Rlf7x6 & Ylf7x6));
assign Ylf7x6 = (Fmf7x6 & Mmf7x6);
assign Mmf7x6 = (Wawnv6 | Tmf7x6);
assign Fmf7x6 = (~(Dtm7z6[3] & Anf7x6));
assign Rlf7x6 = (Hnf7x6 & Onf7x6);
assign Onf7x6 = (~(Dtm7z6[0] & HRDATAD[19]));
assign Hnf7x6 = (~(Dtm7z6[1] & HRDATAS[19]));
assign Wkf7x6 = (~(Fcwnv6 & Ieyhw6));
assign Ieyhw6 = (JTAGNSW ? Aixmz6[19] : Ulxmz6[19]);
assign Mmx7v6 = (~(Vnf7x6 & Cof7x6));
assign Cof7x6 = (~(Idf7x6 & Itb7z6[20]));
assign Vnf7x6 = (Jof7x6 & Qof7x6);
assign Qof7x6 = (~(Xof7x6 & Kef7x6));
assign Xof7x6 = (~(Epf7x6 & Lpf7x6));
assign Lpf7x6 = (Spf7x6 & Zpf7x6);
assign Zpf7x6 = (Wawnv6 | Gqf7x6);
assign Spf7x6 = (~(Dtm7z6[3] & Nqf7x6));
assign Epf7x6 = (Uqf7x6 & Brf7x6);
assign Brf7x6 = (~(Dtm7z6[0] & HRDATAD[20]));
assign Uqf7x6 = (~(Dtm7z6[1] & HRDATAS[20]));
assign Jof7x6 = (~(Fcwnv6 & Ciyhw6));
assign Ciyhw6 = (JTAGNSW ? Aixmz6[20] : Ulxmz6[20]);
assign Fmx7v6 = (~(Irf7x6 & Prf7x6));
assign Prf7x6 = (~(Idf7x6 & Itb7z6[21]));
assign Irf7x6 = (Wrf7x6 & Dsf7x6);
assign Dsf7x6 = (~(Ksf7x6 & Kef7x6));
assign Ksf7x6 = (~(Rsf7x6 & Ysf7x6));
assign Ysf7x6 = (Ftf7x6 & Mtf7x6);
assign Mtf7x6 = (Wawnv6 | Ttf7x6);
assign Ftf7x6 = (~(Dtm7z6[3] & Auf7x6));
assign Rsf7x6 = (Huf7x6 & Ouf7x6);
assign Ouf7x6 = (~(Dtm7z6[0] & HRDATAD[21]));
assign Huf7x6 = (~(Dtm7z6[1] & HRDATAS[21]));
assign Wrf7x6 = (~(Fcwnv6 & Udyhw6));
assign Udyhw6 = (JTAGNSW ? Aixmz6[21] : Ulxmz6[21]);
assign Ylx7v6 = (~(Vuf7x6 & Cvf7x6));
assign Cvf7x6 = (~(Idf7x6 & Itb7z6[22]));
assign Vuf7x6 = (Jvf7x6 & Qvf7x6);
assign Qvf7x6 = (~(Xvf7x6 & Kef7x6));
assign Xvf7x6 = (~(Ewf7x6 & Lwf7x6));
assign Lwf7x6 = (Swf7x6 & Zwf7x6);
assign Zwf7x6 = (Wawnv6 | Gxf7x6);
assign Swf7x6 = (~(Dtm7z6[3] & Nxf7x6));
assign Ewf7x6 = (Uxf7x6 & Byf7x6);
assign Byf7x6 = (~(Dtm7z6[0] & HRDATAD[22]));
assign Uxf7x6 = (~(Dtm7z6[1] & HRDATAS[22]));
assign Jvf7x6 = (~(Fcwnv6 & Ohyhw6));
assign Ohyhw6 = (JTAGNSW ? Aixmz6[22] : Ulxmz6[22]);
assign Rlx7v6 = (~(Iyf7x6 & Pyf7x6));
assign Pyf7x6 = (~(Idf7x6 & Itb7z6[23]));
assign Iyf7x6 = (Wyf7x6 & Dzf7x6);
assign Dzf7x6 = (~(Kzf7x6 & Kef7x6));
assign Kzf7x6 = (~(Rzf7x6 & Yzf7x6));
assign Yzf7x6 = (F0g7x6 & M0g7x6);
assign M0g7x6 = (Wawnv6 | T0g7x6);
assign F0g7x6 = (~(Dtm7z6[3] & A1g7x6));
assign Rzf7x6 = (H1g7x6 & O1g7x6);
assign O1g7x6 = (~(Dtm7z6[0] & HRDATAD[23]));
assign H1g7x6 = (~(Dtm7z6[1] & HRDATAS[23]));
assign Wyf7x6 = (~(Fcwnv6 & Kfyhw6));
assign Kfyhw6 = (JTAGNSW ? Aixmz6[23] : Ulxmz6[23]);
assign Klx7v6 = (~(V1g7x6 & C2g7x6));
assign C2g7x6 = (~(Fcwnv6 & Sjyhw6));
assign Sjyhw6 = (JTAGNSW ? Aixmz6[16] : Ulxmz6[16]);
assign V1g7x6 = (J2g7x6 & Q2g7x6);
assign Q2g7x6 = (~(X2g7x6 & Kef7x6));
assign X2g7x6 = (~(E3g7x6 & L3g7x6));
assign L3g7x6 = (S3g7x6 & Z3g7x6);
assign Z3g7x6 = (Wawnv6 | G4g7x6);
assign S3g7x6 = (~(Dtm7z6[3] & N4g7x6));
assign E3g7x6 = (U4g7x6 & B5g7x6);
assign B5g7x6 = (~(Dtm7z6[0] & HRDATAD[16]));
assign U4g7x6 = (~(Dtm7z6[1] & HRDATAS[16]));
assign J2g7x6 = (~(Idf7x6 & Itb7z6[16]));
assign Idf7x6 = (~(Kef7x6 | Fvd7x6));
assign Kef7x6 = (~(I5g7x6 & P5g7x6));
assign P5g7x6 = (~(Ahe7x6 & W5g7x6));
assign W5g7x6 = (~(Ohe7x6 & D6g7x6));
assign D6g7x6 = (~(K6g7x6 & Ugo7z6[1]));
assign K6g7x6 = (Jie7x6 & Qie7x6);
assign I5g7x6 = (Eje7x6 | Ugo7z6[1]);
assign Eje7x6 = (~(R6g7x6 & Y6g7x6));
assign Y6g7x6 = (Ugo7z6[0] & Jie7x6);
assign R6g7x6 = (Ahe7x6 & Hub7z6[0]);
assign Dlx7v6 = (~(F7g7x6 & M7g7x6));
assign M7g7x6 = (~(L8wnv6 & Itb7z6[25]));
assign F7g7x6 = (T7g7x6 & A8g7x6);
assign A8g7x6 = (~(G9wnv6 & H8g7x6));
assign H8g7x6 = (~(O8g7x6 & V8g7x6));
assign V8g7x6 = (C9g7x6 & J9g7x6);
assign J9g7x6 = (Wawnv6 | Q9g7x6);
assign C9g7x6 = (~(Dtm7z6[3] & X9g7x6));
assign O8g7x6 = (Eag7x6 & Lag7x6);
assign Lag7x6 = (~(Dtm7z6[0] & HRDATAD[25]));
assign Eag7x6 = (~(Dtm7z6[1] & HRDATAS[25]));
assign T7g7x6 = (~(Fcwnv6 & Bsyhw6));
assign Bsyhw6 = (Dz1nv6 ? Ulxmz6[25] : Aixmz6[25]);
assign Wkx7v6 = (~(Sag7x6 & Zag7x6));
assign Zag7x6 = (~(L8wnv6 & Itb7z6[24]));
assign Sag7x6 = (Gbg7x6 & Nbg7x6);
assign Nbg7x6 = (~(G9wnv6 & Ubg7x6));
assign Ubg7x6 = (~(Bcg7x6 & Icg7x6));
assign Icg7x6 = (Pcg7x6 & Wcg7x6);
assign Wcg7x6 = (Wawnv6 | Ddg7x6);
assign Pcg7x6 = (~(Dtm7z6[3] & Kdg7x6));
assign Bcg7x6 = (Rdg7x6 & Ydg7x6);
assign Ydg7x6 = (~(Dtm7z6[0] & HRDATAD[24]));
assign Rdg7x6 = (~(Dtm7z6[1] & HRDATAS[24]));
assign Gbg7x6 = (~(Fcwnv6 & Psyhw6));
assign Psyhw6 = (JTAGNSW ? Aixmz6[24] : Ulxmz6[24]);
assign Pkx7v6 = (Mdonv6 ? Veonv6 : U8oet6);
assign Mdonv6 = (Rsdiw6 | Qteet6);
assign Ikx7v6 = (Sblov6 ? Feg7x6 : Wktet6);
assign Sblov6 = (Meg7x6 & Zy1ft6);
assign Meg7x6 = (Y94iw6 & Teg7x6);
assign Teg7x6 = (~(Afg7x6 & Hfg7x6));
assign Hfg7x6 = (~(Ofg7x6 & Vfg7x6));
assign Vfg7x6 = (Cgg7x6 & Gr2et6);
assign Cgg7x6 = (Wcmov6 & B2jnv6);
assign Ofg7x6 = (Xc1ft6 & Tk1ft6);
assign Afg7x6 = (~(Jgg7x6 & Qgg7x6));
assign Qgg7x6 = (~(Cegiw6 | K6adt6));
assign Cegiw6 = (!Gjdiw6);
assign Jgg7x6 = (Zb1ft6 & Jj1ft6);
assign Feg7x6 = (~(Xc1ft6 & Tk1ft6));
assign Bkx7v6 = (~(Xgg7x6 & Ehg7x6));
assign Ehg7x6 = (~(Lhg7x6 & Shg7x6));
assign Lhg7x6 = (Zhg7x6 & P52nv6);
assign Xgg7x6 = (~(Vveet6 & Gig7x6));
assign Gig7x6 = (~(Zhg7x6 & Nig7x6));
assign Nig7x6 = (~(Cwadt6 & Uig7x6));
assign Uig7x6 = (!Shg7x6);
assign Ujx7v6 = (Eofov6 & Qnfov6);
assign Qnfov6 = (~(Bjg7x6 & Ijg7x6));
assign Ijg7x6 = (~(Fe2nv6 & Pjg7x6));
assign Pjg7x6 = (~(Wjg7x6 & Dkg7x6));
assign Dkg7x6 = (Kkg7x6 & Rkg7x6);
assign Wjg7x6 = (Ykg7x6 & Kd2nv6);
assign Bjg7x6 = (Bcmov6 & Flg7x6);
assign Bcmov6 = (~(Mlg7x6 & Ebdiw6));
assign Mlg7x6 = (Zhg7x6 & Tlg7x6);
assign Tlg7x6 = (~(Amg7x6 & F52iw6));
assign Njx7v6 = (~(Hmg7x6 & Omg7x6));
assign Omg7x6 = (Wi2ov6 | Pcg7z6[31]);
assign Hmg7x6 = (Vmg7x6 & Cng7x6);
assign Cng7x6 = (~(Rj2ov6 & Ykmdt6));
assign Vmg7x6 = (~(Yj2ov6 & Yxf7z6[1]));
assign Gjx7v6 = (~(Jng7x6 & Qng7x6));
assign Qng7x6 = (~(Y3bov6 & Yxf7z6[1]));
assign Jng7x6 = (Xng7x6 & Eog7x6);
assign Eog7x6 = (~(Rj2ov6 & Mcmdt6));
assign Xng7x6 = (~(Yj2ov6 & Yxf7z6[5]));
assign Zix7v6 = (~(Log7x6 & Sog7x6));
assign Sog7x6 = (~(Y3bov6 & Yxf7z6[5]));
assign Log7x6 = (Zog7x6 & Gpg7x6);
assign Gpg7x6 = (~(Rj2ov6 & A4mdt6));
assign Zog7x6 = (~(Yj2ov6 & Yxf7z6[9]));
assign Six7v6 = (~(Npg7x6 & Upg7x6));
assign Upg7x6 = (~(Y3bov6 & Yxf7z6[9]));
assign Npg7x6 = (Bqg7x6 & Iqg7x6);
assign Iqg7x6 = (~(Rj2ov6 & Ovldt6));
assign Bqg7x6 = (~(Yj2ov6 & Yxf7z6[13]));
assign Lix7v6 = (~(Pqg7x6 & Wqg7x6));
assign Wqg7x6 = (~(Y3bov6 & Yxf7z6[13]));
assign Pqg7x6 = (Drg7x6 & Krg7x6);
assign Krg7x6 = (~(Rj2ov6 & Cnldt6));
assign Drg7x6 = (~(Yj2ov6 & Yxf7z6[17]));
assign Eix7v6 = (~(Rrg7x6 & Yrg7x6));
assign Yrg7x6 = (~(Y3bov6 & Yxf7z6[17]));
assign Rrg7x6 = (Fsg7x6 & Msg7x6);
assign Msg7x6 = (~(Rj2ov6 & Qeldt6));
assign Fsg7x6 = (~(Yj2ov6 & Yxf7z6[21]));
assign Xhx7v6 = (~(Tsg7x6 & Atg7x6));
assign Atg7x6 = (~(Y3bov6 & Yxf7z6[21]));
assign Tsg7x6 = (Htg7x6 & Otg7x6);
assign Otg7x6 = (~(Rj2ov6 & E6ldt6));
assign Htg7x6 = (~(Yj2ov6 & Yxf7z6[25]));
assign Qhx7v6 = (~(Vtg7x6 & Cug7x6));
assign Cug7x6 = (~(Y3bov6 & Yxf7z6[25]));
assign Vtg7x6 = (Jug7x6 & Qug7x6);
assign Qug7x6 = (~(Rj2ov6 & Sxkdt6));
assign Jug7x6 = (~(Yj2ov6 & Yxf7z6[29]));
assign Jhx7v6 = (~(Xug7x6 & Evg7x6));
assign Evg7x6 = (~(Yj2ov6 & Yxf7z6[33]));
assign Xug7x6 = (~(Y3bov6 & Yxf7z6[29]));
assign Chx7v6 = (Z6jhw6 ? D5f7z6[1] : Kknnv6);
assign Kknnv6 = (~(Lvg7x6 & Svg7x6));
assign Svg7x6 = (Zvg7x6 & Gwg7x6);
assign Gwg7x6 = (~(Ua0jw6 & Nwg7x6));
assign Nwg7x6 = (~(Xf0jw6 & Uwg7x6));
assign Uwg7x6 = (~(Bxg7x6 & Rc0jw6));
assign Bxg7x6 = (Wb0jw6 & Ixg7x6);
assign Ua0jw6 = (~(I40jw6 | Pxg7x6));
assign Zvg7x6 = (Wxg7x6 & Dyg7x6);
assign Dyg7x6 = (~(P40jw6 & Kyg7x6));
assign Kyg7x6 = (~(S90jw6 & Ryg7x6));
assign Ryg7x6 = (~(Yyg7x6 & M60jw6));
assign Yyg7x6 = (R50jw6 & Fzg7x6);
assign P40jw6 = (Mzg7x6 & Wwi6x6);
assign Mzg7x6 = (Tzg7x6 & Dxi6x6);
assign Dxi6x6 = (A0h7x6 | S90jw6);
assign S90jw6 = (~(H0h7x6 & Uu1jw6));
assign Uu1jw6 = (~(O0h7x6 | Fzg7x6));
assign Fzg7x6 = (~(V0h7x6 & C1h7x6));
assign C1h7x6 = (~(O70jw6 & J1h7x6));
assign V0h7x6 = (V70jw6 ? J1h7x6 : O70jw6);
assign V70jw6 = (Q1h7x6 & X1h7x6);
assign X1h7x6 = (~(E3c7z6[4] & E2h7x6));
assign Q1h7x6 = (~(Ijnnv6 & Onf7z6[4]));
assign O70jw6 = (~(L2h7x6 & S2h7x6));
assign S2h7x6 = (~(Fhc7z6[5] & E2h7x6));
assign L2h7x6 = (~(Ijnnv6 & Onf7z6[5]));
assign O0h7x6 = (~(M60jw6 & R50jw6));
assign R50jw6 = (Z2h7x6 ^ J1h7x6);
assign Z2h7x6 = (~(G3h7x6 & N3h7x6));
assign N3h7x6 = (~(Fhc7z6[7] & E2h7x6));
assign G3h7x6 = (~(Ijnnv6 & Onf7z6[7]));
assign M60jw6 = (U3h7x6 ^ J1h7x6);
assign U3h7x6 = (~(B4h7x6 & I4h7x6));
assign I4h7x6 = (~(Fhc7z6[6] & E2h7x6));
assign B4h7x6 = (~(Ijnnv6 & Onf7z6[6]));
assign H0h7x6 = (P4h7x6 & X80jw6);
assign X80jw6 = (W4h7x6 ^ J1h7x6);
assign W4h7x6 = (~(D5h7x6 & K5h7x6));
assign K5h7x6 = (~(E3c7z6[3] & E2h7x6));
assign D5h7x6 = (~(Ijnnv6 & Onf7z6[3]));
assign P4h7x6 = (J1h7x6 ^ J80jw6);
assign J80jw6 = (~(R5h7x6 & Y5h7x6));
assign Y5h7x6 = (~(E3c7z6[2] & E2h7x6));
assign R5h7x6 = (~(Ijnnv6 & Onf7z6[2]));
assign A0h7x6 = (F6h7x6 | Z90jw6);
assign Z90jw6 = (M6h7x6 ^ Tzziw6);
assign M6h7x6 = (~(T6h7x6 & A7h7x6));
assign A7h7x6 = (~(E3c7z6[1] & E2h7x6));
assign T6h7x6 = (~(Ijnnv6 & Onf7z6[1]));
assign F6h7x6 = (~(Tzziw6 ^ H7h7x6));
assign H7h7x6 = (O7h7x6 & V7h7x6);
assign V7h7x6 = (~(E3c7z6[0] & E2h7x6));
assign O7h7x6 = (~(Ijnnv6 & Onf7z6[0]));
assign Tzg7x6 = (!Kxi6x6);
assign Wxg7x6 = (~(Bxziw6 & C8h7x6));
assign C8h7x6 = (L20jw6 | J8h7x6);
assign J8h7x6 = (Q8h7x6 & Yyziw6);
assign Q8h7x6 = (Dyziw6 & X8h7x6);
assign Bxziw6 = (~(Kxi6x6 | Wwi6x6));
assign Wwi6x6 = (E9h7x6 & L20jw6);
assign L20jw6 = (L9h7x6 & Pv1jw6);
assign Pv1jw6 = (~(S9h7x6 | X8h7x6));
assign X8h7x6 = (~(Z9h7x6 & Gah7x6));
assign Gah7x6 = (~(H00jw6 & J1h7x6));
assign Z9h7x6 = (O00jw6 ? J1h7x6 : H00jw6);
assign O00jw6 = (Nah7x6 & Uah7x6);
assign Uah7x6 = (~(Fhc7z6[12] & E2h7x6));
assign Nah7x6 = (~(Ijnnv6 & Onf7z6[12]));
assign H00jw6 = (~(Bbh7x6 & Ibh7x6));
assign Ibh7x6 = (~(Fhc7z6[13] & E2h7x6));
assign Bbh7x6 = (~(Ijnnv6 & Onf7z6[13]));
assign S9h7x6 = (~(Yyziw6 & Dyziw6));
assign Dyziw6 = (Pbh7x6 ^ J1h7x6);
assign Pbh7x6 = (~(Wbh7x6 & Dch7x6));
assign Dch7x6 = (~(Fhc7z6[15] & E2h7x6));
assign Wbh7x6 = (~(Ijnnv6 & Onf7z6[15]));
assign Yyziw6 = (Kch7x6 ^ J1h7x6);
assign Kch7x6 = (~(Rch7x6 & Ych7x6));
assign Ych7x6 = (~(Fhc7z6[14] & E2h7x6));
assign Rch7x6 = (~(Ijnnv6 & Onf7z6[14]));
assign L9h7x6 = (Fdh7x6 & Q10jw6);
assign Q10jw6 = (Mdh7x6 ^ J1h7x6);
assign Mdh7x6 = (~(Tdh7x6 & Aeh7x6));
assign Aeh7x6 = (~(Fhc7z6[11] & E2h7x6));
assign Tdh7x6 = (~(Ijnnv6 & Onf7z6[11]));
assign Fdh7x6 = (J1h7x6 ^ C10jw6);
assign C10jw6 = (~(Heh7x6 & Oeh7x6));
assign Oeh7x6 = (~(Fhc7z6[10] & E2h7x6));
assign Heh7x6 = (~(Ijnnv6 & Onf7z6[10]));
assign E9h7x6 = (Veh7x6 & S20jw6);
assign S20jw6 = (Cfh7x6 ^ J1h7x6);
assign Cfh7x6 = (~(Jfh7x6 & Qfh7x6));
assign Qfh7x6 = (~(Fhc7z6[9] & E2h7x6));
assign Jfh7x6 = (~(Ijnnv6 & Onf7z6[9]));
assign Veh7x6 = (~(J1h7x6 ^ Xfh7x6));
assign Xfh7x6 = (Egh7x6 & Lgh7x6);
assign Lgh7x6 = (~(Fhc7z6[8] & E2h7x6));
assign Egh7x6 = (~(Ijnnv6 & Onf7z6[8]));
assign Kxi6x6 = (~(Sgh7x6 & Pxg7x6));
assign Pxg7x6 = (~(Zgh7x6 | Xf0jw6));
assign Xf0jw6 = (~(Ghh7x6 & Wv1jw6));
assign Wv1jw6 = (~(Nhh7x6 | Ixg7x6));
assign Ixg7x6 = (~(Uhh7x6 & Bih7x6));
assign Bih7x6 = (~(Td0jw6 & J1h7x6));
assign Uhh7x6 = (Ae0jw6 ? J1h7x6 : Td0jw6);
assign Ae0jw6 = (Iih7x6 & Pih7x6);
assign Pih7x6 = (~(Fhc7z6[20] & E2h7x6));
assign Iih7x6 = (~(Ijnnv6 & Onf7z6[20]));
assign Td0jw6 = (~(Wih7x6 & Djh7x6));
assign Djh7x6 = (~(Fhc7z6[21] & E2h7x6));
assign Wih7x6 = (~(Ijnnv6 & Onf7z6[21]));
assign Nhh7x6 = (~(Rc0jw6 & Wb0jw6));
assign Wb0jw6 = (Kjh7x6 ^ J1h7x6);
assign Kjh7x6 = (~(Rjh7x6 & Yjh7x6));
assign Yjh7x6 = (~(Fhc7z6[23] & E2h7x6));
assign Rjh7x6 = (~(Ijnnv6 & Onf7z6[23]));
assign Rc0jw6 = (Fkh7x6 ^ J1h7x6);
assign Fkh7x6 = (~(Mkh7x6 & Tkh7x6));
assign Tkh7x6 = (~(Fhc7z6[22] & E2h7x6));
assign Mkh7x6 = (~(Ijnnv6 & Onf7z6[22]));
assign Ghh7x6 = (Alh7x6 & Cf0jw6);
assign Cf0jw6 = (Hlh7x6 ^ J1h7x6);
assign Hlh7x6 = (~(Olh7x6 & Vlh7x6));
assign Vlh7x6 = (~(Fhc7z6[19] & E2h7x6));
assign Olh7x6 = (~(Ijnnv6 & Onf7z6[19]));
assign Alh7x6 = (J1h7x6 ^ Oe0jw6);
assign Oe0jw6 = (~(Cmh7x6 & Jmh7x6));
assign Jmh7x6 = (~(Fhc7z6[18] & E2h7x6));
assign Cmh7x6 = (~(Ijnnv6 & Onf7z6[18]));
assign Zgh7x6 = (Qmh7x6 | Eg0jw6);
assign Eg0jw6 = (Xmh7x6 ^ Tzziw6);
assign Xmh7x6 = (~(Enh7x6 & Lnh7x6));
assign Lnh7x6 = (~(Fhc7z6[17] & E2h7x6));
assign Enh7x6 = (~(Ijnnv6 & Onf7z6[17]));
assign Qmh7x6 = (~(Tzziw6 ^ Snh7x6));
assign Snh7x6 = (Znh7x6 & Goh7x6);
assign Goh7x6 = (~(Fhc7z6[16] & E2h7x6));
assign Znh7x6 = (~(Ijnnv6 & Onf7z6[16]));
assign Sgh7x6 = (!I40jw6);
assign Lvg7x6 = (Noh7x6 & Uoh7x6);
assign Uoh7x6 = (~(Gu1jw6 & Bph7x6));
assign Noh7x6 = (~(U30jw6 & I40jw6));
assign I40jw6 = (~(Iph7x6 & U30jw6));
assign Iph7x6 = (Pph7x6 & B40jw6);
assign B40jw6 = (Wph7x6 ^ J1h7x6);
assign Wph7x6 = (~(Dqh7x6 & Kqh7x6));
assign Kqh7x6 = (~(Fhc7z6[25] & E2h7x6));
assign Dqh7x6 = (~(Ijnnv6 & Onf7z6[25]));
assign Pph7x6 = (~(J1h7x6 ^ Rqh7x6));
assign Rqh7x6 = (Yqh7x6 & Frh7x6);
assign Frh7x6 = (~(Fhc7z6[24] & E2h7x6));
assign Yqh7x6 = (~(Ijnnv6 & Onf7z6[24]));
assign U30jw6 = (Mrh7x6 & Trh7x6);
assign Trh7x6 = (Ash7x6 & Fk0jw6);
assign Fk0jw6 = (!Dj0jw6);
assign Dj0jw6 = (Hsh7x6 ^ Tzziw6);
assign Hsh7x6 = (~(Osh7x6 & Vsh7x6));
assign Vsh7x6 = (~(Fhc7z6[26] & E2h7x6));
assign Osh7x6 = (~(Ijnnv6 & Onf7z6[26]));
assign Ash7x6 = (J1h7x6 ^ Kj0jw6);
assign Kj0jw6 = (~(Cth7x6 & Jth7x6));
assign Jth7x6 = (~(Fhc7z6[27] & E2h7x6));
assign Cth7x6 = (~(Ijnnv6 & Onf7z6[27]));
assign Mrh7x6 = (Gu1jw6 & Nu1jw6);
assign Nu1jw6 = (!Bph7x6);
assign Bph7x6 = (~(Qth7x6 & Xth7x6));
assign Xth7x6 = (~(Ii0jw6 & J1h7x6));
assign Qth7x6 = (Pi0jw6 ? J1h7x6 : Ii0jw6);
assign Pi0jw6 = (Euh7x6 & Luh7x6);
assign Luh7x6 = (~(Fhc7z6[28] & E2h7x6));
assign Euh7x6 = (~(Ijnnv6 & Onf7z6[28]));
assign Ii0jw6 = (~(Suh7x6 & Zuh7x6));
assign Zuh7x6 = (~(Fhc7z6[29] & E2h7x6));
assign Suh7x6 = (~(Ijnnv6 & Onf7z6[29]));
assign Gu1jw6 = (Gh0jw6 & Sg0jw6);
assign Sg0jw6 = (~(J1h7x6 & Gvh7x6));
assign Gvh7x6 = (~(Nvh7x6 & Uvh7x6));
assign Uvh7x6 = (~(Fhc7z6[31] & E2h7x6));
assign Nvh7x6 = (~(Ijnnv6 & Onf7z6[31]));
assign Gh0jw6 = (~(Bwh7x6 ^ Tzziw6));
assign Tzziw6 = (!J1h7x6);
assign J1h7x6 = (~(Rabov6 & N427x6));
assign N427x6 = (E327x6 & Fhc7z6[31]);
assign E327x6 = (Uh2ov6 & Mrbdt6);
assign Bwh7x6 = (~(Iwh7x6 & Pwh7x6));
assign Pwh7x6 = (~(Fhc7z6[30] & E2h7x6));
assign E2h7x6 = (Svziw6 | Rabov6);
assign Iwh7x6 = (~(Ijnnv6 & Onf7z6[30]));
assign Vgx7v6 = (K7tnv6 ? Yhzmz6[0] : ETMINTNUM[0]);
assign Ogx7v6 = (K7tnv6 ? Yhzmz6[1] : ETMINTNUM[1]);
assign Hgx7v6 = (K7tnv6 ? Yhzmz6[2] : ETMINTNUM[2]);
assign Agx7v6 = (K7tnv6 ? Yhzmz6[3] : ETMINTNUM[3]);
assign Tfx7v6 = (K7tnv6 ? Yhzmz6[4] : ETMINTNUM[4]);
assign Mfx7v6 = (K7tnv6 ? Zxymz6[5] : ETMINTNUM[5]);
assign Ffx7v6 = (K7tnv6 ? Zxymz6[6] : ETMINTNUM[6]);
assign Yex7v6 = (K7tnv6 ? Zxymz6[7] : ETMINTNUM[7]);
assign Rex7v6 = (K7tnv6 ? Zxymz6[8] : ETMINTNUM[8]);
assign K7tnv6 = (~(Wwh7x6 & Glh7v6));
assign Wwh7x6 = (Zkh7v6 & W3wnv6);
assign Kex7v6 = (~(Dxh7x6 & G1iov6));
assign G1iov6 = (~(Kxh7x6 & Rxh7x6));
assign Kxh7x6 = (Vzgov6 & Om2nv6);
assign Om2nv6 = (!Z3j7z6[7]);
assign Dxh7x6 = (Z3j7z6[7] ? Fyh7x6 : Yxh7x6);
assign Fyh7x6 = (~(Myh7x6 & Tyh7x6));
assign Tyh7x6 = (~(Egfiw6 & Wohov6));
assign Myh7x6 = (Azh7x6 & U4fov6);
assign Azh7x6 = (~(Kphov6 & Hzh7x6));
assign Yxh7x6 = (~(Wohov6 & R62nv6));
assign Dex7v6 = (~(Ozh7x6 & Ayhov6));
assign Ayhov6 = (~(Vzh7x6 & Vzgov6));
assign Vzh7x6 = (C0i7x6 & Vm2nv6);
assign Ozh7x6 = (Z3j7z6[8] ? Q0i7x6 : J0i7x6);
assign Q0i7x6 = (~(X0i7x6 & E1i7x6));
assign E1i7x6 = (~(Kphov6 & L1i7x6));
assign X0i7x6 = (S1i7x6 & U4fov6);
assign S1i7x6 = (~(Qlhov6 & Nhfiw6));
assign J0i7x6 = (~(Qlhov6 & U47iw6));
assign Wdx7v6 = (~(Z1i7x6 & G2i7x6));
assign Z1i7x6 = (Z3j7z6[10] ? U2i7x6 : N2i7x6);
assign U2i7x6 = (~(B3i7x6 & I3i7x6));
assign I3i7x6 = (~(Kphov6 & P3i7x6));
assign B3i7x6 = (W3i7x6 & U4fov6);
assign W3i7x6 = (~(Qlhov6 & Fkfiw6));
assign N2i7x6 = (~(Qlhov6 & H17iw6));
assign Pdx7v6 = (G5eov6 ? Oqbet6 : D4i7x6);
assign D4i7x6 = (K4i7x6 & G2i7x6);
assign G2i7x6 = (~(R4i7x6 & Vzgov6));
assign R4i7x6 = (Y4i7x6 & Qn2nv6);
assign Qn2nv6 = (!Z3j7z6[10]);
assign K4i7x6 = (~(Q0hov6 & H44iw6));
assign Idx7v6 = (~(F5i7x6 & M5i7x6));
assign F5i7x6 = (Z3j7z6[11] ? A6i7x6 : T5i7x6);
assign A6i7x6 = (~(H6i7x6 & O6i7x6));
assign O6i7x6 = (~(Kphov6 & V6i7x6));
assign H6i7x6 = (C7i7x6 & U4fov6);
assign C7i7x6 = (~(Qlhov6 & Olfiw6));
assign T5i7x6 = (~(Qlhov6 & Dz6iw6));
assign Bdx7v6 = (!Z4eov6);
assign Z4eov6 = (Zfcet6 ? Q7i7x6 : J7i7x6);
assign Q7i7x6 = (~(X7i7x6 & M5i7x6));
assign M5i7x6 = (~(E8i7x6 & K4hov6));
assign E8i7x6 = (~(Kxgov6 | Z3j7z6[11]));
assign Kxgov6 = (!Vzgov6);
assign X7i7x6 = (~(Q0hov6 & Iklov6));
assign J7i7x6 = (L8i7x6 & S8i7x6);
assign S8i7x6 = (~(M5bdt6 & Z8i7x6));
assign Z8i7x6 = (~(Jqj7z6[8] & Z3j7z6[11]));
assign L8i7x6 = (~(Q0hov6 & E64iw6));
assign Ucx7v6 = (~(G9i7x6 & N9i7x6));
assign N9i7x6 = (U9i7x6 | Fsliw6);
assign G9i7x6 = (Bai7x6 & Iai7x6);
assign Bai7x6 = (Z3fov6 | Zo2nv6);
assign Ncx7v6 = (!Pai7x6);
assign Pai7x6 = (M6j7z6[8] ? Dbi7x6 : Wai7x6);
assign Dbi7x6 = (~(Kbi7x6 & Iai7x6));
assign Iai7x6 = (~(Rbi7x6 & H0miw6));
assign Rbi7x6 = (Ybi7x6 & Zo2nv6);
assign Zo2nv6 = (!G5j7z6[8]);
assign Kbi7x6 = (~(Fci7x6 & U47iw6));
assign Wai7x6 = (Mci7x6 & Tci7x6);
assign Tci7x6 = (~(Adi7x6 & U47iw6));
assign Mci7x6 = (~(Qkj7z6[8] | Hdi7x6));
assign Hdi7x6 = (Odi7x6 & Tib7z6[8]);
assign Odi7x6 = (~(Jqj7z6[17] & G5j7z6[8]));
assign Gcx7v6 = (~(Vdi7x6 & Cei7x6));
assign Cei7x6 = (~(G5j7z6[9] & Jei7x6));
assign Jei7x6 = (~(Vtliw6 & Qei7x6));
assign Zbx7v6 = (!Xei7x6);
assign Xei7x6 = (M6j7z6[9] ? Lfi7x6 : Efi7x6);
assign Lfi7x6 = (~(Vdi7x6 & Sfi7x6));
assign Sfi7x6 = (~(Fci7x6 & J27iw6));
assign Vdi7x6 = (~(Zfi7x6 & H0miw6));
assign Zfi7x6 = (Ggi7x6 & Gp2nv6);
assign Gp2nv6 = (!G5j7z6[9]);
assign Efi7x6 = (Ngi7x6 & Ugi7x6);
assign Ugi7x6 = (~(Adi7x6 & J27iw6));
assign Ngi7x6 = (~(Qkj7z6[9] | Bhi7x6));
assign Bhi7x6 = (Ihi7x6 & Tib7z6[9]);
assign Ihi7x6 = (~(Jqj7z6[18] & G5j7z6[9]));
assign Sbx7v6 = (~(Phi7x6 & Whi7x6));
assign Whi7x6 = (~(Dii7x6 & U4fov6));
assign Phi7x6 = (Kii7x6 & Rii7x6);
assign Kii7x6 = (Z3fov6 | Lv2nv6);
assign Lbx7v6 = (!Yii7x6);
assign Yii7x6 = (M6j7z6[10] ? Mji7x6 : Fji7x6);
assign Mji7x6 = (~(Tji7x6 & Rii7x6));
assign Rii7x6 = (~(Aki7x6 & H0miw6));
assign Aki7x6 = (Hki7x6 & Lv2nv6);
assign Lv2nv6 = (!G5j7z6[10]);
assign Tji7x6 = (~(Fci7x6 & H17iw6));
assign Fji7x6 = (Oki7x6 & Vki7x6);
assign Vki7x6 = (~(Adi7x6 & H17iw6));
assign Oki7x6 = (~(Qkj7z6[10] | Cli7x6));
assign Cli7x6 = (Jli7x6 & Tib7z6[10]);
assign Jli7x6 = (~(Jqj7z6[19] & G5j7z6[10]));
assign Ebx7v6 = (~(Qli7x6 & Xli7x6));
assign Xli7x6 = (~(Emi7x6 & U4fov6));
assign Qli7x6 = (Lmi7x6 & Smi7x6);
assign Lmi7x6 = (Z3fov6 | Vt2nv6);
assign Xax7v6 = (!Zmi7x6);
assign Zmi7x6 = (M6j7z6[11] ? Nni7x6 : Gni7x6);
assign Nni7x6 = (~(Uni7x6 & Smi7x6));
assign Smi7x6 = (~(Boi7x6 & H0miw6));
assign Boi7x6 = (Rxh7x6 & Vt2nv6);
assign Vt2nv6 = (!G5j7z6[11]);
assign Uni7x6 = (~(Fci7x6 & Dz6iw6));
assign Gni7x6 = (Ioi7x6 & Poi7x6);
assign Poi7x6 = (~(Adi7x6 & Dz6iw6));
assign Ioi7x6 = (~(Qkj7z6[11] | Woi7x6));
assign Woi7x6 = (Dpi7x6 & Tib7z6[11]);
assign Dpi7x6 = (~(Jqj7z6[20] & G5j7z6[11]));
assign Qax7v6 = (~(Kpi7x6 & Rpi7x6));
assign Rpi7x6 = (~(G5j7z6[12] & Ypi7x6));
assign Ypi7x6 = (Fqi7x6 | Mqi7x6);
assign Jax7v6 = (!Tqi7x6);
assign Tqi7x6 = (M6j7z6[12] ? Hri7x6 : Ari7x6);
assign Hri7x6 = (~(Ori7x6 & Kpi7x6));
assign Kpi7x6 = (~(Vri7x6 & H0miw6));
assign Vri7x6 = (C0i7x6 & Csi7x6);
assign Ori7x6 = (~(Fci7x6 & Emhov6));
assign Ari7x6 = (Jsi7x6 & Qsi7x6);
assign Qsi7x6 = (~(Adi7x6 & Emhov6));
assign Jsi7x6 = (~(Qkj7z6[12] | Xsi7x6));
assign Xsi7x6 = (Eti7x6 & Tib7z6[12]);
assign Eti7x6 = (~(Jqj7z6[21] & G5j7z6[12]));
assign Cax7v6 = (~(Lti7x6 & Sti7x6));
assign Sti7x6 = (~(G5j7z6[13] & Zti7x6));
assign Zti7x6 = (Fqi7x6 | Gui7x6);
assign V9x7v6 = (!Nui7x6);
assign Nui7x6 = (M6j7z6[13] ? Bvi7x6 : Uui7x6);
assign Bvi7x6 = (~(Lti7x6 & Ivi7x6));
assign Ivi7x6 = (~(Fci7x6 & Guhov6));
assign Lti7x6 = (~(Pvi7x6 & H0miw6));
assign Pvi7x6 = (Wvi7x6 & Dwi7x6);
assign Uui7x6 = (Kwi7x6 & Rwi7x6);
assign Rwi7x6 = (~(Adi7x6 & Guhov6));
assign Kwi7x6 = (~(Qkj7z6[13] | Ywi7x6));
assign Ywi7x6 = (Fxi7x6 & Tib7z6[13]);
assign Fxi7x6 = (~(Jqj7z6[22] & G5j7z6[13]));
assign O9x7v6 = (~(Mxi7x6 & Txi7x6));
assign Txi7x6 = (~(G5j7z6[14] & Ayi7x6));
assign Ayi7x6 = (Fqi7x6 | Rwhov6);
assign Fqi7x6 = (!Vtliw6);
assign H9x7v6 = (!Hyi7x6);
assign Hyi7x6 = (M6j7z6[14] ? Vyi7x6 : Oyi7x6);
assign Vyi7x6 = (~(Mxi7x6 & Czi7x6));
assign Czi7x6 = (~(Fci7x6 & Bk6iw6));
assign Mxi7x6 = (~(Jzi7x6 & H0miw6));
assign Jzi7x6 = (Y4i7x6 & Qzi7x6);
assign Oyi7x6 = (Xzi7x6 & E0j7x6);
assign E0j7x6 = (~(Adi7x6 & Bk6iw6));
assign Xzi7x6 = (~(Qkj7z6[14] | L0j7x6));
assign L0j7x6 = (S0j7x6 & Tib7z6[14]);
assign S0j7x6 = (~(Jqj7z6[23] & G5j7z6[14]));
assign A9x7v6 = (~(Z0j7x6 & G1j7x6));
assign G1j7x6 = (~(G5j7z6[15] & N1j7x6));
assign N1j7x6 = (~(Vtliw6 & N2hov6));
assign N2hov6 = (V6i7x6 | Fsliw6);
assign Vtliw6 = (U1j7x6 & Z3fov6);
assign U1j7x6 = (~(B2j7x6 & U4fov6));
assign T8x7v6 = (!I2j7x6);
assign I2j7x6 = (M6j7z6[15] ? W2j7x6 : P2j7x6);
assign W2j7x6 = (~(Z0j7x6 & D3j7x6));
assign D3j7x6 = (~(Fci7x6 & Z0iov6));
assign Fci7x6 = (K3j7x6 & Bqi7z6[1]);
assign K3j7x6 = (!Arniw6);
assign Z0j7x6 = (~(R3j7x6 & H0miw6));
assign H0miw6 = (Y3j7x6 & F4j7x6);
assign Y3j7x6 = (Sa2nv6 & P2j7z6[4]);
assign R3j7x6 = (K4hov6 & M4j7x6);
assign P2j7x6 = (T4j7x6 & A5j7x6);
assign A5j7x6 = (~(Adi7x6 & Z0iov6));
assign Adi7x6 = (H5j7x6 & Bqi7z6[1]);
assign H5j7x6 = (!Qsniw6);
assign T4j7x6 = (~(Qkj7z6[15] | O5j7x6));
assign O5j7x6 = (V5j7x6 & Tib7z6[15]);
assign V5j7x6 = (~(Jqj7z6[24] & G5j7z6[15]));
assign M8x7v6 = (~(C6j7x6 & J6j7x6));
assign J6j7x6 = (~(G5j7z6[24] & Q6j7x6));
assign Q6j7x6 = (~(Wimiw6 & X6j7x6));
assign F8x7v6 = (!E7j7x6);
assign E7j7x6 = (M6j7z6[24] ? S7j7x6 : L7j7x6);
assign S7j7x6 = (~(Z7j7x6 & C6j7x6));
assign C6j7x6 = (~(G8j7x6 & Dcmiw6));
assign G8j7x6 = (Ybi7x6 & N8j7x6);
assign Z7j7x6 = (~(U8j7x6 & Wf4iw6));
assign L7j7x6 = (B9j7x6 & I9j7x6);
assign I9j7x6 = (~(P9j7x6 & Wf4iw6));
assign B9j7x6 = (~(Qkj7z6[24] | W9j7x6));
assign W9j7x6 = (Daj7x6 & Tib7z6[24]);
assign Daj7x6 = (~(Jqj7z6[33] & G5j7z6[24]));
assign Y7x7v6 = (~(Kaj7x6 & Raj7x6));
assign Raj7x6 = (~(Yaj7x6 & G5j7z6[25]));
assign Yaj7x6 = (Fbj7x6 & U4fov6);
assign Fbj7x6 = (~(Cfmiw6 & Mbj7x6));
assign R7x7v6 = (!Tbj7x6);
assign Tbj7x6 = (M6j7z6[25] ? Hcj7x6 : Acj7x6);
assign Hcj7x6 = (~(Kaj7x6 & Ocj7x6));
assign Ocj7x6 = (~(U8j7x6 & Iklov6));
assign Kaj7x6 = (~(Vcj7x6 & Dcmiw6));
assign Vcj7x6 = (Ggi7x6 & Cdj7x6);
assign Acj7x6 = (Jdj7x6 & Qdj7x6);
assign Qdj7x6 = (~(P9j7x6 & Iklov6));
assign Jdj7x6 = (~(Qkj7z6[25] | Xdj7x6));
assign Xdj7x6 = (Eej7x6 & Tib7z6[25]);
assign Eej7x6 = (~(Jqj7z6[34] & G5j7z6[25]));
assign K7x7v6 = (~(Lej7x6 & Sej7x6));
assign Sej7x6 = (~(Zej7x6 & G5j7z6[26]));
assign Zej7x6 = (Gfj7x6 & U4fov6);
assign Gfj7x6 = (~(Cfmiw6 & Nfj7x6));
assign D7x7v6 = (!Ufj7x6);
assign Ufj7x6 = (M6j7z6[26] ? Igj7x6 : Bgj7x6);
assign Igj7x6 = (~(Lej7x6 & Pgj7x6));
assign Pgj7x6 = (~(U8j7x6 & E64iw6));
assign Lej7x6 = (~(Wgj7x6 & Dcmiw6));
assign Wgj7x6 = (Hki7x6 & Dhj7x6);
assign Bgj7x6 = (Khj7x6 & Rhj7x6);
assign Rhj7x6 = (~(P9j7x6 & E64iw6));
assign Khj7x6 = (~(Qkj7z6[26] | Yhj7x6));
assign Yhj7x6 = (Fij7x6 & Tib7z6[26]);
assign Fij7x6 = (~(Jqj7z6[35] & G5j7z6[26]));
assign W6x7v6 = (~(Mij7x6 & Tij7x6));
assign Tij7x6 = (~(Ajj7x6 & G5j7z6[27]));
assign Ajj7x6 = (Hjj7x6 & U4fov6);
assign Hjj7x6 = (~(Cfmiw6 & Hzh7x6));
assign P6x7v6 = (!Ojj7x6);
assign Ojj7x6 = (M6j7z6[27] ? Ckj7x6 : Vjj7x6);
assign Ckj7x6 = (~(Mij7x6 & Jkj7x6));
assign Jkj7x6 = (~(U8j7x6 & H44iw6));
assign Mij7x6 = (~(Qkj7x6 & Dcmiw6));
assign Qkj7x6 = (Rxh7x6 & Xkj7x6);
assign Vjj7x6 = (Elj7x6 & Llj7x6);
assign Llj7x6 = (~(P9j7x6 & H44iw6));
assign Elj7x6 = (~(Qkj7z6[27] | Slj7x6));
assign Slj7x6 = (Zlj7x6 & Tib7z6[27]);
assign Zlj7x6 = (~(Jqj7z6[36] & G5j7z6[27]));
assign I6x7v6 = (~(Gmj7x6 & Nmj7x6));
assign Nmj7x6 = (~(G5j7z6[28] & Umj7x6));
assign Umj7x6 = (S9miw6 | Mqi7x6);
assign S9miw6 = (!Wimiw6);
assign Wimiw6 = (Z3fov6 & Bnj7x6);
assign Bnj7x6 = (~(U4fov6 & Inj7x6));
assign B6x7v6 = (!Pnj7x6);
assign Pnj7x6 = (M6j7z6[28] ? Doj7x6 : Wnj7x6);
assign Doj7x6 = (~(Koj7x6 & Gmj7x6));
assign Gmj7x6 = (~(Roj7x6 & Dcmiw6));
assign Roj7x6 = (C0i7x6 & Yoj7x6);
assign Koj7x6 = (~(U8j7x6 & W14iw6));
assign Wnj7x6 = (Fpj7x6 & Mpj7x6);
assign Mpj7x6 = (~(P9j7x6 & W14iw6));
assign Fpj7x6 = (~(Qkj7z6[28] | Tpj7x6));
assign Tpj7x6 = (Aqj7x6 & Tib7z6[28]);
assign Aqj7x6 = (~(Jqj7z6[37] & G5j7z6[28]));
assign U5x7v6 = (~(Hqj7x6 & Oqj7x6));
assign Oqj7x6 = (~(Vqj7x6 & G5j7z6[29]));
assign Vqj7x6 = (Crj7x6 & U4fov6);
assign Crj7x6 = (~(Cfmiw6 & Jrj7x6));
assign N5x7v6 = (!Qrj7x6);
assign Qrj7x6 = (M6j7z6[29] ? Esj7x6 : Xrj7x6);
assign Esj7x6 = (~(Hqj7x6 & Lsj7x6));
assign Lsj7x6 = (~(U8j7x6 & Zz3iw6));
assign Hqj7x6 = (~(Ssj7x6 & Dcmiw6));
assign Ssj7x6 = (Wvi7x6 & Zsj7x6);
assign Xrj7x6 = (Gtj7x6 & Ntj7x6);
assign Ntj7x6 = (~(P9j7x6 & Zz3iw6));
assign Gtj7x6 = (~(Qkj7z6[29] | Utj7x6));
assign Utj7x6 = (Buj7x6 & Tib7z6[29]);
assign Buj7x6 = (~(Jqj7z6[38] & G5j7z6[29]));
assign G5x7v6 = (~(Iuj7x6 & Puj7x6));
assign Puj7x6 = (~(Wuj7x6 & G5j7z6[30]));
assign Wuj7x6 = (Dvj7x6 & U4fov6);
assign Dvj7x6 = (~(Cfmiw6 & P3i7x6));
assign Z4x7v6 = (!Kvj7x6);
assign Kvj7x6 = (M6j7z6[30] ? Yvj7x6 : Rvj7x6);
assign Yvj7x6 = (~(Iuj7x6 & Fwj7x6));
assign Fwj7x6 = (~(U8j7x6 & Ro3iw6));
assign Iuj7x6 = (~(Mwj7x6 & Dcmiw6));
assign Mwj7x6 = (Y4i7x6 & Twj7x6);
assign Rvj7x6 = (Axj7x6 & Hxj7x6);
assign Hxj7x6 = (~(P9j7x6 & Ro3iw6));
assign Axj7x6 = (~(Qkj7z6[30] | Oxj7x6));
assign Oxj7x6 = (Vxj7x6 & Tib7z6[30]);
assign Vxj7x6 = (~(Jqj7z6[39] & G5j7z6[30]));
assign S4x7v6 = (~(Cyj7x6 & Jyj7x6));
assign Jyj7x6 = (~(Qyj7x6 & G5j7z6[31]));
assign Qyj7x6 = (Xyj7x6 & U4fov6);
assign Xyj7x6 = (~(Cfmiw6 & V6i7x6));
assign Cfmiw6 = (~(Sh2nv6 | Inj7x6));
assign L4x7v6 = (!Ezj7x6);
assign Ezj7x6 = (M6j7z6[31] ? Szj7x6 : Lzj7x6);
assign Szj7x6 = (~(Cyj7x6 & Zzj7x6));
assign Zzj7x6 = (~(U8j7x6 & X0hov6));
assign U8j7x6 = (~(Arniw6 | Dv3iw6));
assign Arniw6 = (~(Pceiw6 & G0k7x6));
assign Pceiw6 = (Toi7z6[7] & Pb8iw6);
assign Cyj7x6 = (~(N0k7x6 & Dcmiw6));
assign Dcmiw6 = (~(U0k7x6 | P2j7z6[4]));
assign N0k7x6 = (K4hov6 & B1k7x6);
assign K4hov6 = (I1k7x6 & Rc3nv6);
assign I1k7x6 = (P2j7z6[0] & P2j7z6[1]);
assign Lzj7x6 = (P1k7x6 & W1k7x6);
assign W1k7x6 = (~(P9j7x6 & X0hov6));
assign P9j7x6 = (~(Qsniw6 | Dv3iw6));
assign Qsniw6 = (~(Ddeiw6 & G0k7x6));
assign Ddeiw6 = (Pb8iw6 & D2k7x6);
assign P1k7x6 = (~(Qkj7z6[31] | K2k7x6));
assign K2k7x6 = (R2k7x6 & Tib7z6[31]);
assign R2k7x6 = (~(Jqj7z6[40] & G5j7z6[31]));
assign E4x7v6 = (~(Y2k7x6 & F3k7x6));
assign F3k7x6 = (~(G5j7z6[40] & M3k7x6));
assign M3k7x6 = (~(Kqmiw6 & X6j7x6));
assign X6j7x6 = (~(U4fov6 & T3k7x6));
assign Kqmiw6 = (!A4k7x6);
assign X3x7v6 = (!H4k7x6);
assign H4k7x6 = (M6j7z6[40] ? V4k7x6 : O4k7x6);
assign V4k7x6 = (~(C5k7x6 & Y2k7x6));
assign Y2k7x6 = (~(J5k7x6 & A5iov6));
assign J5k7x6 = (Ybi7x6 & Q5k7x6);
assign C5k7x6 = (~(M4iov6 & U47iw6));
assign O4k7x6 = (X5k7x6 & E6k7x6);
assign E6k7x6 = (~(C6iov6 & U47iw6));
assign X5k7x6 = (~(Qkj7z6[40] | L6k7x6));
assign L6k7x6 = (S6k7x6 & Tib7z6[40]);
assign S6k7x6 = (~(Jqj7z6[49] & G5j7z6[40]));
assign Q3x7v6 = (~(Z6k7x6 & G7k7x6));
assign G7k7x6 = (~(G5j7z6[41] & N7k7x6));
assign N7k7x6 = (~(D3iov6 & Qei7x6));
assign Qei7x6 = (~(U4fov6 & U7k7x6));
assign J3x7v6 = (!B8k7x6);
assign B8k7x6 = (M6j7z6[41] ? P8k7x6 : I8k7x6);
assign P8k7x6 = (~(Z6k7x6 & W8k7x6));
assign W8k7x6 = (~(M4iov6 & J27iw6));
assign Z6k7x6 = (~(D9k7x6 & A5iov6));
assign D9k7x6 = (Ggi7x6 & K9k7x6);
assign I8k7x6 = (R9k7x6 & Y9k7x6);
assign Y9k7x6 = (~(C6iov6 & J27iw6));
assign R9k7x6 = (~(Qkj7z6[41] | Fak7x6));
assign Fak7x6 = (Mak7x6 & Tib7z6[41]);
assign Mak7x6 = (~(Jqj7z6[50] & G5j7z6[41]));
assign C3x7v6 = (~(Tak7x6 & Abk7x6));
assign Abk7x6 = (~(G5j7z6[42] & Hbk7x6));
assign Hbk7x6 = (~(D3iov6 & Obk7x6));
assign V2x7v6 = (!Vbk7x6);
assign Vbk7x6 = (M6j7z6[42] ? Jck7x6 : Cck7x6);
assign Jck7x6 = (~(Tak7x6 & Qck7x6));
assign Qck7x6 = (~(M4iov6 & H17iw6));
assign Tak7x6 = (~(Xck7x6 & A5iov6));
assign Xck7x6 = (Hki7x6 & Edk7x6);
assign Cck7x6 = (Ldk7x6 & Sdk7x6);
assign Sdk7x6 = (~(C6iov6 & H17iw6));
assign Ldk7x6 = (~(Qkj7z6[42] | Zdk7x6));
assign Zdk7x6 = (Gek7x6 & Tib7z6[42]);
assign Gek7x6 = (~(Jqj7z6[51] & G5j7z6[42]));
assign O2x7v6 = (~(Nek7x6 & Uek7x6));
assign Uek7x6 = (~(G5j7z6[43] & Bfk7x6));
assign Bfk7x6 = (~(D3iov6 & Ifk7x6));
assign Ifk7x6 = (~(Pfk7x6 & U4fov6));
assign H2x7v6 = (!Wfk7x6);
assign Wfk7x6 = (M6j7z6[43] ? Kgk7x6 : Dgk7x6);
assign Kgk7x6 = (~(Nek7x6 & Rgk7x6));
assign Rgk7x6 = (~(M4iov6 & Dz6iw6));
assign Nek7x6 = (~(Ygk7x6 & A5iov6));
assign Ygk7x6 = (Rxh7x6 & Fhk7x6);
assign Dgk7x6 = (Mhk7x6 & Thk7x6);
assign Thk7x6 = (~(C6iov6 & Dz6iw6));
assign Mhk7x6 = (~(Qkj7z6[43] | Aik7x6));
assign Aik7x6 = (Hik7x6 & Tib7z6[43]);
assign Hik7x6 = (~(Jqj7z6[52] & G5j7z6[43]));
assign A2x7v6 = (~(Oik7x6 & Vik7x6));
assign Vik7x6 = (~(G5j7z6[44] & Cjk7x6));
assign Cjk7x6 = (A4k7x6 | Mqi7x6);
assign A4k7x6 = (~(Z3fov6 & Jjk7x6));
assign Jjk7x6 = (Fsliw6 | Qjk7x6);
assign T1x7v6 = (!Xjk7x6);
assign Xjk7x6 = (M6j7z6[44] ? Lkk7x6 : Ekk7x6);
assign Lkk7x6 = (~(Skk7x6 & Oik7x6));
assign Oik7x6 = (~(Zkk7x6 & A5iov6));
assign Zkk7x6 = (C0i7x6 & Glk7x6);
assign Skk7x6 = (~(M4iov6 & Emhov6));
assign Ekk7x6 = (Nlk7x6 & Ulk7x6);
assign Ulk7x6 = (~(C6iov6 & Emhov6));
assign Nlk7x6 = (~(Qkj7z6[44] | Bmk7x6));
assign Bmk7x6 = (Imk7x6 & Tib7z6[44]);
assign Imk7x6 = (~(Jqj7z6[53] & G5j7z6[44]));
assign M1x7v6 = (~(Pmk7x6 & Wmk7x6));
assign Wmk7x6 = (~(G5j7z6[45] & Dnk7x6));
assign Dnk7x6 = (Knk7x6 | Gui7x6);
assign F1x7v6 = (!Rnk7x6);
assign Rnk7x6 = (M6j7z6[45] ? Fok7x6 : Ynk7x6);
assign Fok7x6 = (~(Pmk7x6 & Mok7x6));
assign Mok7x6 = (~(M4iov6 & Guhov6));
assign Pmk7x6 = (~(Tok7x6 & A5iov6));
assign Tok7x6 = (Wvi7x6 & Apk7x6);
assign Ynk7x6 = (Hpk7x6 & Opk7x6);
assign Opk7x6 = (~(C6iov6 & Guhov6));
assign Hpk7x6 = (~(Qkj7z6[45] | Vpk7x6));
assign Vpk7x6 = (Cqk7x6 & Tib7z6[45]);
assign Cqk7x6 = (~(Jqj7z6[54] & G5j7z6[45]));
assign Y0x7v6 = (~(Jqk7x6 & Qqk7x6));
assign Qqk7x6 = (~(G5j7z6[46] & Xqk7x6));
assign Xqk7x6 = (Knk7x6 | Rwhov6);
assign Rwhov6 = (U4fov6 & Erk7x6);
assign Knk7x6 = (!D3iov6);
assign D3iov6 = (~(Lrk7x6 & U4fov6));
assign Lrk7x6 = (~(Sugov6 & Qjk7x6));
assign R0x7v6 = (!Srk7x6);
assign Srk7x6 = (M6j7z6[46] ? Gsk7x6 : Zrk7x6);
assign Gsk7x6 = (~(Jqk7x6 & Nsk7x6));
assign Nsk7x6 = (~(M4iov6 & Bk6iw6));
assign M4iov6 = (~(Nmoiw6 | Nq6iw6));
assign Jqk7x6 = (~(Usk7x6 & A5iov6));
assign A5iov6 = (~(U0k7x6 | E7iov6));
assign U0k7x6 = (~(Btk7x6 & Sa2nv6));
assign Btk7x6 = (P2j7z6[5] & Wfjov6);
assign Usk7x6 = (Y4i7x6 & Itk7x6);
assign Zrk7x6 = (Ptk7x6 & Wtk7x6);
assign Wtk7x6 = (~(C6iov6 & Bk6iw6));
assign C6iov6 = (~(Dooiw6 | Nq6iw6));
assign Ptk7x6 = (~(Qkj7z6[46] | Duk7x6));
assign Duk7x6 = (Kuk7x6 & Tib7z6[46]);
assign Kuk7x6 = (~(Jqj7z6[55] & G5j7z6[46]));
assign K0x7v6 = (~(Ruk7x6 & Yuk7x6));
assign Yuk7x6 = (~(Fvk7x6 & U4fov6));
assign Ruk7x6 = (Mvk7x6 & Tvk7x6);
assign Mvk7x6 = (Z3fov6 | Up2nv6);
assign D0x7v6 = (!Awk7x6);
assign Awk7x6 = (M6j7z6[56] ? Owk7x6 : Hwk7x6);
assign Owk7x6 = (~(Vwk7x6 & Tvk7x6));
assign Tvk7x6 = (~(Cxk7x6 & Ybi7x6));
assign Ybi7x6 = (~(Jxk7x6 | P2j7z6[0]));
assign Cxk7x6 = (R4hov6 & Up2nv6);
assign Up2nv6 = (!G5j7z6[56]);
assign Vwk7x6 = (~(W3hov6 & Wf4iw6));
assign Hwk7x6 = (Qxk7x6 & Xxk7x6);
assign Xxk7x6 = (~(T5hov6 & Wf4iw6));
assign Qxk7x6 = (~(Qkj7z6[56] | Eyk7x6));
assign Eyk7x6 = (Lyk7x6 & Tib7z6[56]);
assign Lyk7x6 = (~(Jqj7z6[65] & G5j7z6[56]));
assign Wzw7v6 = (~(Syk7x6 & Zyk7x6));
assign Zyk7x6 = (~(Gzk7x6 & U4fov6));
assign Syk7x6 = (Nzk7x6 & Uzk7x6);
assign Nzk7x6 = (Z3fov6 | Bq2nv6);
assign Pzw7v6 = (!B0l7x6);
assign B0l7x6 = (M6j7z6[57] ? P0l7x6 : I0l7x6);
assign P0l7x6 = (~(W0l7x6 & Uzk7x6));
assign Uzk7x6 = (~(D1l7x6 & Ggi7x6));
assign Ggi7x6 = (~(Jxk7x6 | Bgiov6));
assign Jxk7x6 = (~(K1l7x6 & P2j7z6[3]));
assign K1l7x6 = (Rgjov6 & U1iov6);
assign D1l7x6 = (R4hov6 & Bq2nv6);
assign Bq2nv6 = (!G5j7z6[57]);
assign W0l7x6 = (~(W3hov6 & Iklov6));
assign I0l7x6 = (R1l7x6 & Y1l7x6);
assign Y1l7x6 = (~(T5hov6 & Iklov6));
assign R1l7x6 = (~(Qkj7z6[57] | F2l7x6));
assign F2l7x6 = (M2l7x6 & Tib7z6[57]);
assign M2l7x6 = (~(Jqj7z6[66] & G5j7z6[57]));
assign Izw7v6 = (~(T2l7x6 & A3l7x6));
assign A3l7x6 = (~(G5j7z6[58] & H3l7x6));
assign H3l7x6 = (~(G2hov6 & Obk7x6));
assign Obk7x6 = (~(U4fov6 & O3l7x6));
assign Bzw7v6 = (!V3l7x6);
assign V3l7x6 = (M6j7z6[58] ? J4l7x6 : C4l7x6);
assign J4l7x6 = (~(T2l7x6 & Q4l7x6));
assign Q4l7x6 = (~(W3hov6 & E64iw6));
assign T2l7x6 = (~(X4l7x6 & Hki7x6));
assign Hki7x6 = (~(E5l7x6 | P2j7z6[0]));
assign X4l7x6 = (R4hov6 & Iq2nv6);
assign C4l7x6 = (L5l7x6 & S5l7x6);
assign S5l7x6 = (~(T5hov6 & E64iw6));
assign L5l7x6 = (~(Qkj7z6[58] | Z5l7x6));
assign Z5l7x6 = (G6l7x6 & Tib7z6[58]);
assign G6l7x6 = (~(Jqj7z6[67] & G5j7z6[58]));
assign Uyw7v6 = (~(N6l7x6 & U6l7x6));
assign U6l7x6 = (B7l7x6 | Fsliw6);
assign N6l7x6 = (I7l7x6 & P7l7x6);
assign I7l7x6 = (~(G5j7z6[59] & Kwhov6));
assign Nyw7v6 = (!W7l7x6);
assign W7l7x6 = (M6j7z6[59] ? K8l7x6 : D8l7x6);
assign K8l7x6 = (~(P7l7x6 & R8l7x6));
assign R8l7x6 = (~(W3hov6 & H44iw6));
assign P7l7x6 = (~(Y8l7x6 & Rxh7x6));
assign Rxh7x6 = (~(E5l7x6 | Bgiov6));
assign E5l7x6 = (~(F9l7x6 & P2j7z6[3]));
assign F9l7x6 = (P2j7z6[1] & U1iov6);
assign Y8l7x6 = (R4hov6 & So2nv6);
assign D8l7x6 = (M9l7x6 & T9l7x6);
assign T9l7x6 = (~(T5hov6 & H44iw6));
assign M9l7x6 = (~(Qkj7z6[59] | Aal7x6));
assign Aal7x6 = (Hal7x6 & Tib7z6[59]);
assign Hal7x6 = (~(Jqj7z6[68] & G5j7z6[59]));
assign Gyw7v6 = (~(Oal7x6 & Val7x6));
assign Val7x6 = (~(G5j7z6[52] & Cbl7x6));
assign Cbl7x6 = (~(G2hov6 & L2miw6));
assign L2miw6 = (Fsliw6 | Cshov6);
assign Zxw7v6 = (!Jbl7x6);
assign Jbl7x6 = (M6j7z6[52] ? Xbl7x6 : Qbl7x6);
assign Xbl7x6 = (~(Ecl7x6 & Oal7x6));
assign Oal7x6 = (~(Lcl7x6 & Uuhov6));
assign Lcl7x6 = (R4hov6 & Scl7x6);
assign Ecl7x6 = (~(X7niw6 & Bl5iw6));
assign Qbl7x6 = (Zcl7x6 & Gdl7x6);
assign Gdl7x6 = (~(S8niw6 & Bl5iw6));
assign Zcl7x6 = (~(Qkj7z6[52] | Ndl7x6));
assign Ndl7x6 = (Udl7x6 & Tib7z6[52]);
assign Udl7x6 = (~(Jqj7z6[61] & G5j7z6[52]));
assign Sxw7v6 = (~(Bel7x6 & Iel7x6));
assign Iel7x6 = (~(G5j7z6[53] & Pel7x6));
assign Pel7x6 = (~(G2hov6 & Qlniw6));
assign Lxw7v6 = (!Wel7x6);
assign Wel7x6 = (M6j7z6[53] ? Kfl7x6 : Dfl7x6);
assign Kfl7x6 = (~(Bel7x6 & Rfl7x6));
assign Rfl7x6 = (~(X7niw6 & Ej5iw6));
assign Bel7x6 = (~(Yfl7x6 & Gnniw6));
assign Yfl7x6 = (R4hov6 & Fgl7x6);
assign Dfl7x6 = (Mgl7x6 & Tgl7x6);
assign Tgl7x6 = (~(S8niw6 & Ej5iw6));
assign Mgl7x6 = (~(Qkj7z6[53] | Ahl7x6));
assign Ahl7x6 = (Hhl7x6 & Tib7z6[53]);
assign Hhl7x6 = (~(Jqj7z6[62] & G5j7z6[53]));
assign Exw7v6 = (~(Ohl7x6 & Vhl7x6));
assign Vhl7x6 = (~(G5j7z6[54] & Cil7x6));
assign Cil7x6 = (~(G2hov6 & F6miw6));
assign F6miw6 = (Fsliw6 | Rphov6);
assign Xww7v6 = (!Jil7x6);
assign Jil7x6 = (M6j7z6[54] ? Xil7x6 : Qil7x6);
assign Xil7x6 = (~(Ohl7x6 & Ejl7x6));
assign Ejl7x6 = (~(X7niw6 & D85iw6));
assign Ohl7x6 = (~(Ljl7x6 & Gnhov6));
assign Ljl7x6 = (R4hov6 & Sjl7x6);
assign Qil7x6 = (Zjl7x6 & Gkl7x6);
assign Gkl7x6 = (~(S8niw6 & D85iw6));
assign Zjl7x6 = (~(Qkj7z6[54] | Nkl7x6));
assign Nkl7x6 = (Ukl7x6 & Tib7z6[54]);
assign Ukl7x6 = (~(Jqj7z6[63] & G5j7z6[54]));
assign Qww7v6 = (~(Bll7x6 & Ill7x6));
assign Ill7x6 = (~(G5j7z6[55] & Pll7x6));
assign Pll7x6 = (~(G2hov6 & Rpniw6));
assign Rpniw6 = (J6oiw6 | Fsliw6);
assign G2hov6 = (!Kwhov6);
assign Jww7v6 = (!Wll7x6);
assign Wll7x6 = (M6j7z6[55] ? Kml7x6 : Dml7x6);
assign Kml7x6 = (~(Bll7x6 & Rml7x6));
assign Rml7x6 = (~(X7niw6 & Cx4iw6));
assign X7niw6 = (~(Nmoiw6 | Ie5iw6));
assign Bll7x6 = (~(Orniw6 & Yml7x6));
assign Yml7x6 = (R4hov6 & Fnl7x6);
assign Orniw6 = (Mnl7x6 & P2j7z6[1]);
assign Dml7x6 = (Tnl7x6 & Aol7x6);
assign Aol7x6 = (~(S8niw6 & Cx4iw6));
assign S8niw6 = (~(Dooiw6 | Ie5iw6));
assign Tnl7x6 = (~(Qkj7z6[55] | Hol7x6));
assign Hol7x6 = (Ool7x6 & Tib7z6[55]);
assign Ool7x6 = (~(Jqj7z6[64] & G5j7z6[55]));
assign Cww7v6 = (~(Vol7x6 & Cpl7x6));
assign Cpl7x6 = (~(G5j7z6[60] & Jpl7x6));
assign Jpl7x6 = (Kwhov6 | Mqi7x6);
assign Mqi7x6 = (Qpl7x6 & U4fov6);
assign Vvw7v6 = (!Xpl7x6);
assign Xpl7x6 = (M6j7z6[60] ? Lql7x6 : Eql7x6);
assign Lql7x6 = (~(Sql7x6 & Vol7x6));
assign Vol7x6 = (~(Zql7x6 & R4hov6));
assign Zql7x6 = (C0i7x6 & Grl7x6);
assign Sql7x6 = (~(W3hov6 & W14iw6));
assign Eql7x6 = (Nrl7x6 & Url7x6);
assign Url7x6 = (~(T5hov6 & W14iw6));
assign Nrl7x6 = (~(Qkj7z6[60] | Bsl7x6));
assign Bsl7x6 = (Isl7x6 & Tib7z6[60]);
assign Isl7x6 = (~(Jqj7z6[69] & G5j7z6[60]));
assign Ovw7v6 = (~(Psl7x6 & Wsl7x6));
assign Wsl7x6 = (~(G5j7z6[61] & Dtl7x6));
assign Dtl7x6 = (Kwhov6 | Gui7x6);
assign Gui7x6 = (Ktl7x6 & U4fov6);
assign Kwhov6 = (~(Rtl7x6 & Z3fov6));
assign Z3fov6 = (~(U4fov6 & Sh2nv6));
assign Rtl7x6 = (~(Ytl7x6 & U4fov6));
assign U4fov6 = (!Fsliw6);
assign Hvw7v6 = (!Ful7x6);
assign Ful7x6 = (M6j7z6[61] ? Tul7x6 : Mul7x6);
assign Tul7x6 = (~(Psl7x6 & Avl7x6));
assign Avl7x6 = (~(W3hov6 & Zz3iw6));
assign Psl7x6 = (~(Hvl7x6 & Wvi7x6));
assign Wvi7x6 = (Ovl7x6 & Rc3nv6);
assign Ovl7x6 = (P2j7z6[0] & Rgjov6);
assign Hvl7x6 = (R4hov6 & Vvl7x6);
assign Mul7x6 = (Cwl7x6 & Jwl7x6);
assign Jwl7x6 = (~(T5hov6 & Zz3iw6));
assign Cwl7x6 = (~(Qkj7z6[61] | Qwl7x6));
assign Qwl7x6 = (Xwl7x6 & Tib7z6[61]);
assign Xwl7x6 = (~(Jqj7z6[70] & G5j7z6[61]));
assign Avw7v6 = (~(Exl7x6 & Lxl7x6));
assign Lxl7x6 = (~(Sxl7x6 & Zxl7x6));
assign Zxl7x6 = (~(Jqj7z6[3] & Z3j7z6[1]));
assign Sxl7x6 = (E6a7z6 & Yfdov6);
assign Exl7x6 = (Qlhov6 ? Nyl7x6 : Gyl7x6);
assign Qlhov6 = (~(Uyl7x6 | Nq6iw6));
assign Uyl7x6 = (!Bzl7x6);
assign Nyl7x6 = (~(Izl7x6 & Bk6iw6));
assign Izl7x6 = (Pzl7x6 | Yfdov6);
assign Gyl7x6 = (~(Z3j7z6[14] & Pzl7x6));
assign Tuw7v6 = (~(Wzl7x6 & Pzl7x6));
assign Pzl7x6 = (~(D0m7x6 & Vzgov6));
assign Vzgov6 = (~(Ga3nv6 | K0m7x6));
assign D0m7x6 = (Gnniw6 & R0m7x6);
assign Wzl7x6 = (Z3j7z6[1] ? F1m7x6 : Y0m7x6);
assign F1m7x6 = (~(M1m7x6 & T1m7x6));
assign T1m7x6 = (~(Qlniw6 & A2m7x6));
assign A2m7x6 = (Fsliw6 | Kphov6);
assign Kphov6 = (Sugov6 & H2m7x6);
assign Qlniw6 = (I2oiw6 | Fsliw6);
assign Fsliw6 = (Dtjiw6 & B52nv6);
assign Dtjiw6 = (O2m7x6 & V2m7x6);
assign V2m7x6 = (C3m7x6 & J3m7x6);
assign J3m7x6 = (Q3m7x6 & Bqi7z6[0]);
assign Q3m7x6 = (Bl5iw6 & Gr5iw6);
assign C3m7x6 = (X3m7x6 & Wagiw6);
assign X3m7x6 = (Bqi7z6[3] & Bqi7z6[1]);
assign O2m7x6 = (E4m7x6 & L4m7x6);
assign L4m7x6 = (S4m7x6 & Z4m7x6);
assign S4m7x6 = (Fcgiw6 & Sufiw6);
assign E4m7x6 = (G5m7x6 & T68iw6);
assign G5m7x6 = (Zy4iw6 & N5m7x6);
assign M1m7x6 = (~(L19iw6 & Wohov6));
assign Y0m7x6 = (~(Wohov6 & B52nv6));
assign Wohov6 = (Bzl7x6 & Bqi7z6[0]);
assign Muw7v6 = (~(U5m7x6 & B6m7x6));
assign B6m7x6 = (~(Byi7z6[1] & I6m7x6));
assign I6m7x6 = (~(P6m7x6 & W6m7x6));
assign P6m7x6 = (Bqi7z6[0] & B52nv6);
assign Fuw7v6 = (~(D7m7x6 & K7m7x6));
assign K7m7x6 = (~(R7m7x6 & Y7m7x6));
assign R7m7x6 = (~(Xsinv6 | F8m7x6));
assign D7m7x6 = (~(Byi7z6[31] & M8m7x6));
assign M8m7x6 = (~(W6m7x6 & Gg2iw6));
assign Ytw7v6 = (~(T8m7x6 & A9m7x6));
assign A9m7x6 = (~(H9m7x6 & Etinv6));
assign H9m7x6 = (~(O9m7x6 | Y7m7x6));
assign Y7m7x6 = (Ffadt6 & V9m7x6);
assign T8m7x6 = (~(Byi7z6[30] & Cam7x6));
assign Cam7x6 = (~(W6m7x6 & Nf3iw6));
assign W6m7x6 = (Kgbiw6 & T68iw6);
assign Kgbiw6 = (Eec7x6 & Toi7z6[2]);
assign Rtw7v6 = (!Jam7x6);
assign Jam7x6 = (M6j7z6[62] ? Xam7x6 : Qam7x6);
assign Xam7x6 = (~(Pvhov6 & Ebm7x6));
assign Ebm7x6 = (~(W3hov6 & Ro3iw6));
assign W3hov6 = (~(Nmoiw6 | Dv3iw6));
assign Nmoiw6 = (~(Feeiw6 & G0k7x6));
assign Feeiw6 = (Toi7z6[2] & Toi7z6[7]);
assign Pvhov6 = (~(Lbm7x6 & Y4i7x6));
assign Y4i7x6 = (Sbm7x6 & Rc3nv6);
assign Sbm7x6 = (P2j7z6[1] & Bgiov6);
assign Lbm7x6 = (R4hov6 & Zbm7x6);
assign R4hov6 = (Gcm7x6 & Ncm7x6);
assign Ncm7x6 = (E7iov6 & Owjov6);
assign Gcm7x6 = (Sa2nv6 & P2j7z6[6]);
assign Qam7x6 = (Ucm7x6 & Bdm7x6);
assign Bdm7x6 = (~(T5hov6 & Ro3iw6));
assign T5hov6 = (~(Dooiw6 | Dv3iw6));
assign Dooiw6 = (~(Meeiw6 & G0k7x6));
assign G0k7x6 = (Teeiw6 & Idm7x6);
assign Idm7x6 = (Toi7z6[9] & Hfeiw6);
assign Hfeiw6 = (!Toi7z6[8]);
assign Teeiw6 = (~(Pdm7x6 | X88iw6));
assign X88iw6 = (!Wdm7x6);
assign Meeiw6 = (Toi7z6[2] & D2k7x6);
assign Ucm7x6 = (~(Qkj7z6[62] | Dem7x6));
assign Dem7x6 = (Kem7x6 & Tib7z6[62]);
assign Kem7x6 = (~(Jqj7z6[71] & G5j7z6[62]));
assign Ktw7v6 = (Rem7x6 ? Gvd7z6[0] : Vjc7z6[1]);
assign Dtw7v6 = (Rem7x6 ? Gvd7z6[6] : Vjc7z6[31]);
assign Wsw7v6 = (Rem7x6 ? Gvd7z6[5] : Vjc7z6[6]);
assign Psw7v6 = (Rem7x6 ? Gvd7z6[4] : Vjc7z6[5]);
assign Isw7v6 = (Rem7x6 ? Gvd7z6[3] : Vjc7z6[4]);
assign Bsw7v6 = (Rem7x6 ? Gvd7z6[2] : Vjc7z6[3]);
assign Urw7v6 = (Rem7x6 ? Gvd7z6[1] : Vjc7z6[2]);
assign Nrw7v6 = (~(Yem7x6 & Ffm7x6));
assign Ffm7x6 = (~(Ebdiw6 & Zhg7x6));
assign Yem7x6 = (Mfm7x6 & Tfm7x6);
assign Tfm7x6 = (~(Agm7x6 & Hgm7x6));
assign Hgm7x6 = (~(Ogm7x6 & Rkg7x6));
assign Rkg7x6 = (Vgm7x6 | Chm7x6);
assign Vgm7x6 = (~(Eofov6 & Jhm7x6));
assign Jhm7x6 = (~(Zamov6 & Vs9ov6));
assign Ogm7x6 = (Qhm7x6 | Rd2nv6);
assign Rd2nv6 = (~(Zgadt6 & Xhm7x6));
assign Xhm7x6 = (~(Zamov6 & Ga3nv6));
assign Qhm7x6 = (~(Q7hov6 & Eim7x6));
assign Eim7x6 = (~(Lim7x6 & Zamov6));
assign Agm7x6 = (Amg7x6 ? Vm2nv6 : Ldo7v6);
assign Vm2nv6 = (!Z3j7z6[8]);
assign Mfm7x6 = (~(Bxi7z6[0] & Sim7x6));
assign Sim7x6 = (~(O8fov6 & U42nv6));
assign Grw7v6 = (~(Zim7x6 & Gjm7x6));
assign Gjm7x6 = (~(Njm7x6 & Fe2nv6));
assign Njm7x6 = (~(F02nv6 | Ykg7x6));
assign Ykg7x6 = (Ujm7x6 & Bkm7x6);
assign Bkm7x6 = (~(Ikm7x6 & Zodet6));
assign Ikm7x6 = (~(Cr97z6 | Yfadt6));
assign Ujm7x6 = (~(Sa2nv6 & Jnfov6));
assign Jnfov6 = (~(Pkm7x6 & Wkm7x6));
assign Wkm7x6 = (Dlm7x6 & Klm7x6);
assign Klm7x6 = (~(Rlm7x6 & Ylm7x6));
assign Ylm7x6 = (W2eet6 & Fmm7x6);
assign Fmm7x6 = (Byi7z6[1] | Byi7z6[30]);
assign Rlm7x6 = (Mmm7x6 & Mjniw6);
assign Dlm7x6 = (Tmm7x6 & Anm7x6);
assign Anm7x6 = (~(Hnm7x6 & Onm7x6));
assign Onm7x6 = (Tnzdt6 & Vnm7x6);
assign Vnm7x6 = (~(Com7x6 & Jom7x6));
assign Jom7x6 = (~(Qom7x6 & Mjniw6));
assign Mjniw6 = (~(Qroiw6 | Rgjov6));
assign Qroiw6 = (~(Xom7x6 & P2j7z6[0]));
assign Qom7x6 = (Byi7z6[1] & Dc3nv6);
assign Com7x6 = (~(Epm7x6 & Dc3nv6));
assign Epm7x6 = (Lpm7x6 & Rgjov6);
assign Lpm7x6 = (~(Spm7x6 & Zpm7x6));
assign Zpm7x6 = (~(Mnl7x6 & Gqm7x6));
assign Gqm7x6 = (Bzi7z6[11] | Bzi7z6[12]);
assign Spm7x6 = (~(Nqm7x6 & Uqm7x6));
assign Uqm7x6 = (Bzi7z6[3] | Bzi7z6[4]);
assign Hnm7x6 = (Fe2nv6 & X0eet6);
assign Tmm7x6 = (~(Brm7x6 & Irm7x6));
assign Irm7x6 = (Brdet6 & Prm7x6);
assign Prm7x6 = (Bzi7z6[0] | Bzi7z6[1]);
assign Brm7x6 = (Mmm7x6 & Uuhov6);
assign Uuhov6 = (Nqm7x6 & Rgjov6);
assign Pkm7x6 = (Wrm7x6 & Dsm7x6);
assign Dsm7x6 = (~(Ksm7x6 & Rsm7x6));
assign Rsm7x6 = (Yydet6 & Ysm7x6);
assign Ysm7x6 = (Ftm7x6 | Bzi7z6[10]);
assign Ftm7x6 = (Bzi7z6[8] | Bzi7z6[9]);
assign Ksm7x6 = (Mmm7x6 & Gnniw6);
assign Gnniw6 = (Mnl7x6 & Rgjov6);
assign Mnl7x6 = (Mtm7x6 & P2j7z6[0]);
assign Mtm7x6 = (P2j7z6[2] & Z7iov6);
assign Wrm7x6 = (~(Ttm7x6 & Mmm7x6));
assign Mmm7x6 = (Aum7x6 & Fe2nv6);
assign Aum7x6 = (Dc3nv6 & Tnzdt6);
assign Ttm7x6 = (Gnhov6 & Hum7x6);
assign Hum7x6 = (~(Oum7x6 & Vum7x6));
assign Vum7x6 = (~(Bzi7z6[19] & Zsdet6));
assign Oum7x6 = (Cvm7x6 & Jvm7x6);
assign Jvm7x6 = (~(Zudet6 & Qvm7x6));
assign Qvm7x6 = (Bzi7z6[25] | Bzi7z6[24]);
assign Cvm7x6 = (~(Ywdet6 & Xvm7x6));
assign Xvm7x6 = (Ewm7x6 | Bzi7z6[16]);
assign Ewm7x6 = (Bzi7z6[17] | Bzi7z6[18]);
assign Gnhov6 = (Nqm7x6 & P2j7z6[1]);
assign Nqm7x6 = (Lwm7x6 & P2j7z6[2]);
assign Lwm7x6 = (Bgiov6 & Z7iov6);
assign Zim7x6 = (~(Bxi7z6[3] & Swm7x6));
assign Swm7x6 = (~(O8fov6 & P52nv6));
assign Zqw7v6 = (~(Zwm7x6 & Gxm7x6));
assign Gxm7x6 = (~(Nxm7x6 & Nxeov6));
assign Zwm7x6 = (Uxm7x6 & Bym7x6);
assign Bym7x6 = (~(Sriiw6 & Iym7x6));
assign Iym7x6 = (~(Fjadt6 & Pym7x6));
assign Uxm7x6 = (~(Fjb7z6[1] & Lriiw6));
assign Sqw7v6 = (~(Wym7x6 & Dzm7x6));
assign Dzm7x6 = (Kzm7x6 & Rzm7x6);
assign Rzm7x6 = (~(J6bov6 & Alf7z6[1]));
assign J6bov6 = (Yzm7x6 & F0n7x6);
assign F0n7x6 = (!C6bov6);
assign Kzm7x6 = (~(C6bov6 & Se2jw6));
assign Se2jw6 = (~(M0n7x6 & T0n7x6));
assign T0n7x6 = (~(A1n7x6 & H1n7x6));
assign H1n7x6 = (~(O1n7x6 & V1n7x6));
assign V1n7x6 = (C2n7x6 & J2n7x6);
assign J2n7x6 = (A1v6x6 | J2v6x6);
assign J2v6x6 = (Q2n7x6 & X2n7x6);
assign X2n7x6 = (E3n7x6 & L3n7x6);
assign L3n7x6 = (Mkw6x6 | Vf27x6);
assign Vf27x6 = (Sx07x6 & Kf07x6);
assign Kf07x6 = (S3n7x6 & Z3n7x6);
assign Z3n7x6 = (~(Cve7z6[11] & Sb17x6));
assign S3n7x6 = (~(Cve7z6[27] & Kbx6x6));
assign Sx07x6 = (G4n7x6 & N4n7x6);
assign N4n7x6 = (~(Cve7z6[3] & We07x6));
assign G4n7x6 = (~(Cve7z6[19] & Dbx6x6));
assign E3n7x6 = (~(Xzx6x6 & U4n7x6));
assign U4n7x6 = (~(Id17x6 & Yk27x6));
assign Yk27x6 = (B5n7x6 & I5n7x6);
assign I5n7x6 = (~(Cve7z6[15] & Sb17x6));
assign B5n7x6 = (~(Kbx6x6 & Neo7v6));
assign Id17x6 = (P5n7x6 & W5n7x6);
assign W5n7x6 = (~(Cve7z6[7] & We07x6));
assign P5n7x6 = (~(Cve7z6[23] & Dbx6x6));
assign Q2n7x6 = (D6n7x6 & K6n7x6);
assign K6n7x6 = (E1x6x6 | Hwz6x6);
assign Hwz6x6 = (R6n7x6 & Vzw6x6);
assign Vzw6x6 = (Y6n7x6 & F7n7x6);
assign F7n7x6 = (~(Cve7z6[22] & Sb17x6));
assign Y6n7x6 = (~(Cve7z6[6] & Kbx6x6));
assign R6n7x6 = (Vh07x6 & M7n7x6);
assign M7n7x6 = (~(Cve7z6[30] & We07x6));
assign Vh07x6 = (~(Cve7z6[14] & Dbx6x6));
assign D6n7x6 = (Juv6x6 | Lh27x6);
assign Lh27x6 = (T7n7x6 & Svv6x6);
assign Svv6x6 = (A8n7x6 & H8n7x6);
assign H8n7x6 = (~(Cve7z6[18] & Sb17x6));
assign A8n7x6 = (~(Cve7z6[2] & Kbx6x6));
assign T7n7x6 = (Hh07x6 & O8n7x6);
assign O8n7x6 = (~(Cve7z6[26] & We07x6));
assign Hh07x6 = (~(Cve7z6[10] & Dbx6x6));
assign A1v6x6 = (~(V8n7x6 & C9n7x6));
assign C2n7x6 = (Q2v6x6 | V8v6x6);
assign V8v6x6 = (J9n7x6 & Q9n7x6);
assign Q9n7x6 = (X9n7x6 & Ean7x6);
assign Ean7x6 = (Juv6x6 | Kk27x6);
assign Kk27x6 = (Lan7x6 & Cxz6x6);
assign Cxz6x6 = (San7x6 & Zan7x6);
assign Zan7x6 = (~(Cve7z6[19] & Sb17x6));
assign Cve7z6[19] = (Dte7z6[9] & Fhc7z6[19]);
assign San7x6 = (~(Cve7z6[3] & Kbx6x6));
assign Cve7z6[3] = (Dte7z6[9] & E3c7z6[3]);
assign Lan7x6 = (Y807x6 & Gbn7x6);
assign Gbn7x6 = (~(Cve7z6[27] & We07x6));
assign Cve7z6[27] = (Dte7z6[9] & Fhc7z6[27]);
assign Y807x6 = (~(Cve7z6[11] & Dbx6x6));
assign Cve7z6[11] = (Dte7z6[9] & Fhc7z6[11]);
assign X9n7x6 = (E1x6x6 | Ex07x6);
assign Ex07x6 = (Nbn7x6 & J7x6x6);
assign J7x6x6 = (Ubn7x6 & Bcn7x6);
assign Bcn7x6 = (~(Cve7z6[23] & Sb17x6));
assign Cve7z6[23] = (Dte7z6[9] & Fhc7z6[23]);
assign Ubn7x6 = (~(Cve7z6[7] & Kbx6x6));
assign Cve7z6[7] = (Dte7z6[9] & Fhc7z6[7]);
assign Nbn7x6 = (Af27x6 & Icn7x6);
assign Icn7x6 = (~(We07x6 & Neo7v6));
assign Af27x6 = (~(Cve7z6[15] & Dbx6x6));
assign Cve7z6[15] = (Dte7z6[9] & Fhc7z6[15]);
assign J9n7x6 = (Pcn7x6 & Wcn7x6);
assign Wcn7x6 = (Mkw6x6 | Pj27x6);
assign Pj27x6 = (K017x6 & N607x6);
assign N607x6 = (Ddn7x6 & Kdn7x6);
assign Kdn7x6 = (~(Cve7z6[12] & Sb17x6));
assign Ddn7x6 = (~(Cve7z6[28] & Kbx6x6));
assign K017x6 = (Rdn7x6 & Ydn7x6);
assign Ydn7x6 = (~(Cve7z6[4] & We07x6));
assign Rdn7x6 = (~(Cve7z6[20] & Dbx6x6));
assign Pcn7x6 = (~(Xzx6x6 & Jw07x6));
assign Jw07x6 = (~(Zi17x6 & Pq27x6));
assign Pq27x6 = (Fen7x6 & Men7x6);
assign Men7x6 = (~(Sb17x6 & Cve7z6[16]));
assign Fen7x6 = (~(Cve7z6[0] & Kbx6x6));
assign Zi17x6 = (Ten7x6 & Afn7x6);
assign Afn7x6 = (~(Cve7z6[8] & We07x6));
assign Ten7x6 = (~(Cve7z6[24] & Dbx6x6));
assign Q2v6x6 = (C9n7x6 | V8n7x6);
assign V8n7x6 = (!Hfn7x6);
assign O1n7x6 = (Ofn7x6 & Vfn7x6);
assign Vfn7x6 = (C2v6x6 | C9v6x6);
assign C9v6x6 = (Cgn7x6 & Jgn7x6);
assign Jgn7x6 = (~(Vlw6x6 & Bq27x6));
assign Bq27x6 = (~(Qgn7x6 & Tkw6x6));
assign Tkw6x6 = (Xgn7x6 & Ehn7x6);
assign Ehn7x6 = (~(Cve7z6[20] & Sb17x6));
assign Cve7z6[20] = (Dte7z6[9] & Fhc7z6[20]);
assign Xgn7x6 = (~(Cve7z6[4] & Kbx6x6));
assign Cve7z6[4] = (Dte7z6[9] & E3c7z6[4]);
assign Qgn7x6 = (Zc07x6 & Lhn7x6);
assign Lhn7x6 = (~(Cve7z6[28] & We07x6));
assign Cve7z6[28] = (Dte7z6[9] & Fhc7z6[28]);
assign Zc07x6 = (~(Cve7z6[12] & Dbx6x6));
assign Cve7z6[12] = (Dte7z6[9] & Fhc7z6[12]);
assign Cgn7x6 = (Shn7x6 & Zhn7x6);
assign Zhn7x6 = (Lvv6x6 | Bz07x6);
assign Lvv6x6 = (!Xzx6x6);
assign Shn7x6 = (~(Zvv6x6 & Wz07x6));
assign Wz07x6 = (~(Ja17x6 & Ui27x6));
assign Ui27x6 = (Gin7x6 & Nin7x6);
assign Nin7x6 = (~(Cve7z6[0] & We07x6));
assign Cve7z6[0] = (Dte7z6[9] & E3c7z6[0]);
assign Gin7x6 = (~(Cve7z6[16] & Dbx6x6));
assign Cve7z6[16] = (Dte7z6[9] & Fhc7z6[16]);
assign Ja17x6 = (Uin7x6 & Bjn7x6);
assign Bjn7x6 = (~(Cve7z6[24] & Sb17x6));
assign Cve7z6[24] = (Dte7z6[9] & Fhc7z6[24]);
assign Uin7x6 = (~(Cve7z6[8] & Kbx6x6));
assign Cve7z6[8] = (Dte7z6[9] & Fhc7z6[8]);
assign C2v6x6 = (C9n7x6 | Hfn7x6);
assign Ofn7x6 = (M0v6x6 | X2v6x6);
assign X2v6x6 = (Ijn7x6 & Pjn7x6);
assign Pjn7x6 = (Wjn7x6 & Dkn7x6);
assign Dkn7x6 = (Mkw6x6 | Y2z6x6);
assign Y2z6x6 = (U517x6 & Ha07x6);
assign Ha07x6 = (Kkn7x6 & Rkn7x6);
assign Rkn7x6 = (~(Cve7z6[10] & Sb17x6));
assign Cve7z6[10] = (Dte7z6[9] & Fhc7z6[10]);
assign Kkn7x6 = (~(Cve7z6[26] & Kbx6x6));
assign Cve7z6[26] = (Dte7z6[9] & Fhc7z6[26]);
assign U517x6 = (Ykn7x6 & Fln7x6);
assign Fln7x6 = (~(Cve7z6[2] & We07x6));
assign Cve7z6[2] = (Dte7z6[9] & E3c7z6[2]);
assign Ykn7x6 = (~(Cve7z6[18] & Dbx6x6));
assign Cve7z6[18] = (Dte7z6[9] & Fhc7z6[18]);
assign Mkw6x6 = (!V307x6);
assign V307x6 = (~(Fwbov6 | Cnv6x6));
assign Wjn7x6 = (~(Xzx6x6 & Mln7x6));
assign Mln7x6 = (~(I617x6 & Xg27x6));
assign Xg27x6 = (Tln7x6 & Amn7x6);
assign Amn7x6 = (~(Cve7z6[14] & Sb17x6));
assign Cve7z6[14] = (Dte7z6[9] & Fhc7z6[14]);
assign Tln7x6 = (~(Cve7z6[30] & Kbx6x6));
assign Cve7z6[30] = (Dte7z6[9] & Fhc7z6[30]);
assign I617x6 = (Hmn7x6 & Omn7x6);
assign Omn7x6 = (~(Cve7z6[6] & We07x6));
assign Cve7z6[6] = (Dte7z6[9] & Fhc7z6[6]);
assign Hmn7x6 = (~(Cve7z6[22] & Dbx6x6));
assign Cve7z6[22] = (Dte7z6[9] & Fhc7z6[22]);
assign Xzx6x6 = (~(Fwbov6 | Zuw6x6));
assign Ijn7x6 = (Vmn7x6 & Cnn7x6);
assign Cnn7x6 = (E1x6x6 | Quv6x6);
assign Quv6x6 = (Jnn7x6 & Asw6x6);
assign Asw6x6 = (Qnn7x6 & Xnn7x6);
assign Xnn7x6 = (~(Cve7z6[21] & Sb17x6));
assign Cve7z6[21] = (Dte7z6[9] & Fhc7z6[21]);
assign Qnn7x6 = (~(Cve7z6[5] & Kbx6x6));
assign Cve7z6[5] = (Dte7z6[9] & Fhc7z6[5]);
assign Jnn7x6 = (X407x6 & Eon7x6);
assign Eon7x6 = (~(Cve7z6[29] & We07x6));
assign Cve7z6[29] = (Dte7z6[9] & Fhc7z6[29]);
assign X407x6 = (~(Cve7z6[13] & Dbx6x6));
assign Cve7z6[13] = (Dte7z6[9] & Fhc7z6[13]);
assign E1x6x6 = (!Zvv6x6);
assign Zvv6x6 = (~(Lon7x6 | Cnv6x6));
assign Vmn7x6 = (Juv6x6 | A4z6x6);
assign A4z6x6 = (Son7x6 & Bz07x6);
assign Bz07x6 = (Zon7x6 & Gpn7x6);
assign Gpn7x6 = (~(Cve7z6[17] & Sb17x6));
assign Cve7z6[17] = (Dte7z6[9] & Fhc7z6[17]);
assign Zon7x6 = (~(Cve7z6[1] & Kbx6x6));
assign Cve7z6[1] = (Dte7z6[9] & E3c7z6[1]);
assign Son7x6 = (J407x6 & Npn7x6);
assign Npn7x6 = (~(Cve7z6[25] & We07x6));
assign We07x6 = (~(Upn7x6 | Bqn7x6));
assign Cve7z6[25] = (Dte7z6[9] & Fhc7z6[25]);
assign J407x6 = (~(Cve7z6[9] & Dbx6x6));
assign Cve7z6[9] = (Dte7z6[9] & Fhc7z6[9]);
assign Juv6x6 = (!Vlw6x6);
assign Vlw6x6 = (~(Zuw6x6 | Lon7x6));
assign M0v6x6 = (~(C9n7x6 & Hfn7x6));
assign Hfn7x6 = (~(Vkx6x6 ^ Lon7x6));
assign C9n7x6 = (Fwbov6 ^ Iqn7x6);
assign A1n7x6 = (~(Dzu6x6 ^ Pqn7x6));
assign M0n7x6 = (~(Xrbov6 & Wqn7x6));
assign Wqn7x6 = (Dzu6x6 | Pqn7x6);
assign Pqn7x6 = (Drn7x6 & Eav6x6);
assign Eav6x6 = (~(Krn7x6 | Rbx6x6));
assign Rbx6x6 = (~(Rrn7x6 & Okx6x6));
assign Okx6x6 = (~(Dbx6x6 & Zav6x6));
assign Dbx6x6 = (Upn7x6 & Yrn7x6);
assign Rrn7x6 = (~(Ajy6x6 | Sb17x6));
assign Sb17x6 = (Bqn7x6 & Fsn7x6);
assign Ajy6x6 = (Kbx6x6 & Zav6x6);
assign Krn7x6 = (~(Vfv6x6 & Py17x6));
assign Py17x6 = (Zav6x6 | Kbx6x6);
assign Vfv6x6 = (Msn7x6 & Wubov6);
assign Msn7x6 = (Tsn7x6 & Atn7x6);
assign Drn7x6 = (Zav6x6 ? Qgv6x6 : Kuz6x6);
assign Qgv6x6 = (Sav6x6 & Vkx6x6);
assign Sav6x6 = (Zuw6x6 & Iqn7x6);
assign Dzu6x6 = (~(Htn7x6 & Wubov6));
assign Wubov6 = (Otn7x6 & Vtn7x6);
assign Vtn7x6 = (~(Cun7x6 & Jun7x6));
assign Jun7x6 = (Tsn7x6 & Fwbov6);
assign Fwbov6 = (!Lon7x6);
assign Cun7x6 = (~(Ntbov6 | Kvbov6));
assign Otn7x6 = (~(Lsbov6 & Utbov6));
assign Lsbov6 = (Kvbov6 & Tsn7x6);
assign Tsn7x6 = (~(Dte7z6[6] & Dte7z6[7]));
assign Htn7x6 = (Atn7x6 & Zav6x6);
assign Zav6x6 = (~(Lon7x6 & Ntbov6));
assign Ntbov6 = (~(Kbx6x6 & Yt07x6));
assign Yt07x6 = (Kuz6x6 & Jry6x6);
assign Jry6x6 = (!Vkx6x6);
assign Vkx6x6 = (~(Qun7x6 & Xun7x6));
assign Xun7x6 = (~(Dte7z6[11] & Kxb7z6[0]));
assign Qun7x6 = (~(Ple7z6[0] & Dte7z6[10]));
assign Kuz6x6 = (Evn7x6 & Cnv6x6);
assign Cnv6x6 = (!Zuw6x6);
assign Zuw6x6 = (~(Lvn7x6 & Svn7x6));
assign Svn7x6 = (~(Dte7z6[11] & Kxb7z6[2]));
assign Lvn7x6 = (~(Ple7z6[2] & Dte7z6[10]));
assign Evn7x6 = (!Iqn7x6);
assign Iqn7x6 = (~(Zvn7x6 & Gwn7x6));
assign Gwn7x6 = (~(Dte7z6[11] & Kxb7z6[1]));
assign Zvn7x6 = (~(Ple7z6[1] & Dte7z6[10]));
assign Kbx6x6 = (Bqn7x6 & Upn7x6);
assign Upn7x6 = (!Fsn7x6);
assign Fsn7x6 = (~(Nwn7x6 & Uwn7x6));
assign Uwn7x6 = (~(Dte7z6[11] & Kxb7z6[4]));
assign Nwn7x6 = (~(Ple7z6[4] & Dte7z6[10]));
assign Bqn7x6 = (!Yrn7x6);
assign Yrn7x6 = (~(Bxn7x6 & Ixn7x6));
assign Ixn7x6 = (~(Dte7z6[11] & Kxb7z6[3]));
assign Bxn7x6 = (~(Ple7z6[3] & Dte7z6[10]));
assign Atn7x6 = (~(Lon7x6 & Utbov6));
assign Utbov6 = (~(Pxn7x6 & Zsbov6));
assign Zsbov6 = (Wxn7x6 & Dyn7x6);
assign Dyn7x6 = (~(Dte7z6[11] & Kyn7x6));
assign Kyn7x6 = (Kxb7z6[6] | Kxb7z6[7]);
assign Wxn7x6 = (~(Dte7z6[10] & Ryn7x6));
assign Ryn7x6 = (Ple7z6[6] | Ple7z6[7]);
assign Pxn7x6 = (Yyn7x6 & Fzn7x6);
assign Fzn7x6 = (~(Ple7z6[5] & Dte7z6[10]));
assign Yyn7x6 = (~(Dte7z6[11] & Kxb7z6[5]));
assign Lon7x6 = (~(Dte7z6[7] | Dte7z6[6]));
assign Xrbov6 = (!Byu6x6);
assign Byu6x6 = (~(Mzn7x6 & Dte7z6[7]));
assign Mzn7x6 = (Neo7v6 & Tzn7x6);
assign Tzn7x6 = (!Dte7z6[6]);
assign C6bov6 = (M1lhw6 | Qf2ov6);
assign M1lhw6 = (Y3bov6 & Rfkov6);
assign Rfkov6 = (!Mpe7z6[5]);
assign Wym7x6 = (A0o7x6 & H0o7x6);
assign H0o7x6 = (~(L0g7z6[17] & E7bov6));
assign A0o7x6 = (~(L0g7z6[1] & L7bov6));
assign Lqw7v6 = (O0o7x6 ? Aw77z6 : Bni7z6[1]);
assign Eqw7v6 = (O0o7x6 ? Um77z6 : Bni7z6[31]);
assign Xpw7v6 = (O0o7x6 ? Cn77z6 : Bni7z6[30]);
assign Qpw7v6 = (O0o7x6 ? Kn77z6 : Bni7z6[29]);
assign Jpw7v6 = (O0o7x6 ? Sn77z6 : Bni7z6[28]);
assign Cpw7v6 = (O0o7x6 ? Ao77z6 : Bni7z6[27]);
assign Vow7v6 = (O0o7x6 ? Io77z6 : Bni7z6[26]);
assign Oow7v6 = (O0o7x6 ? Qo77z6 : Bni7z6[25]);
assign How7v6 = (O0o7x6 ? Yo77z6 : Bni7z6[24]);
assign Aow7v6 = (O0o7x6 ? Gp77z6 : Bni7z6[23]);
assign Tnw7v6 = (O0o7x6 ? Op77z6 : Bni7z6[22]);
assign Mnw7v6 = (O0o7x6 ? Wp77z6 : Bni7z6[21]);
assign Fnw7v6 = (O0o7x6 ? Eq77z6 : Bni7z6[20]);
assign Ymw7v6 = (O0o7x6 ? Mq77z6 : Bni7z6[19]);
assign Rmw7v6 = (O0o7x6 ? Uq77z6 : Bni7z6[18]);
assign Kmw7v6 = (O0o7x6 ? Cr77z6 : Bni7z6[17]);
assign Dmw7v6 = (O0o7x6 ? Kr77z6 : Bni7z6[16]);
assign Wlw7v6 = (O0o7x6 ? Sr77z6 : Bni7z6[15]);
assign Plw7v6 = (O0o7x6 ? As77z6 : Bni7z6[14]);
assign Ilw7v6 = (O0o7x6 ? Is77z6 : Bni7z6[13]);
assign Blw7v6 = (O0o7x6 ? Qs77z6 : Bni7z6[12]);
assign Ukw7v6 = (O0o7x6 ? Ys77z6 : Bni7z6[11]);
assign Nkw7v6 = (O0o7x6 ? Gt77z6 : Bni7z6[10]);
assign Gkw7v6 = (O0o7x6 ? Ot77z6 : Bni7z6[9]);
assign Zjw7v6 = (O0o7x6 ? Wt77z6 : Bni7z6[8]);
assign Sjw7v6 = (O0o7x6 ? Eu77z6 : Bni7z6[7]);
assign Ljw7v6 = (O0o7x6 ? Mu77z6 : Bni7z6[6]);
assign Ejw7v6 = (O0o7x6 ? Uu77z6 : Bni7z6[5]);
assign Xiw7v6 = (O0o7x6 ? Cv77z6 : Bni7z6[4]);
assign Qiw7v6 = (O0o7x6 ? Kv77z6 : Bni7z6[3]);
assign Jiw7v6 = (O0o7x6 ? Sv77z6 : Bni7z6[2]);
assign O0o7x6 = (~(Wpk8v6 | V0o7x6));
assign V0o7x6 = (C1o7x6 & Jgliw6);
assign C1o7x6 = (~(Kslov6 & J1o7x6));
assign J1o7x6 = (~(F02nv6 & C0wnv6));
assign Wpk8v6 = (Q1o7x6 & X1o7x6);
assign Q1o7x6 = (E2o7x6 & Jgliw6);
assign E2o7x6 = (~(L2o7x6 & Xolhw6));
assign Xolhw6 = (!Z9onv6);
assign Ciw7v6 = (~(S2o7x6 & Z2o7x6));
assign Z2o7x6 = (~(G3o7x6 & Mq4ft6));
assign G3o7x6 = (N3o7x6 & Wdtnv6);
assign N3o7x6 = (Po4ft6 | E9hnv6);
assign S2o7x6 = (~(K6fov6 & Po4ft6));
assign Ohw7v6 = (U3o7x6 ? Zdp7z6[0] : E9hnv6);
assign U3o7x6 = (Kygnv6 & B4o7x6);
assign E9hnv6 = (I4o7x6 & P4o7x6);
assign P4o7x6 = (W4o7x6 & D5o7x6);
assign W4o7x6 = (~(I7p7z6[0] | W22ft6));
assign I4o7x6 = (~(K5o7x6 | Cx5ov6));
assign Hhw7v6 = (Ypinv6 ? Sk4ft6 : R5o7x6);
assign R5o7x6 = (Y5o7x6 & F6o7x6);
assign F6o7x6 = (~(M6o7x6 & T6o7x6));
assign T6o7x6 = (~(I7p7z6[1] & A7o7x6));
assign M6o7x6 = (D5o7x6 | M12ft6);
assign Ahw7v6 = (K94iw6 ? Um4ft6 : H7o7x6);
assign H7o7x6 = (Y5o7x6 & O7o7x6);
assign Tgw7v6 = (~(V7o7x6 & C8o7x6));
assign C8o7x6 = (J8o7x6 & Q8o7x6);
assign J8o7x6 = (~(Lafov6 | Vhw7v6));
assign Vhw7v6 = (X8o7x6 & E9o7x6);
assign E9o7x6 = (HTMDHBURST[0] & L9o7x6);
assign X8o7x6 = (Y5o7x6 & I7p7z6[3]);
assign V7o7x6 = (S9o7x6 & Z9o7x6);
assign S9o7x6 = (~(W94ft6 & Gao7x6));
assign Gao7x6 = (~(Na9ov6 & Nao7x6));
assign Mgw7v6 = (~(Uao7x6 & Bbo7x6));
assign Bbo7x6 = (~(Ibo7x6 & X15ft6));
assign Ibo7x6 = (Pbo7x6 & Wdtnv6);
assign Pbo7x6 = (A05ft6 | Gpgnv6);
assign Gpgnv6 = (Wbo7x6 & O18ov6);
assign Wbo7x6 = (~(Dco7x6 | Cq2ft6));
assign Uao7x6 = (~(K6fov6 & A05ft6));
assign Fgw7v6 = (~(Kco7x6 & Rco7x6));
assign Rco7x6 = (~(Yco7x6 & Gb5ft6));
assign Yco7x6 = (Fdo7x6 & Wdtnv6);
assign Fdo7x6 = (J95ft6 | Rdgnv6);
assign Kco7x6 = (~(K6fov6 & J95ft6));
assign K6fov6 = (~(Fzunv6 | Mdo7x6));
assign Fzunv6 = (Ac77z6 & Pfo7v6);
assign Rfw7v6 = (Tdo7x6 ? Zdp7z6[2] : Rdgnv6);
assign Tdo7x6 = (Kygnv6 & Aeo7x6);
assign Rdgnv6 = (Heo7x6 & Oeo7x6);
assign Oeo7x6 = (Veo7x6 & B4fiw6);
assign Heo7x6 = (Cfo7x6 & Jfo7x6);
assign Kfw7v6 = (~(Qfo7x6 & Xfo7x6));
assign Xfo7x6 = (B4o7x6 | Ego7x6);
assign Dfw7v6 = (~(Lgo7x6 & Sgo7x6));
assign Sgo7x6 = (B1rnv6 | Zgo7x6);
assign Wew7v6 = (~(Gho7x6 & Nho7x6));
assign Nho7x6 = (Aeo7x6 | Uho7x6);
assign Pew7v6 = (~(Bio7x6 & Iio7x6));
assign Iio7x6 = (U0rnv6 | Pio7x6);
assign Iew7v6 = (Ypinv6 ? M55ft6 : Wio7x6);
assign Wio7x6 = (Djo7x6 & Kjo7x6);
assign Djo7x6 = (~(Rjo7x6 & Yjo7x6));
assign Yjo7x6 = (~(Hmp7z6[1] & Fko7x6));
assign Rjo7x6 = (Mko7x6 | Dm2ft6);
assign Bew7v6 = (Alo7x6 ? Tko7x6 : Wlr7z6[1]);
assign Tko7x6 = (~(Hlo7x6 & Olo7x6));
assign Olo7x6 = (Vlo7x6 & Cmo7x6);
assign Cmo7x6 = (~(Jmo7x6 & A97ov6));
assign Vlo7x6 = (~(Qmo7x6 & Ca7ov6));
assign Hlo7x6 = (Xmo7x6 & Eno7x6);
assign Eno7x6 = (~(Lno7x6 & Ja7ov6));
assign Xmo7x6 = (~(Sno7x6 & H97ov6));
assign Udw7v6 = (Alo7x6 ? Zno7x6 : Wlr7z6[2]);
assign Zno7x6 = (~(Goo7x6 & Noo7x6));
assign Noo7x6 = (Uoo7x6 & Bpo7x6);
assign Bpo7x6 = (~(Jmo7x6 & Iz6ov6));
assign Uoo7x6 = (~(Qmo7x6 & K07ov6));
assign Goo7x6 = (Ipo7x6 & Ppo7x6);
assign Ppo7x6 = (~(Lno7x6 & R07ov6));
assign Ipo7x6 = (~(Sno7x6 & Pz6ov6));
assign Ndw7v6 = (Alo7x6 ? Wpo7x6 : Wlr7z6[3]);
assign Wpo7x6 = (~(Dqo7x6 & Kqo7x6));
assign Kqo7x6 = (Rqo7x6 & Yqo7x6);
assign Yqo7x6 = (~(Jmo7x6 & Sb7ov6));
assign Rqo7x6 = (~(Qmo7x6 & Uc7ov6));
assign Dqo7x6 = (Fro7x6 & Mro7x6);
assign Mro7x6 = (~(Lno7x6 & Bd7ov6));
assign Fro7x6 = (~(Sno7x6 & Zb7ov6));
assign Gdw7v6 = (Alo7x6 ? Tro7x6 : Wlr7z6[4]);
assign Tro7x6 = (~(Aso7x6 & Hso7x6));
assign Hso7x6 = (Oso7x6 & Vso7x6);
assign Vso7x6 = (~(Jmo7x6 & U57ov6));
assign Oso7x6 = (~(Qmo7x6 & W67ov6));
assign Aso7x6 = (Cto7x6 & Jto7x6);
assign Jto7x6 = (~(Lno7x6 & D77ov6));
assign Cto7x6 = (~(Sno7x6 & B67ov6));
assign Zcw7v6 = (Alo7x6 ? Qto7x6 : Wlr7z6[5]);
assign Qto7x6 = (~(Xto7x6 & Euo7x6));
assign Euo7x6 = (Luo7x6 & Suo7x6);
assign Suo7x6 = (~(Jmo7x6 & Og7ov6));
assign Luo7x6 = (~(Qmo7x6 & Qh7ov6));
assign Xto7x6 = (Zuo7x6 & Gvo7x6);
assign Gvo7x6 = (~(Lno7x6 & Xh7ov6));
assign Zuo7x6 = (~(Sno7x6 & Vg7ov6));
assign Scw7v6 = (Alo7x6 ? Nvo7x6 : Wlr7z6[6]);
assign Nvo7x6 = (~(Uvo7x6 & Bwo7x6));
assign Bwo7x6 = (Iwo7x6 & Pwo7x6);
assign Pwo7x6 = (~(Jmo7x6 & An7ov6));
assign Iwo7x6 = (~(Qmo7x6 & Co7ov6));
assign Uvo7x6 = (Wwo7x6 & Dxo7x6);
assign Dxo7x6 = (~(Lno7x6 & Jo7ov6));
assign Wwo7x6 = (~(Sno7x6 & Hn7ov6));
assign Lcw7v6 = (Alo7x6 ? Kxo7x6 : Wlr7z6[7]);
assign Kxo7x6 = (~(Rxo7x6 & Yxo7x6));
assign Yxo7x6 = (Fyo7x6 & Myo7x6);
assign Myo7x6 = (~(Qmo7x6 & Ax4ov6));
assign Fyo7x6 = (~(Jmo7x6 & Ox4ov6));
assign Rxo7x6 = (Tyo7x6 & Azo7x6);
assign Azo7x6 = (~(Sno7x6 & Yv4ov6));
assign Tyo7x6 = (~(Lno7x6 & Qy4ov6));
assign Ecw7v6 = (Alo7x6 ? Hzo7x6 : Wlr7z6[8]);
assign Hzo7x6 = (~(Ozo7x6 & Vzo7x6));
assign Vzo7x6 = (C0p7x6 & J0p7x6);
assign J0p7x6 = (~(Q0p7x6 & C37ov6));
assign C0p7x6 = (~(X0p7x6 & H27ov6));
assign Ozo7x6 = (E1p7x6 & L1p7x6);
assign L1p7x6 = (~(S1p7x6 & J37ov6));
assign E1p7x6 = (~(Z1p7x6 & A27ov6));
assign Xbw7v6 = (Alo7x6 ? G2p7x6 : Wlr7z6[9]);
assign G2p7x6 = (~(N2p7x6 & U2p7x6));
assign U2p7x6 = (B3p7x6 & I3p7x6);
assign I3p7x6 = (~(Z1p7x6 & A97ov6));
assign B3p7x6 = (~(Q0p7x6 & Ca7ov6));
assign N2p7x6 = (P3p7x6 & W3p7x6);
assign W3p7x6 = (~(S1p7x6 & Ja7ov6));
assign P3p7x6 = (~(X0p7x6 & H97ov6));
assign Qbw7v6 = (Alo7x6 ? D4p7x6 : Wlr7z6[10]);
assign D4p7x6 = (~(K4p7x6 & R4p7x6));
assign R4p7x6 = (Y4p7x6 & F5p7x6);
assign F5p7x6 = (~(Z1p7x6 & Iz6ov6));
assign Y4p7x6 = (~(Q0p7x6 & K07ov6));
assign K4p7x6 = (M5p7x6 & T5p7x6);
assign T5p7x6 = (~(S1p7x6 & R07ov6));
assign M5p7x6 = (~(X0p7x6 & Pz6ov6));
assign Jbw7v6 = (Alo7x6 ? A6p7x6 : Wlr7z6[11]);
assign A6p7x6 = (~(H6p7x6 & O6p7x6));
assign O6p7x6 = (V6p7x6 & C7p7x6);
assign C7p7x6 = (~(Z1p7x6 & Sb7ov6));
assign V6p7x6 = (~(Q0p7x6 & Uc7ov6));
assign H6p7x6 = (J7p7x6 & Q7p7x6);
assign Q7p7x6 = (~(S1p7x6 & Bd7ov6));
assign J7p7x6 = (~(X0p7x6 & Zb7ov6));
assign Cbw7v6 = (Alo7x6 ? X7p7x6 : Wlr7z6[12]);
assign X7p7x6 = (~(E8p7x6 & L8p7x6));
assign L8p7x6 = (S8p7x6 & Z8p7x6);
assign Z8p7x6 = (~(Z1p7x6 & U57ov6));
assign S8p7x6 = (~(Q0p7x6 & W67ov6));
assign E8p7x6 = (G9p7x6 & N9p7x6);
assign N9p7x6 = (~(S1p7x6 & D77ov6));
assign G9p7x6 = (~(X0p7x6 & B67ov6));
assign Vaw7v6 = (Alo7x6 ? U9p7x6 : Wlr7z6[13]);
assign U9p7x6 = (~(Bap7x6 & Iap7x6));
assign Iap7x6 = (Pap7x6 & Wap7x6);
assign Wap7x6 = (~(Z1p7x6 & Og7ov6));
assign Pap7x6 = (~(Q0p7x6 & Qh7ov6));
assign Bap7x6 = (Dbp7x6 & Kbp7x6);
assign Kbp7x6 = (~(S1p7x6 & Xh7ov6));
assign Dbp7x6 = (~(X0p7x6 & Vg7ov6));
assign Oaw7v6 = (Alo7x6 ? Rbp7x6 : Wlr7z6[14]);
assign Rbp7x6 = (~(Ybp7x6 & Fcp7x6));
assign Fcp7x6 = (Mcp7x6 & Tcp7x6);
assign Tcp7x6 = (~(Z1p7x6 & An7ov6));
assign Mcp7x6 = (~(Q0p7x6 & Co7ov6));
assign Ybp7x6 = (Adp7x6 & Hdp7x6);
assign Hdp7x6 = (~(S1p7x6 & Jo7ov6));
assign Adp7x6 = (~(X0p7x6 & Hn7ov6));
assign Haw7v6 = (Alo7x6 ? Odp7x6 : Wlr7z6[15]);
assign Odp7x6 = (~(Vdp7x6 & Cep7x6));
assign Cep7x6 = (Jep7x6 & Qep7x6);
assign Qep7x6 = (~(Q0p7x6 & Ax4ov6));
assign Jep7x6 = (~(Z1p7x6 & Ox4ov6));
assign Vdp7x6 = (Xep7x6 & Efp7x6);
assign Efp7x6 = (~(X0p7x6 & Yv4ov6));
assign Xep7x6 = (~(S1p7x6 & Qy4ov6));
assign Aaw7v6 = (~(Lfp7x6 & Sfp7x6));
assign Sfp7x6 = (Zfp7x6 & Ggp7x6);
assign Ggp7x6 = (~(Jy4ov6 & A27ov6));
assign Zfp7x6 = (Ngp7x6 & Ugp7x6);
assign Ugp7x6 = (~(Hx4ov6 & H27ov6));
assign Ngp7x6 = (~(Tw4ov6 & J37ov6));
assign Lfp7x6 = (Bhp7x6 & Ihp7x6);
assign Ihp7x6 = (~(Rv4ov6 & C37ov6));
assign Bhp7x6 = (~(Wlr7z6[16] & Xy4ov6));
assign T9w7v6 = (~(Php7x6 & Whp7x6));
assign Whp7x6 = (Dip7x6 & Kip7x6);
assign Kip7x6 = (~(Tw4ov6 & Ja7ov6));
assign Dip7x6 = (Rip7x6 & Yip7x6);
assign Yip7x6 = (~(Jy4ov6 & A97ov6));
assign Rip7x6 = (~(Rv4ov6 & Ca7ov6));
assign Php7x6 = (Fjp7x6 & Mjp7x6);
assign Mjp7x6 = (~(Hx4ov6 & H97ov6));
assign Fjp7x6 = (~(Wlr7z6[17] & Xy4ov6));
assign M9w7v6 = (~(Tjp7x6 & Akp7x6));
assign Akp7x6 = (Hkp7x6 & Okp7x6);
assign Okp7x6 = (~(Tw4ov6 & R07ov6));
assign Hkp7x6 = (Vkp7x6 & Clp7x6);
assign Clp7x6 = (~(Jy4ov6 & Iz6ov6));
assign Vkp7x6 = (~(Rv4ov6 & K07ov6));
assign Tjp7x6 = (Jlp7x6 & Qlp7x6);
assign Qlp7x6 = (~(Hx4ov6 & Pz6ov6));
assign Jlp7x6 = (~(Wlr7z6[18] & Xy4ov6));
assign F9w7v6 = (~(Xlp7x6 & Emp7x6));
assign Emp7x6 = (Lmp7x6 & Smp7x6);
assign Smp7x6 = (~(Tw4ov6 & Bd7ov6));
assign Lmp7x6 = (Zmp7x6 & Gnp7x6);
assign Gnp7x6 = (~(Jy4ov6 & Sb7ov6));
assign Zmp7x6 = (~(Rv4ov6 & Uc7ov6));
assign Xlp7x6 = (Nnp7x6 & Unp7x6);
assign Unp7x6 = (~(Hx4ov6 & Zb7ov6));
assign Nnp7x6 = (~(Wlr7z6[19] & Xy4ov6));
assign Y8w7v6 = (~(Bop7x6 & Iop7x6));
assign Iop7x6 = (Pop7x6 & Wop7x6);
assign Wop7x6 = (~(Tw4ov6 & D77ov6));
assign Pop7x6 = (Dpp7x6 & Kpp7x6);
assign Kpp7x6 = (~(Jy4ov6 & U57ov6));
assign Dpp7x6 = (~(Rv4ov6 & W67ov6));
assign Bop7x6 = (Rpp7x6 & Ypp7x6);
assign Ypp7x6 = (~(Hx4ov6 & B67ov6));
assign Rpp7x6 = (~(Wlr7z6[20] & Xy4ov6));
assign R8w7v6 = (~(Fqp7x6 & Mqp7x6));
assign Mqp7x6 = (Tqp7x6 & Arp7x6);
assign Arp7x6 = (~(Tw4ov6 & Xh7ov6));
assign Tqp7x6 = (Hrp7x6 & Orp7x6);
assign Orp7x6 = (~(Jy4ov6 & Og7ov6));
assign Hrp7x6 = (~(Rv4ov6 & Qh7ov6));
assign Fqp7x6 = (Vrp7x6 & Csp7x6);
assign Csp7x6 = (~(Hx4ov6 & Vg7ov6));
assign Vrp7x6 = (~(Wlr7z6[21] & Xy4ov6));
assign K8w7v6 = (~(Jsp7x6 & Qsp7x6));
assign Qsp7x6 = (Xsp7x6 & Etp7x6);
assign Etp7x6 = (~(Rv4ov6 & Co7ov6));
assign Xsp7x6 = (Ltp7x6 & Stp7x6);
assign Stp7x6 = (~(Jy4ov6 & An7ov6));
assign Ltp7x6 = (~(Hx4ov6 & Hn7ov6));
assign Jsp7x6 = (Ztp7x6 & Gup7x6);
assign Gup7x6 = (~(Tw4ov6 & Jo7ov6));
assign Ztp7x6 = (~(Wlr7z6[22] & Xy4ov6));
assign D8w7v6 = (~(Nup7x6 & Uup7x6));
assign Uup7x6 = (Bvp7x6 & Ivp7x6);
assign Ivp7x6 = (~(Hx4ov6 & Yv4ov6));
assign Yv4ov6 = (~(Pvp7x6 & Wvp7x6));
assign Wvp7x6 = (~(Dwp7x6 & Kwp7x6));
assign Pvp7x6 = (~(Rwp7x6 & Hp67x6));
assign Bvp7x6 = (Ywp7x6 & Fxp7x6);
assign Fxp7x6 = (~(Rv4ov6 & Ax4ov6));
assign Ax4ov6 = (~(Mxp7x6 & Txp7x6));
assign Txp7x6 = (~(Dwp7x6 & Ht1ov6));
assign Mxp7x6 = (~(Rwp7x6 & Kn67x6));
assign Ywp7x6 = (~(Jy4ov6 & Ox4ov6));
assign Ox4ov6 = (~(Ayp7x6 & Hyp7x6));
assign Hyp7x6 = (~(Dwp7x6 & Oyp7x6));
assign Ayp7x6 = (~(Rwp7x6 & Dh57x6));
assign Nup7x6 = (Vyp7x6 & Czp7x6);
assign Czp7x6 = (~(Tw4ov6 & Qy4ov6));
assign Qy4ov6 = (~(Jzp7x6 & Qzp7x6));
assign Qzp7x6 = (~(Dwp7x6 & Xzp7x6));
assign Jzp7x6 = (~(Rwp7x6 & Rh57x6));
assign Vyp7x6 = (~(Wlr7z6[23] & Xy4ov6));
assign W7w7v6 = (~(E0q7x6 & L0q7x6));
assign L0q7x6 = (S0q7x6 & Z0q7x6);
assign Z0q7x6 = (~(Jy4ov6 & J37ov6));
assign S0q7x6 = (G1q7x6 & N1q7x6);
assign N1q7x6 = (~(Hx4ov6 & A27ov6));
assign G1q7x6 = (~(Tw4ov6 & C37ov6));
assign E0q7x6 = (U1q7x6 & B2q7x6);
assign B2q7x6 = (~(Rv4ov6 & H27ov6));
assign U1q7x6 = (~(Wlr7z6[24] & Xy4ov6));
assign P7w7v6 = (~(I2q7x6 & P2q7x6));
assign P2q7x6 = (W2q7x6 & D3q7x6);
assign D3q7x6 = (~(Jy4ov6 & Ja7ov6));
assign Ja7ov6 = (~(K3q7x6 & R3q7x6));
assign R3q7x6 = (~(Dwp7x6 & Y3q7x6));
assign K3q7x6 = (~(Rwp7x6 & Ob67x6));
assign W2q7x6 = (F4q7x6 & M4q7x6);
assign M4q7x6 = (~(Hx4ov6 & A97ov6));
assign A97ov6 = (~(T4q7x6 & A5q7x6));
assign A5q7x6 = (~(Dwp7x6 & H5q7x6));
assign T4q7x6 = (~(Rwp7x6 & Ab67x6));
assign F4q7x6 = (~(Tw4ov6 & Ca7ov6));
assign Ca7ov6 = (~(O5q7x6 & V5q7x6));
assign V5q7x6 = (~(Dwp7x6 & C6q7x6));
assign O5q7x6 = (~(Rwp7x6 & Vv77x6));
assign I2q7x6 = (J6q7x6 & Q6q7x6);
assign Q6q7x6 = (~(Rv4ov6 & H97ov6));
assign H97ov6 = (~(X6q7x6 & E7q7x6));
assign E7q7x6 = (~(Dwp7x6 & L7q7x6));
assign X6q7x6 = (~(Rwp7x6 & Ex77x6));
assign J6q7x6 = (~(Wlr7z6[25] & Xy4ov6));
assign I7w7v6 = (~(S7q7x6 & Z7q7x6));
assign Z7q7x6 = (G8q7x6 & N8q7x6);
assign N8q7x6 = (~(Jy4ov6 & R07ov6));
assign R07ov6 = (~(U8q7x6 & B9q7x6));
assign B9q7x6 = (~(Dwp7x6 & I9q7x6));
assign U8q7x6 = (~(Rwp7x6 & Ddfov6));
assign G8q7x6 = (P9q7x6 & W9q7x6);
assign W9q7x6 = (~(Hx4ov6 & Iz6ov6));
assign Iz6ov6 = (~(Daq7x6 & Kaq7x6));
assign Kaq7x6 = (~(Dwp7x6 & Raq7x6));
assign Daq7x6 = (~(Rwp7x6 & Kdfov6));
assign P9q7x6 = (~(Tw4ov6 & K07ov6));
assign K07ov6 = (~(Yaq7x6 & Fbq7x6));
assign Fbq7x6 = (~(Dwp7x6 & Mbq7x6));
assign Yaq7x6 = (~(Rwp7x6 & Bcfov6));
assign S7q7x6 = (Tbq7x6 & Acq7x6);
assign Acq7x6 = (~(Rv4ov6 & Pz6ov6));
assign Pz6ov6 = (~(Hcq7x6 & Ocq7x6));
assign Ocq7x6 = (~(Dwp7x6 & Vcq7x6));
assign Hcq7x6 = (~(Rwp7x6 & Icfov6));
assign Tbq7x6 = (~(Wlr7z6[26] & Xy4ov6));
assign B7w7v6 = (~(Cdq7x6 & Jdq7x6));
assign Jdq7x6 = (Qdq7x6 & Xdq7x6);
assign Xdq7x6 = (~(Jy4ov6 & Bd7ov6));
assign Bd7ov6 = (~(Eeq7x6 & Leq7x6));
assign Leq7x6 = (~(Dwp7x6 & Seq7x6));
assign Eeq7x6 = (~(Rwp7x6 & Hnlov6));
assign Qdq7x6 = (Zeq7x6 & Gfq7x6);
assign Gfq7x6 = (~(Hx4ov6 & Sb7ov6));
assign Sb7ov6 = (~(Nfq7x6 & Ufq7x6));
assign Ufq7x6 = (~(Dwp7x6 & Bgq7x6));
assign Nfq7x6 = (~(Rwp7x6 & Onlov6));
assign Zeq7x6 = (~(Tw4ov6 & Uc7ov6));
assign Uc7ov6 = (~(Igq7x6 & Pgq7x6));
assign Pgq7x6 = (~(Dwp7x6 & Wgq7x6));
assign Igq7x6 = (~(Rwp7x6 & Fmlov6));
assign Cdq7x6 = (Dhq7x6 & Khq7x6);
assign Khq7x6 = (~(Rv4ov6 & Zb7ov6));
assign Zb7ov6 = (~(Rhq7x6 & Yhq7x6));
assign Yhq7x6 = (~(Dwp7x6 & Fiq7x6));
assign Rhq7x6 = (~(Rwp7x6 & Mmlov6));
assign Dhq7x6 = (~(Wlr7z6[27] & Xy4ov6));
assign U6w7v6 = (~(Miq7x6 & Tiq7x6));
assign Tiq7x6 = (Ajq7x6 & Hjq7x6);
assign Hjq7x6 = (~(Jy4ov6 & D77ov6));
assign D77ov6 = (~(Ojq7x6 & Vjq7x6));
assign Vjq7x6 = (~(Dwp7x6 & Ckq7x6));
assign Ojq7x6 = (~(Rwp7x6 & Ax57x6));
assign Ajq7x6 = (Jkq7x6 & Qkq7x6);
assign Qkq7x6 = (~(Hx4ov6 & U57ov6));
assign U57ov6 = (~(Xkq7x6 & Elq7x6));
assign Elq7x6 = (~(Dwp7x6 & Llq7x6));
assign Xkq7x6 = (~(Rwp7x6 & Tw57x6));
assign Jkq7x6 = (~(Tw4ov6 & W67ov6));
assign W67ov6 = (~(Slq7x6 & Zlq7x6));
assign Zlq7x6 = (~(Dwp7x6 & Gmq7x6));
assign Slq7x6 = (~(Rwp7x6 & T977x6));
assign Miq7x6 = (Nmq7x6 & Umq7x6);
assign Umq7x6 = (~(Rv4ov6 & B67ov6));
assign B67ov6 = (~(Bnq7x6 & Inq7x6));
assign Inq7x6 = (~(Dwp7x6 & Pnq7x6));
assign Bnq7x6 = (~(Rwp7x6 & Cb77x6));
assign Nmq7x6 = (~(Wlr7z6[28] & Xy4ov6));
assign N6w7v6 = (~(Wnq7x6 & Doq7x6));
assign Doq7x6 = (Koq7x6 & Roq7x6);
assign Roq7x6 = (~(Jy4ov6 & Xh7ov6));
assign Xh7ov6 = (~(Yoq7x6 & Fpq7x6));
assign Fpq7x6 = (~(Dwp7x6 & Mpq7x6));
assign Yoq7x6 = (~(Rwp7x6 & Xr57x6));
assign Koq7x6 = (Tpq7x6 & Aqq7x6);
assign Aqq7x6 = (~(Hx4ov6 & Og7ov6));
assign Og7ov6 = (~(Hqq7x6 & Oqq7x6));
assign Oqq7x6 = (~(Dwp7x6 & Vqq7x6));
assign Hqq7x6 = (~(Rwp7x6 & Qr57x6));
assign Tpq7x6 = (~(Tw4ov6 & Qh7ov6));
assign Qh7ov6 = (~(Crq7x6 & Jrq7x6));
assign Jrq7x6 = (~(Dwp7x6 & Qrq7x6));
assign Crq7x6 = (~(Rwp7x6 & T277x6));
assign Wnq7x6 = (Xrq7x6 & Esq7x6);
assign Esq7x6 = (~(Rv4ov6 & Vg7ov6));
assign Vg7ov6 = (~(Lsq7x6 & Ssq7x6));
assign Ssq7x6 = (~(Dwp7x6 & Zsq7x6));
assign Lsq7x6 = (~(Rwp7x6 & C477x6));
assign Xrq7x6 = (~(Wlr7z6[29] & Xy4ov6));
assign G6w7v6 = (~(Gtq7x6 & Ntq7x6));
assign Ntq7x6 = (Utq7x6 & Buq7x6);
assign Buq7x6 = (~(Jy4ov6 & Jo7ov6));
assign Jo7ov6 = (~(Iuq7x6 & Puq7x6));
assign Puq7x6 = (~(Dwp7x6 & Wuq7x6));
assign Iuq7x6 = (~(Rwp7x6 & Um57x6));
assign Jy4ov6 = (Dvq7x6 & Ncp7z6[0]);
assign Dvq7x6 = (Ncp7z6[1] & Kvq7x6);
assign Utq7x6 = (Rvq7x6 & Yvq7x6);
assign Yvq7x6 = (~(Hx4ov6 & An7ov6));
assign An7ov6 = (~(Fwq7x6 & Mwq7x6));
assign Mwq7x6 = (~(Dwp7x6 & Twq7x6));
assign Fwq7x6 = (~(Rwp7x6 & Nm57x6));
assign Hx4ov6 = (Axq7x6 & Ncp7z6[1]);
assign Axq7x6 = (Kvq7x6 & T69ov6);
assign Rvq7x6 = (~(Tw4ov6 & Co7ov6));
assign Co7ov6 = (~(Hxq7x6 & Oxq7x6));
assign Oxq7x6 = (~(Dwp7x6 & Vxq7x6));
assign Hxq7x6 = (~(Rwp7x6 & Tv67x6));
assign Tw4ov6 = (Cyq7x6 & Kvq7x6);
assign Gtq7x6 = (Jyq7x6 & Qyq7x6);
assign Qyq7x6 = (~(Rv4ov6 & Hn7ov6));
assign Hn7ov6 = (~(Xyq7x6 & Ezq7x6));
assign Ezq7x6 = (~(Dwp7x6 & Lzq7x6));
assign Xyq7x6 = (~(Rwp7x6 & Cx67x6));
assign Rv4ov6 = (Szq7x6 & Ncp7z6[0]);
assign Szq7x6 = (Kvq7x6 & M69ov6);
assign Kvq7x6 = (Zzq7x6 & Bbp7z6[1]);
assign Zzq7x6 = (~(Xy4ov6 | Bbp7z6[0]));
assign Jyq7x6 = (~(Wlr7z6[30] & Xy4ov6));
assign Z5w7v6 = (Alo7x6 ? G0r7x6 : Dfr7z6[0]);
assign G0r7x6 = (N0r7x6 & Z9o7x6);
assign N0r7x6 = (~(M55ft6 & U0r7x6));
assign S5w7v6 = (Alo7x6 ? B1r7x6 : Dfr7z6[1]);
assign B1r7x6 = (U0r7x6 & Z9o7x6);
assign L5w7v6 = (Alo7x6 ? L42ft6 : Vr5ft6);
assign E5w7v6 = (Alo7x6 ? Bbp7z6[0] : Xcr7z6[0]);
assign X4w7v6 = (Alo7x6 ? Bbp7z6[1] : Xcr7z6[1]);
assign Q4w7v6 = (Alo7x6 ? I1r7x6 : Wlr7z6[0]);
assign I1r7x6 = (~(P1r7x6 & W1r7x6));
assign W1r7x6 = (D2r7x6 & K2r7x6);
assign K2r7x6 = (~(Qmo7x6 & C37ov6));
assign C37ov6 = (~(R2r7x6 & Y2r7x6));
assign Y2r7x6 = (~(Dwp7x6 & Yqonv6));
assign R2r7x6 = (~(Rwp7x6 & Fd9ov6));
assign Qmo7x6 = (X0p7x6 | F3r7x6);
assign F3r7x6 = (M3r7x6 & Ncp7z6[0]);
assign M3r7x6 = (~(M69ov6 | Bbp7z6[1]));
assign X0p7x6 = (T3r7x6 & Ncp7z6[0]);
assign T3r7x6 = (Ncp7z6[1] & A4r7x6);
assign D2r7x6 = (~(Lno7x6 & J37ov6));
assign J37ov6 = (~(H4r7x6 & O4r7x6));
assign O4r7x6 = (~(Dwp7x6 & V4r7x6));
assign H4r7x6 = (~(Rwp7x6 & Ve9ov6));
assign Lno7x6 = (Q0p7x6 | C5r7x6);
assign C5r7x6 = (J5r7x6 & Ncp7z6[1]);
assign J5r7x6 = (~(Ncp7z6[0] | Bbp7z6[1]));
assign Q0p7x6 = (Q5r7x6 & Ncp7z6[1]);
assign Q5r7x6 = (A4r7x6 & T69ov6);
assign P1r7x6 = (X5r7x6 & E6r7x6);
assign E6r7x6 = (~(Jmo7x6 & A27ov6));
assign A27ov6 = (~(L6r7x6 & S6r7x6));
assign S6r7x6 = (~(Dwp7x6 & Kqonv6));
assign L6r7x6 = (~(Rwp7x6 & Jf9ov6));
assign Jmo7x6 = (S1p7x6 | Z6r7x6);
assign Z6r7x6 = (G7r7x6 & Ncp7z6[0]);
assign S1p7x6 = (N7r7x6 & Ncp7z6[0]);
assign N7r7x6 = (A4r7x6 & M69ov6);
assign X5r7x6 = (~(Sno7x6 & H27ov6));
assign H27ov6 = (~(U7r7x6 & B8r7x6));
assign B8r7x6 = (~(Dwp7x6 & I8r7x6));
assign Dwp7x6 = (~(P8r7x6 | Kygnv6));
assign P8r7x6 = (!L42ft6);
assign U7r7x6 = (~(Rwp7x6 & Td9ov6));
assign Rwp7x6 = (~(Kygnv6 | L42ft6));
assign Sno7x6 = (Z1p7x6 | W8r7x6);
assign W8r7x6 = (G7r7x6 & T69ov6);
assign G7r7x6 = (~(Ncp7z6[1] | Bbp7z6[1]));
assign Z1p7x6 = (Cyq7x6 & A4r7x6);
assign A4r7x6 = (Bbp7z6[0] ^ Bbp7z6[1]);
assign Cyq7x6 = (T69ov6 & M69ov6);
assign M69ov6 = (!Ncp7z6[1]);
assign T69ov6 = (!Ncp7z6[0]);
assign J4w7v6 = (K94iw6 ? O75ft6 : D9r7x6);
assign C4w7v6 = (~(K9r7x6 & Kkg7x6));
assign Kkg7x6 = (~(Ffadt6 & Jg2nv6));
assign Jg2nv6 = (~(R9r7x6 & Y9r7x6));
assign Y9r7x6 = (Far7x6 & Bc2nv6);
assign Bc2nv6 = (~(Mar7x6 & Tar7x6));
assign Tar7x6 = (~(Etinv6 & Abr7x6));
assign Abr7x6 = (~(Uxeov6 & Hbr7x6));
assign Hbr7x6 = (~(Sfoov6 & Obr7x6));
assign Obr7x6 = (~(Vbr7x6 & Ccr7x6));
assign Vbr7x6 = (Jcr7x6 & Qcr7x6);
assign Qcr7x6 = (Xcr7x6 | Mbiov6);
assign Xcr7x6 = (Edr7x6 & Ldr7x6);
assign Jcr7x6 = (Ldr7x6 | Edr7x6);
assign Edr7x6 = (Sdr7x6 & Zdr7x6);
assign Zdr7x6 = (~(Ger7x6 & Ociov6));
assign Sdr7x6 = (~(Ner7x6 & Cdiov6));
assign Ner7x6 = (Uer7x6 & CURRPRI[5]);
assign Uer7x6 = (~(Qdiov6 & Bfr7x6));
assign Sfoov6 = (Fvjov6 & W9iov6);
assign W9iov6 = (K0m7x6 | Rxgov6);
assign Rxgov6 = (~(P2j7z6[1] & Q7niw6));
assign Q7niw6 = (Xom7x6 & Bgiov6);
assign Xom7x6 = (U1iov6 & Z7iov6);
assign K0m7x6 = (!Dc3nv6);
assign Mar7x6 = (Ifr7x6 & Ui2nv6);
assign Ifr7x6 = (~(Pfr7x6 & Ev2nv6));
assign Pfr7x6 = (~(Xg2nv6 & Nxeov6));
assign Far7x6 = (Bj2nv6 & Lh2nv6);
assign Lh2nv6 = (~(Nmadt6 & Wfr7x6));
assign Wfr7x6 = (~(Dgr7x6 & Kgr7x6));
assign Kgr7x6 = (L7iov6 & Rviov6);
assign L7iov6 = (Rgr7x6 & Ygr7x6);
assign Ygr7x6 = (~(Rviov6 & Itjov6));
assign Dgr7x6 = (B2iov6 & G8iov6);
assign G8iov6 = (Fhr7x6 & Mhr7x6);
assign Mhr7x6 = (~(Thr7x6 | Lsiov6));
assign Thr7x6 = (Rviov6 & Air7x6);
assign Air7x6 = (E6jov6 | Hir7x6);
assign Hir7x6 = (Itjov6 & Ptjov6);
assign Fhr7x6 = (Oir7x6 & Vir7x6);
assign Vir7x6 = (Rgr7x6 | Apjov6);
assign Rgr7x6 = (!Tojov6);
assign Oir7x6 = (~(Hsgov6 & D9jov6));
assign B2iov6 = (Cjr7x6 & Jjr7x6);
assign Jjr7x6 = (Qjr7x6 & Xjr7x6);
assign Xjr7x6 = (~(Hsgov6 & Ekr7x6));
assign Ekr7x6 = (Sdjov6 | Lkr7x6);
assign Lkr7x6 = (Skr7x6 & Dnjov6);
assign Sdjov6 = (D9jov6 & Zkr7x6);
assign Qjr7x6 = (~(Sliov6 | Bniov6));
assign Bniov6 = (Glr7x6 & Tojov6);
assign Glr7x6 = (~(Apjov6 | Nlr7x6));
assign Sliov6 = (Ulr7x6 & Bmr7x6);
assign Bmr7x6 = (Cjjov6 & Jjjov6);
assign Ulr7x6 = (Osgov6 & Imr7x6);
assign Imr7x6 = (!Qjjov6);
assign Cjr7x6 = (Pmr7x6 & Wmr7x6);
assign Wmr7x6 = (~(Lsiov6 & Gtiov6));
assign Lsiov6 = (Dnr7x6 & Osgov6);
assign Dnr7x6 = (Knr7x6 & Cjjov6);
assign Pmr7x6 = (Rnr7x6 & Ynr7x6);
assign Ynr7x6 = (~(Mpiov6 & Ekjov6));
assign Mpiov6 = (Tojov6 & Apjov6);
assign Tojov6 = (Osgov6 & For7x6);
assign Osgov6 = (Mor7x6 & Tor7x6);
assign Rnr7x6 = (~(Rviov6 & Apr7x6));
assign Apr7x6 = (~(Hpr7x6 & Opr7x6));
assign Opr7x6 = (~(K2jov6 | C5jov6));
assign C5jov6 = (Vpr7x6 & Itjov6);
assign Vpr7x6 = (Ptjov6 & Cqr7x6);
assign K2jov6 = (Jqr7x6 & Itjov6);
assign Jqr7x6 = (Qqr7x6 & Kujov6);
assign Hpr7x6 = (Xqr7x6 & Zrjov6);
assign Zrjov6 = (~(Cyiov6 & Err7x6));
assign Cyiov6 = (Lrr7x6 & Srr7x6);
assign Xqr7x6 = (~(E6jov6 & S6jov6));
assign E6jov6 = (Zrr7x6 & Lrr7x6);
assign Bj2nv6 = (~(Vrinv6 & Gsr7x6));
assign Gsr7x6 = (~(Nsr7x6 & Usr7x6));
assign Usr7x6 = (!K73et6);
assign R9r7x6 = (Ub2nv6 & Btr7x6);
assign Btr7x6 = (~(Doadt6 & Itr7x6));
assign Itr7x6 = (~(Ptr7x6 & Wtr7x6));
assign Wtr7x6 = (~(Dur7x6 | Cwlnv6));
assign Ptr7x6 = (Kur7x6 & Rur7x6);
assign Rur7x6 = (~(Yur7x6 & Fvr7x6));
assign Yur7x6 = (Dcnov6 & Nf4ov6);
assign Dcnov6 = (~(Mvr7x6 & Tvr7x6));
assign Tvr7x6 = (~(Vs9ov6 & H0tiw6));
assign H0tiw6 = (!S6cdt6);
assign Mvr7x6 = (~(Awr7x6 & Hwr7x6));
assign Awr7x6 = (Owr7x6 & Vwr7x6);
assign Vwr7x6 = (~(E1wnv6 & S2onv6));
assign Owr7x6 = (~(F02nv6 & Sdh7v6));
assign Ub2nv6 = (Cxr7x6 & V82nv6);
assign V82nv6 = (~(Jxr7x6 & Qxr7x6));
assign Qxr7x6 = (Xxr7x6 & Eyr7x6);
assign Eyr7x6 = (Lyr7x6 & Syr7x6);
assign Syr7x6 = (Zyr7x6 & Gzr7x6);
assign Gzr7x6 = (~(Nzr7x6 | Uzr7x6));
assign Nzr7x6 = (~(B0s7x6 & Yseov6));
assign Zyr7x6 = (I0s7x6 & P0s7x6);
assign Lyr7x6 = (W0s7x6 & D1s7x6);
assign D1s7x6 = (~(K1s7x6 | R1s7x6));
assign W0s7x6 = (~(Y1s7x6 | F2s7x6));
assign Xxr7x6 = (M2s7x6 & T2s7x6);
assign T2s7x6 = (A3s7x6 & H3s7x6);
assign H3s7x6 = (O3s7x6 & V3s7x6);
assign O3s7x6 = (~(C4s7x6 | J4s7x6));
assign A3s7x6 = (~(Q4s7x6 | X4s7x6));
assign M2s7x6 = (E5s7x6 & L5s7x6);
assign L5s7x6 = (~(S5s7x6 | Z5s7x6));
assign E5s7x6 = (~(G6s7x6 | N6s7x6));
assign Jxr7x6 = (U6s7x6 & B7s7x6);
assign B7s7x6 = (I7s7x6 & P7s7x6);
assign P7s7x6 = (W7s7x6 & D8s7x6);
assign D8s7x6 = (~(K8s7x6 | R8s7x6));
assign K8s7x6 = (Y8s7x6 | F9s7x6);
assign W7s7x6 = (~(M9s7x6 | T9s7x6));
assign I7s7x6 = (Aas7x6 & Has7x6);
assign Has7x6 = (~(Oas7x6 | Vas7x6));
assign Aas7x6 = (~(Cbs7x6 | Jbs7x6));
assign U6s7x6 = (Qbs7x6 & Xbs7x6);
assign Xbs7x6 = (Ecs7x6 & Lcs7x6);
assign Lcs7x6 = (~(Scs7x6 | Zcs7x6));
assign Scs7x6 = (Gds7x6 | Nds7x6);
assign Ecs7x6 = (Uds7x6 & Bes7x6);
assign Bes7x6 = (~(Ies7x6 & Pes7x6));
assign Ies7x6 = (~(Wes7x6 & Dfs7x6));
assign Dfs7x6 = (Kfs7x6 & Rfs7x6);
assign Rfs7x6 = (Yfs7x6 & Fgs7x6);
assign Fgs7x6 = (Mgs7x6 & Tgs7x6);
assign Tgs7x6 = (Ahs7x6 & Vueov6);
assign Ahs7x6 = (~(Fhcet6 | Zfcet6));
assign Mgs7x6 = (Hhs7x6 & Ohs7x6);
assign Ohs7x6 = (~(M6j7z6[11] & Ohj7z6[11]));
assign Hhs7x6 = (~(M6j7z6[13] & Ohj7z6[13]));
assign Yfs7x6 = (Vhs7x6 & Cis7x6);
assign Cis7x6 = (Jis7x6 & Qis7x6);
assign Qis7x6 = (~(M6j7z6[15] & Ohj7z6[15]));
assign Jis7x6 = (~(M6j7z6[17] & Ohj7z6[17]));
assign Vhs7x6 = (Xis7x6 & Ejs7x6);
assign Ejs7x6 = (~(M6j7z6[19] & Ohj7z6[19]));
assign Xis7x6 = (~(M6j7z6[1] & Ohj7z6[1]));
assign Kfs7x6 = (Ljs7x6 & Sjs7x6);
assign Sjs7x6 = (Zjs7x6 & Gks7x6);
assign Gks7x6 = (Nks7x6 & Uks7x6);
assign Uks7x6 = (~(M6j7z6[25] & Ohj7z6[25]));
assign Nks7x6 = (Bls7x6 & Ils7x6);
assign Ils7x6 = (~(M6j7z6[21] & Ohj7z6[21]));
assign Bls7x6 = (~(M6j7z6[23] & Ohj7z6[23]));
assign Zjs7x6 = (Pls7x6 & Wls7x6);
assign Wls7x6 = (~(M6j7z6[27] & Ohj7z6[27]));
assign Pls7x6 = (~(M6j7z6[29] & Ohj7z6[29]));
assign Ljs7x6 = (Dms7x6 & Kms7x6);
assign Kms7x6 = (Rms7x6 & Yms7x6);
assign Yms7x6 = (~(M6j7z6[31] & Ohj7z6[31]));
assign Rms7x6 = (~(M6j7z6[33] & Ohj7z6[33]));
assign Dms7x6 = (Fns7x6 & Mns7x6);
assign Mns7x6 = (~(M6j7z6[35] & Ohj7z6[35]));
assign Fns7x6 = (~(M6j7z6[37] & Ohj7z6[37]));
assign Wes7x6 = (Tns7x6 & Aos7x6);
assign Aos7x6 = (Hos7x6 & Oos7x6);
assign Oos7x6 = (Vos7x6 & Cps7x6);
assign Cps7x6 = (Jps7x6 & Qps7x6);
assign Qps7x6 = (~(M6j7z6[41] & Ohj7z6[41]));
assign Jps7x6 = (Xps7x6 & Eqs7x6);
assign Eqs7x6 = (~(M6j7z6[39] & Ohj7z6[39]));
assign Xps7x6 = (~(M6j7z6[3] & Ohj7z6[3]));
assign Vos7x6 = (Lqs7x6 & Sqs7x6);
assign Sqs7x6 = (~(M6j7z6[43] & Ohj7z6[43]));
assign Lqs7x6 = (~(M6j7z6[45] & Ohj7z6[45]));
assign Hos7x6 = (Zqs7x6 & Grs7x6);
assign Grs7x6 = (Nrs7x6 & Urs7x6);
assign Urs7x6 = (~(M6j7z6[47] & Ohj7z6[47]));
assign Nrs7x6 = (~(M6j7z6[49] & Ohj7z6[49]));
assign Zqs7x6 = (Bss7x6 & Iss7x6);
assign Iss7x6 = (~(M6j7z6[51] & Ohj7z6[51]));
assign Bss7x6 = (~(M6j7z6[53] & Ohj7z6[53]));
assign Tns7x6 = (Pss7x6 & Wss7x6);
assign Wss7x6 = (Dts7x6 & Kts7x6);
assign Kts7x6 = (Rts7x6 & Yts7x6);
assign Yts7x6 = (~(M6j7z6[55] & Ohj7z6[55]));
assign Rts7x6 = (~(M6j7z6[57] & Ohj7z6[57]));
assign Dts7x6 = (Fus7x6 & Mus7x6);
assign Mus7x6 = (~(M6j7z6[59] & Ohj7z6[59]));
assign Fus7x6 = (~(M6j7z6[5] & Ohj7z6[5]));
assign Pss7x6 = (Tus7x6 & Avs7x6);
assign Avs7x6 = (Hvs7x6 & Ovs7x6);
assign Ovs7x6 = (~(M6j7z6[61] & Ohj7z6[61]));
assign Hvs7x6 = (~(M6j7z6[63] & Ohj7z6[63]));
assign Tus7x6 = (Vvs7x6 & Cws7x6);
assign Cws7x6 = (~(M6j7z6[7] & Ohj7z6[7]));
assign Vvs7x6 = (~(M6j7z6[9] & Ohj7z6[9]));
assign Uds7x6 = (Yfdov6 | Jws7x6);
assign Yfdov6 = (!Z3j7z6[14]);
assign Qbs7x6 = (Qws7x6 & Xws7x6);
assign Xws7x6 = (Exs7x6 & Lxs7x6);
assign Lxs7x6 = (~(Micet6 & Z3j7z6[12]));
assign Qws7x6 = (Fvjov6 & Sxs7x6);
assign Cxr7x6 = (~(Zxs7x6 & Gys7x6));
assign Gys7x6 = (Nys7x6 & Nxeov6);
assign Nys7x6 = (~(Uys7x6 & Bzs7x6));
assign Bzs7x6 = (~(C92nv6 & Izs7x6));
assign Uys7x6 = (Ev2nv6 & Xg2nv6);
assign Zxs7x6 = (Pzs7x6 & Wzs7x6);
assign Wzs7x6 = (~(Dxgov6 & D0t7x6));
assign D0t7x6 = (~(C92nv6 & Uxeov6));
assign C92nv6 = (K0t7x6 & R0t7x6);
assign R0t7x6 = (~(Y0t7x6 & F1t7x6));
assign F1t7x6 = (~(Mbiov6 & M1t7x6));
assign K0t7x6 = (M1t7x6 | Mbiov6);
assign Mbiov6 = (Mrgov6 & H1m8v6);
assign Mrgov6 = (Hsgov6 ? A2t7x6 : T1t7x6);
assign A2t7x6 = (!H2t7x6);
assign M1t7x6 = (O2t7x6 & V2t7x6);
assign V2t7x6 = (~(C3t7x6 & Cdiov6));
assign Cdiov6 = (Rwl8v6 & C7hov6);
assign C7hov6 = (~(J3t7x6 & Q3t7x6));
assign Q3t7x6 = (~(X3t7x6 & E4t7x6));
assign X3t7x6 = (Rviov6 | L4t7x6);
assign L4t7x6 = (S4t7x6 & Tor7x6);
assign Rviov6 = (Tor7x6 & Z4t7x6);
assign J3t7x6 = (~(Hsgov6 & G5t7x6));
assign C3t7x6 = (N5t7x6 & U5t7x6);
assign U5t7x6 = (~(Qdiov6 & B6t7x6));
assign O2t7x6 = (~(I6t7x6 & Ociov6));
assign Ociov6 = (!Qdiov6);
assign Qdiov6 = (Zyl8v6 & Asgov6);
assign Asgov6 = (Hsgov6 ? W6t7x6 : P6t7x6);
assign Hsgov6 = (!Tor7x6);
assign Tor7x6 = (~(D7t7x6 & K7t7x6));
assign K7t7x6 = (~(R7t7x6 & Y7t7x6));
assign R7t7x6 = (~(F8t7x6 | M8t7x6));
assign D7t7x6 = (~(T8t7x6 & A9t7x6));
assign A9t7x6 = (~(T1t7x6 & H2t7x6));
assign T8t7x6 = (H9t7x6 & O9t7x6);
assign O9t7x6 = (~(V9t7x6 & Cat7x6));
assign Cat7x6 = (H2t7x6 | T1t7x6);
assign T1t7x6 = (!Jat7x6);
assign Jat7x6 = (Mor7x6 ? Xat7x6 : Qat7x6);
assign H2t7x6 = (D9jov6 ? Lbt7x6 : Ebt7x6);
assign V9t7x6 = (Sbt7x6 & Zbt7x6);
assign Zbt7x6 = (~(W6t7x6 & Gct7x6));
assign Gct7x6 = (~(Nct7x6 & G5t7x6));
assign Nct7x6 = (P6t7x6 & Uct7x6);
assign Sbt7x6 = (~(Bdt7x6 & Idt7x6));
assign Idt7x6 = (~(G5t7x6 & Uct7x6));
assign Uct7x6 = (~(E4t7x6 & Pdt7x6));
assign Pdt7x6 = (Z4t7x6 | S4t7x6);
assign E4t7x6 = (~(Wdt7x6 & Z4t7x6));
assign G5t7x6 = (!Det7x6);
assign Det7x6 = (D9jov6 ? Ret7x6 : Ket7x6);
assign D9jov6 = (!Dnjov6);
assign H9t7x6 = (~(Yet7x6 & Fft7x6));
assign Yet7x6 = (Z4t7x6 & Lrr7x6);
assign W6t7x6 = (Dnjov6 ? Tft7x6 : Mft7x6);
assign Dnjov6 = (~(Agt7x6 & F8t7x6));
assign F8t7x6 = (Hgt7x6 | Ogt7x6);
assign Agt7x6 = (~(Vgt7x6 & Cht7x6));
assign Cht7x6 = (Jht7x6 & Qht7x6);
assign Qht7x6 = (~(Xht7x6 & Eit7x6));
assign Eit7x6 = (~(Lit7x6 | Sit7x6));
assign Lit7x6 = (Mft7x6 & Zit7x6);
assign Xht7x6 = (Ket7x6 & Gjt7x6);
assign Gjt7x6 = (!Ret7x6);
assign Ret7x6 = (Zkr7x6 ? Ujt7x6 : Njt7x6);
assign Ket7x6 = (Abjov6 ? Ikt7x6 : Bkt7x6);
assign Jht7x6 = (~(Pkt7x6 & Tft7x6));
assign Pkt7x6 = (~(Mft7x6 | Sit7x6));
assign Sit7x6 = (~(Wkt7x6 | Lbt7x6));
assign Vgt7x6 = (Dlt7x6 & Klt7x6);
assign Klt7x6 = (~(Lbt7x6 & Wkt7x6));
assign Wkt7x6 = (!Ebt7x6);
assign Ebt7x6 = (Skr7x6 ? Ylt7x6 : Rlt7x6);
assign Rlt7x6 = (!Fmt7x6);
assign Lbt7x6 = (Zkr7x6 ? Tmt7x6 : Mmt7x6);
assign Mmt7x6 = (Fajov6 ? Hnt7x6 : Ant7x6);
assign Dlt7x6 = (~(Y7t7x6 & Abjov6));
assign Tft7x6 = (!Zit7x6);
assign Zit7x6 = (Skr7x6 ? Vnt7x6 : Ont7x6);
assign Skr7x6 = (!Abjov6);
assign Abjov6 = (~(Cot7x6 & M8t7x6));
assign M8t7x6 = (~(Jot7x6 & Qot7x6));
assign Jot7x6 = (Xot7x6 & B0s7x6);
assign Cot7x6 = (~(Ept7x6 & Lpt7x6));
assign Lpt7x6 = (~(Ylt7x6 & Spt7x6));
assign Ept7x6 = (~(Zpt7x6 | Y7t7x6));
assign Y7t7x6 = (Gqt7x6 & Exs7x6);
assign Exs7x6 = (Nqt7x6 & Uqt7x6);
assign Uqt7x6 = (~(Brt7x6 & Pes7x6));
assign Gqt7x6 = (Irt7x6 & Prt7x6);
assign Zpt7x6 = (Fmt7x6 & Wrt7x6);
assign Wrt7x6 = (Spt7x6 | Ylt7x6);
assign Ylt7x6 = (Qcjov6 ? Kst7x6 : Dst7x6);
assign Kst7x6 = (!Rst7x6);
assign Spt7x6 = (~(Yst7x6 & Ftt7x6));
assign Ftt7x6 = (Mtt7x6 | Bkt7x6);
assign Bkt7x6 = (Qcjov6 ? Aut7x6 : Ttt7x6);
assign Ttt7x6 = (Xot7x6 ? Lgj7z6[156] : Lgj7z6[159]);
assign Mtt7x6 = (~(Ikt7x6 & Hut7x6));
assign Hut7x6 = (~(Ont7x6 & Out7x6));
assign Ikt7x6 = (!Vut7x6);
assign Vut7x6 = (Vbjov6 ? Jvt7x6 : Cvt7x6);
assign Cvt7x6 = (Irt7x6 ? Xvt7x6 : Qvt7x6);
assign Yst7x6 = (Out7x6 | Ont7x6);
assign Out7x6 = (!Vnt7x6);
assign Fmt7x6 = (Vbjov6 ? Lwt7x6 : Ewt7x6);
assign Vnt7x6 = (Qcjov6 ? Zwt7x6 : Swt7x6);
assign Qcjov6 = (~(Gxt7x6 | Qot7x6));
assign Qot7x6 = (~(Zcs7x6 | Jcjov6));
assign Gxt7x6 = (Nxt7x6 & Uxt7x6);
assign Uxt7x6 = (Byt7x6 & Iyt7x6);
assign Iyt7x6 = (~(Pyt7x6 & Wyt7x6));
assign Wyt7x6 = (Dzt7x6 & Kzt7x6);
assign Dzt7x6 = (Zwt7x6 | Rzt7x6);
assign Pyt7x6 = (~(Yzt7x6 | Aut7x6));
assign Aut7x6 = (Jcjov6 ? Lgj7z6[165] : Lgj7z6[162]);
assign Yzt7x6 = (Ccjov6 ? M0u7x6 : F0u7x6);
assign Byt7x6 = (~(T0u7x6 & Rzt7x6));
assign T0u7x6 = (Zwt7x6 & Kzt7x6);
assign Kzt7x6 = (~(Rst7x6 & Dst7x6));
assign Nxt7x6 = (A1u7x6 & H1u7x6);
assign H1u7x6 = (Dst7x6 | Rst7x6);
assign Rst7x6 = (Jcjov6 ? Lgj7z6[167] : Lgj7z6[164]);
assign Dst7x6 = (Ccjov6 ? V1u7x6 : O1u7x6);
assign A1u7x6 = (~(Xot7x6 & B0s7x6));
assign Zwt7x6 = (Jcjov6 ? J2u7x6 : C2u7x6);
assign Jcjov6 = (Q2u7x6 & X2u7x6);
assign X2u7x6 = (E3u7x6 & Pes7x6);
assign E3u7x6 = (~(Zcs7x6 & L3u7x6));
assign Zcs7x6 = (S3u7x6 & M6j7z6[54]);
assign S3u7x6 = (Ohj7z6[54] & Pes7x6);
assign Q2u7x6 = (M6j7z6[55] & Ohj7z6[55]);
assign Swt7x6 = (!Rzt7x6);
assign Rzt7x6 = (Xot7x6 ? Lgj7z6[157] : Lgj7z6[160]);
assign Xot7x6 = (!Ccjov6);
assign Ccjov6 = (Z3u7x6 & G4u7x6);
assign G4u7x6 = (N4u7x6 & Pes7x6);
assign N4u7x6 = (B0s7x6 | U4u7x6);
assign B0s7x6 = (~(B5u7x6 & M6j7z6[52]));
assign B5u7x6 = (Ohj7z6[52] & Pes7x6);
assign Z3u7x6 = (M6j7z6[53] & Ohj7z6[53]);
assign Ont7x6 = (Vbjov6 ? P5u7x6 : I5u7x6);
assign Vbjov6 = (W5u7x6 & D6u7x6);
assign D6u7x6 = (~(K6u7x6 & R6u7x6));
assign R6u7x6 = (Y6u7x6 & F7u7x6);
assign F7u7x6 = (~(M7u7x6 & T7u7x6));
assign T7u7x6 = (A8u7x6 & H8u7x6);
assign A8u7x6 = (O8u7x6 | P5u7x6);
assign M7u7x6 = (V8u7x6 & Jvt7x6);
assign Jvt7x6 = (Prt7x6 ? J9u7x6 : C9u7x6);
assign V8u7x6 = (Irt7x6 ? Lgj7z6[144] : Lgj7z6[147]);
assign Y6u7x6 = (~(Q9u7x6 & P5u7x6));
assign Q9u7x6 = (O8u7x6 & H8u7x6);
assign H8u7x6 = (X9u7x6 | Ewt7x6);
assign O8u7x6 = (!I5u7x6);
assign K6u7x6 = (Eau7x6 & Lau7x6);
assign Lau7x6 = (Brt7x6 | Hbjov6);
assign Eau7x6 = (~(Ewt7x6 & X9u7x6));
assign X9u7x6 = (!Lwt7x6);
assign Lwt7x6 = (Objov6 ? Lgj7z6[155] : Lgj7z6[152]);
assign Objov6 = (!Prt7x6);
assign Ewt7x6 = (Irt7x6 ? Lgj7z6[146] : Lgj7z6[149]);
assign W5u7x6 = (~(Nqt7x6 & Prt7x6));
assign Nqt7x6 = (!Sau7x6);
assign P5u7x6 = (Prt7x6 ? Gbu7x6 : Zau7x6);
assign Prt7x6 = (~(Nbu7x6 & Ubu7x6));
assign Ubu7x6 = (Bcu7x6 & Pes7x6);
assign Bcu7x6 = (~(Sau7x6 & Icu7x6));
assign Sau7x6 = (Pcu7x6 & M6j7z6[50]);
assign Pcu7x6 = (Ohj7z6[50] & Pes7x6);
assign Nbu7x6 = (M6j7z6[51] & Ohj7z6[51]);
assign I5u7x6 = (Hbjov6 ? Ddu7x6 : Wcu7x6);
assign Hbjov6 = (!Irt7x6);
assign Irt7x6 = (~(Kdu7x6 & Rdu7x6));
assign Rdu7x6 = (Ydu7x6 & Pes7x6);
assign Ydu7x6 = (~(Feu7x6 & Brt7x6));
assign Brt7x6 = (M6j7z6[48] & Ohj7z6[48]);
assign Kdu7x6 = (M6j7z6[49] & Ohj7z6[49]);
assign Mft7x6 = (Zkr7x6 ? Teu7x6 : Meu7x6);
assign Zkr7x6 = (!Y9jov6);
assign Y9jov6 = (~(Afu7x6 & Ogt7x6));
assign Ogt7x6 = (~(Hfu7x6 & Ofu7x6));
assign Hfu7x6 = (~(Zdjov6 | R1s7x6));
assign Afu7x6 = (~(Vfu7x6 & Cgu7x6));
assign Cgu7x6 = (~(Tmt7x6 & Jgu7x6));
assign Jgu7x6 = (~(Qgu7x6 & Xgu7x6));
assign Tmt7x6 = (!Ehu7x6);
assign Vfu7x6 = (Lhu7x6 & Hgt7x6);
assign Hgt7x6 = (~(Shu7x6 & Zhu7x6));
assign Shu7x6 = (Giu7x6 & P0s7x6);
assign Lhu7x6 = (~(Niu7x6 & Uiu7x6));
assign Uiu7x6 = (~(Bju7x6 & Ehu7x6));
assign Ehu7x6 = (Nejov6 ? Pju7x6 : Iju7x6);
assign Bju7x6 = (Xgu7x6 & Qgu7x6);
assign Qgu7x6 = (~(Wju7x6 & Meu7x6));
assign Wju7x6 = (!Teu7x6);
assign Xgu7x6 = (~(Dku7x6 & Kku7x6));
assign Kku7x6 = (!Ujt7x6);
assign Ujt7x6 = (Nejov6 ? Yku7x6 : Rku7x6);
assign Yku7x6 = (Flu7x6 ? Lgj7z6[186] : Lgj7z6[189]);
assign Dku7x6 = (Njt7x6 & Mlu7x6);
assign Mlu7x6 = (~(Tlu7x6 & Teu7x6));
assign Tlu7x6 = (!Meu7x6);
assign Njt7x6 = (!Amu7x6);
assign Amu7x6 = (Pmjov6 ? Omu7x6 : Hmu7x6);
assign Hmu7x6 = (Giu7x6 ? Cnu7x6 : Vmu7x6);
assign Niu7x6 = (Fajov6 ? Qnu7x6 : Jnu7x6);
assign Fajov6 = (!Pmjov6);
assign Teu7x6 = (Nejov6 ? Eou7x6 : Xnu7x6);
assign Nejov6 = (~(Lou7x6 | Ofu7x6));
assign Ofu7x6 = (I0s7x6 & Flu7x6);
assign Lou7x6 = (Sou7x6 & Zou7x6);
assign Zou7x6 = (Zdjov6 | R1s7x6);
assign Sou7x6 = (Gpu7x6 & Npu7x6);
assign Npu7x6 = (~(Upu7x6 & Bqu7x6));
assign Bqu7x6 = (Iqu7x6 | Iju7x6);
assign Upu7x6 = (~(Pqu7x6 & Wqu7x6));
assign Wqu7x6 = (~(Dru7x6 & Kru7x6));
assign Kru7x6 = (Flu7x6 ? Yru7x6 : Rru7x6);
assign Dru7x6 = (Rku7x6 & Fsu7x6);
assign Fsu7x6 = (Xnu7x6 | Msu7x6);
assign Rku7x6 = (Zdjov6 ? Lgj7z6[183] : Lgj7z6[180]);
assign Pqu7x6 = (~(Msu7x6 & Xnu7x6));
assign Msu7x6 = (!Eou7x6);
assign Gpu7x6 = (~(Iju7x6 & Iqu7x6));
assign Iqu7x6 = (!Pju7x6);
assign Pju7x6 = (Gejov6 ? Lgj7z6[191] : Lgj7z6[188]);
assign Iju7x6 = (Zdjov6 ? Lgj7z6[185] : Lgj7z6[182]);
assign Eou7x6 = (Gejov6 ? Lgj7z6[190] : Lgj7z6[187]);
assign Gejov6 = (!Flu7x6);
assign Flu7x6 = (~(Tsu7x6 & Atu7x6));
assign Atu7x6 = (Htu7x6 & Pes7x6);
assign Htu7x6 = (~(Otu7x6 & Vtu7x6));
assign Otu7x6 = (!I0s7x6);
assign I0s7x6 = (~(Cuu7x6 & M6j7z6[62]));
assign Cuu7x6 = (Ohj7z6[62] & Pes7x6);
assign Tsu7x6 = (M6j7z6[63] & Ohj7z6[63]);
assign Xnu7x6 = (Zdjov6 ? Lgj7z6[184] : Lgj7z6[181]);
assign Zdjov6 = (Juu7x6 & Quu7x6);
assign Quu7x6 = (Xuu7x6 & Pes7x6);
assign Xuu7x6 = (~(R1s7x6 & Evu7x6));
assign R1s7x6 = (Lvu7x6 & M6j7z6[60]);
assign Lvu7x6 = (Ohj7z6[60] & Pes7x6);
assign Juu7x6 = (M6j7z6[61] & Ohj7z6[61]);
assign Meu7x6 = (Pmjov6 ? Zvu7x6 : Svu7x6);
assign Pmjov6 = (~(Gwu7x6 | Zhu7x6));
assign Zhu7x6 = (~(Uzr7x6 | Nwu7x6));
assign Gwu7x6 = (Uwu7x6 & Bxu7x6);
assign Bxu7x6 = (~(Giu7x6 & P0s7x6));
assign Uwu7x6 = (Ixu7x6 & Pxu7x6);
assign Pxu7x6 = (~(Wxu7x6 & Dyu7x6));
assign Dyu7x6 = (~(Jnu7x6 & Hnt7x6));
assign Jnu7x6 = (!Ant7x6);
assign Wxu7x6 = (~(Kyu7x6 & Ryu7x6));
assign Ryu7x6 = (~(Yyu7x6 & Fzu7x6));
assign Fzu7x6 = (Giu7x6 ? Lgj7z6[168] : Lgj7z6[171]);
assign Yyu7x6 = (Omu7x6 & Mzu7x6);
assign Mzu7x6 = (Svu7x6 | Tzu7x6);
assign Omu7x6 = (Nwu7x6 ? H0v7x6 : A0v7x6);
assign Kyu7x6 = (~(Tzu7x6 & Svu7x6));
assign Tzu7x6 = (!Zvu7x6);
assign Ixu7x6 = (~(Qnu7x6 & Ant7x6));
assign Ant7x6 = (Bfjov6 ? V0v7x6 : O0v7x6);
assign Bfjov6 = (!Nwu7x6);
assign Qnu7x6 = (!Hnt7x6);
assign Hnt7x6 = (R9jov6 ? J1v7x6 : C1v7x6);
assign Zvu7x6 = (Nwu7x6 ? Lgj7z6[178] : Lgj7z6[175]);
assign Nwu7x6 = (Q1v7x6 & X1v7x6);
assign X1v7x6 = (E2v7x6 & Pes7x6);
assign E2v7x6 = (~(Uzr7x6 & L2v7x6));
assign Uzr7x6 = (S2v7x6 & M6j7z6[58]);
assign S2v7x6 = (Ohj7z6[58] & Pes7x6);
assign Q1v7x6 = (M6j7z6[59] & Ohj7z6[59]);
assign Svu7x6 = (Giu7x6 ? Lgj7z6[169] : Lgj7z6[172]);
assign Giu7x6 = (!R9jov6);
assign R9jov6 = (Z2v7x6 & G3v7x6);
assign G3v7x6 = (N3v7x6 & Pes7x6);
assign N3v7x6 = (P0s7x6 | U3v7x6);
assign P0s7x6 = (~(B4v7x6 & M6j7z6[56]));
assign B4v7x6 = (Ohj7z6[56] & Pes7x6);
assign Z2v7x6 = (M6j7z6[57] & Ohj7z6[57]);
assign P6t7x6 = (!Bdt7x6);
assign Bdt7x6 = (Mor7x6 ? P4v7x6 : I4v7x6);
assign Mor7x6 = (!Z4t7x6);
assign Z4t7x6 = (~(W4v7x6 & D5v7x6));
assign D5v7x6 = (~(K5v7x6 & R5v7x6));
assign R5v7x6 = (Y5v7x6 & F6v7x6);
assign F6v7x6 = (~(M6v7x6 & T6v7x6));
assign M6v7x6 = (P4v7x6 & A7v7x6);
assign Y5v7x6 = (~(Fft7x6 & Lrr7x6));
assign K5v7x6 = (H7v7x6 & O7v7x6);
assign O7v7x6 = (~(V7v7x6 & C8v7x6));
assign C8v7x6 = (J8v7x6 & A7v7x6);
assign A7v7x6 = (~(Qat7x6 & Q8v7x6));
assign J8v7x6 = (P4v7x6 | T6v7x6);
assign V7v7x6 = (Wdt7x6 & S4t7x6);
assign S4t7x6 = (For7x6 ? E9v7x6 : X8v7x6);
assign Wdt7x6 = (Lrr7x6 ? S9v7x6 : L9v7x6);
assign H7v7x6 = (Q8v7x6 | Qat7x6);
assign Qat7x6 = (Itjov6 ? Gav7x6 : Z9v7x6);
assign Q8v7x6 = (!Xat7x6);
assign Xat7x6 = (For7x6 ? Uav7x6 : Nav7x6);
assign Uav7x6 = (Bbv7x6 & Ibv7x6);
assign W4v7x6 = (Pbv7x6 | Wbv7x6);
assign P4v7x6 = (For7x6 ? Kcv7x6 : Dcv7x6);
assign For7x6 = (!Cjjov6);
assign Cjjov6 = (~(Wbv7x6 & Rcv7x6));
assign Rcv7x6 = (~(Ycv7x6 & Fdv7x6));
assign Fdv7x6 = (~(Mdv7x6 & Bbv7x6));
assign Bbv7x6 = (Apjov6 | Tdv7x6);
assign Mdv7x6 = (Aev7x6 & Ibv7x6);
assign Ibv7x6 = (~(Hev7x6 & Apjov6));
assign Aev7x6 = (~(Oev7x6 & Nav7x6));
assign Nav7x6 = (!Vev7x6);
assign Oev7x6 = (Cfv7x6 & Jfv7x6);
assign Jfv7x6 = (Qfv7x6 | Xfv7x6);
assign Ycv7x6 = (Egv7x6 & Pbv7x6);
assign Pbv7x6 = (~(Lgv7x6 & Sgv7x6));
assign Lgv7x6 = (~(Zgv7x6 | Ghv7x6));
assign Egv7x6 = (~(Nhv7x6 & Vev7x6));
assign Vev7x6 = (Knr7x6 ? Biv7x6 : Uhv7x6);
assign Nhv7x6 = (~(Iiv7x6 | Xfv7x6));
assign Xfv7x6 = (Piv7x6 & Dcv7x6);
assign Piv7x6 = (!Kcv7x6);
assign Iiv7x6 = (Qfv7x6 & Cfv7x6);
assign Cfv7x6 = (~(Wiv7x6 & Kcv7x6));
assign Qfv7x6 = (~(E9v7x6 & Djv7x6));
assign Djv7x6 = (!X8v7x6);
assign X8v7x6 = (Knr7x6 ? Rjv7x6 : Kjv7x6);
assign E9v7x6 = (Apjov6 ? Fkv7x6 : Yjv7x6);
assign Wbv7x6 = (~(Mkv7x6 & Tkv7x6));
assign Mkv7x6 = (~(Alv7x6 | Hlv7x6));
assign Kcv7x6 = (Apjov6 ? Vlv7x6 : Olv7x6);
assign Apjov6 = (~(Alv7x6 & Cmv7x6));
assign Cmv7x6 = (~(Jmv7x6 & Qmv7x6));
assign Qmv7x6 = (Xmv7x6 & Env7x6);
assign Env7x6 = (~(Lnv7x6 & Snv7x6));
assign Snv7x6 = (Znv7x6 & Gov7x6);
assign Znv7x6 = (Olv7x6 | Nov7x6);
assign Lnv7x6 = (Uov7x6 & Yjv7x6);
assign Yjv7x6 = (Hpjov6 ? Ipv7x6 : Bpv7x6);
assign Uov7x6 = (!Fkv7x6);
assign Fkv7x6 = (Hqiov6 ? Wpv7x6 : Ppv7x6);
assign Xmv7x6 = (~(Dqv7x6 & Nov7x6));
assign Nov7x6 = (!Vlv7x6);
assign Dqv7x6 = (Olv7x6 & Gov7x6);
assign Gov7x6 = (Hev7x6 | Tdv7x6);
assign Jmv7x6 = (Kqv7x6 & Rqv7x6);
assign Rqv7x6 = (~(Tdv7x6 & Hev7x6));
assign Hev7x6 = (Hqiov6 ? Frv7x6 : Yqv7x6);
assign Yqv7x6 = (!Mrv7x6);
assign Tdv7x6 = (Nlr7x6 ? Asv7x6 : Trv7x6);
assign Nlr7x6 = (!Hpjov6);
assign Asv7x6 = (!Hsv7x6);
assign Kqv7x6 = (Hlv7x6 | Ekjov6);
assign Alv7x6 = (Osv7x6 | Vsv7x6);
assign Vlv7x6 = (Ekjov6 ? Jtv7x6 : Ctv7x6);
assign Ekjov6 = (!Hqiov6);
assign Hqiov6 = (Qtv7x6 | Tkv7x6);
assign Tkv7x6 = (~(Xtv7x6 | Euv7x6));
assign Qtv7x6 = (Luv7x6 & Suv7x6);
assign Suv7x6 = (~(Mrv7x6 & Zuv7x6));
assign Luv7x6 = (Gvv7x6 & Hlv7x6);
assign Hlv7x6 = (~(Nvv7x6 & Uvv7x6));
assign Uvv7x6 = (~(Vqiov6 | Jbs7x6));
assign Nvv7x6 = (~(Oqiov6 | Cbs7x6));
assign Gvv7x6 = (~(Frv7x6 & Bwv7x6));
assign Bwv7x6 = (Zuv7x6 | Mrv7x6);
assign Mrv7x6 = (Wwv7x6 ? Pwv7x6 : Iwv7x6);
assign Zuv7x6 = (~(Dxv7x6 & Kxv7x6));
assign Kxv7x6 = (~(Rxv7x6 & Ppv7x6));
assign Ppv7x6 = (Wwv7x6 ? Fyv7x6 : Yxv7x6);
assign Fyv7x6 = (Tyv7x6 ? Q88iw6 : Myv7x6);
assign Rxv7x6 = (~(Wpv7x6 | Azv7x6));
assign Azv7x6 = (Ctv7x6 & Hzv7x6);
assign Wpv7x6 = (C0w7x6 ? Vzv7x6 : Ozv7x6);
assign Vzv7x6 = (Oqiov6 ? J0w7x6 : Ua8iw6);
assign Dxv7x6 = (Hzv7x6 | Ctv7x6);
assign Frv7x6 = (C0w7x6 ? X0w7x6 : Q0w7x6);
assign Jtv7x6 = (!Hzv7x6);
assign Hzv7x6 = (Wwv7x6 ? L1w7x6 : E1w7x6);
assign Wwv7x6 = (!Xriov6);
assign Xriov6 = (Xtv7x6 & S1w7x6);
assign S1w7x6 = (~(Z1w7x6 & G2w7x6));
assign G2w7x6 = (N2w7x6 & Euv7x6);
assign Euv7x6 = (Jriov6 | Nds7x6);
assign Nds7x6 = (U2w7x6 & M6j7z6[36]);
assign U2w7x6 = (Ohj7z6[36] & Pes7x6);
assign N2w7x6 = (~(B3w7x6 & L1w7x6));
assign B3w7x6 = (I3w7x6 & P3w7x6);
assign Z1w7x6 = (W3w7x6 & D4w7x6);
assign D4w7x6 = (~(K4w7x6 & R4w7x6));
assign R4w7x6 = (Y4w7x6 & P3w7x6);
assign P3w7x6 = (Iwv7x6 | F5w7x6);
assign Y4w7x6 = (I3w7x6 | L1w7x6);
assign I3w7x6 = (!E1w7x6);
assign K4w7x6 = (M5w7x6 & Yxv7x6);
assign Yxv7x6 = (Qriov6 ? A6w7x6 : T5w7x6);
assign M5w7x6 = (Tyv7x6 ? Lgj7z6[108] : Lgj7z6[111]);
assign W3w7x6 = (~(F5w7x6 & Iwv7x6));
assign Iwv7x6 = (Qriov6 ? O6w7x6 : H6w7x6);
assign F5w7x6 = (!Pwv7x6);
assign Pwv7x6 = (Jriov6 ? V6w7x6 : Yd7iw6);
assign Jriov6 = (!Tyv7x6);
assign Xtv7x6 = (Qriov6 | Oas7x6);
assign L1w7x6 = (Tyv7x6 ? Lgj7z6[109] : Lgj7z6[112]);
assign Tyv7x6 = (~(C7w7x6 & J7w7x6));
assign J7w7x6 = (Q7w7x6 & Pes7x6);
assign Q7w7x6 = (~(X7w7x6 & E8w7x6));
assign X7w7x6 = (M6j7z6[36] & Ohj7z6[36]);
assign C7w7x6 = (M6j7z6[37] & Ohj7z6[37]);
assign E1w7x6 = (Qriov6 ? Lgj7z6[118] : Lgj7z6[115]);
assign Qriov6 = (L8w7x6 & S8w7x6);
assign S8w7x6 = (Z8w7x6 & Pes7x6);
assign Z8w7x6 = (~(Oas7x6 & G9w7x6));
assign Oas7x6 = (N9w7x6 & M6j7z6[38]);
assign N9w7x6 = (Ohj7z6[38] & Pes7x6);
assign L8w7x6 = (M6j7z6[39] & Ohj7z6[39]);
assign Ctv7x6 = (C0w7x6 ? Baw7x6 : U9w7x6);
assign C0w7x6 = (!Criov6);
assign Criov6 = (Iaw7x6 & Paw7x6);
assign Paw7x6 = (~(Waw7x6 & Dbw7x6));
assign Dbw7x6 = (Oqiov6 | Cbs7x6);
assign Waw7x6 = (Kbw7x6 & Rbw7x6);
assign Rbw7x6 = (~(Ybw7x6 & Fcw7x6));
assign Fcw7x6 = (Mcw7x6 | X0w7x6);
assign Ybw7x6 = (~(Tcw7x6 & Adw7x6));
assign Adw7x6 = (~(Hdw7x6 & Odw7x6));
assign Odw7x6 = (Oqiov6 ? Lgj7z6[99] : Lgj7z6[96]);
assign Hdw7x6 = (Ozv7x6 & Vdw7x6);
assign Vdw7x6 = (U9w7x6 | Cew7x6);
assign Ozv7x6 = (Xew7x6 ? Qew7x6 : Jew7x6);
assign Tcw7x6 = (~(Cew7x6 & U9w7x6));
assign Cew7x6 = (!Baw7x6);
assign Kbw7x6 = (~(X0w7x6 & Mcw7x6));
assign Mcw7x6 = (!Q0w7x6);
assign Q0w7x6 = (Vqiov6 ? Lgj7z6[107] : Lgj7z6[104]);
assign X0w7x6 = (Oqiov6 ? Lgj7z6[101] : Lgj7z6[98]);
assign Iaw7x6 = (Jbs7x6 | Vqiov6);
assign Baw7x6 = (Oqiov6 ? Efw7x6 : Ju7iw6);
assign Oqiov6 = (Lfw7x6 & Sfw7x6);
assign Sfw7x6 = (Zfw7x6 & Pes7x6);
assign Zfw7x6 = (~(Cbs7x6 & Ggw7x6));
assign Cbs7x6 = (Ngw7x6 & M6j7z6[32]);
assign Ngw7x6 = (Ohj7z6[32] & Pes7x6);
assign Lfw7x6 = (M6j7z6[33] & Ohj7z6[33]);
assign U9w7x6 = (Xew7x6 ? Bhw7x6 : Ugw7x6);
assign Xew7x6 = (!Vqiov6);
assign Vqiov6 = (Ihw7x6 & Phw7x6);
assign Phw7x6 = (Whw7x6 & Pes7x6);
assign Whw7x6 = (~(Jbs7x6 & Diw7x6));
assign Jbs7x6 = (Kiw7x6 & M6j7z6[34]);
assign Kiw7x6 = (Ohj7z6[34] & Pes7x6);
assign Ihw7x6 = (M6j7z6[35] & Ohj7z6[35]);
assign Olv7x6 = (Hpjov6 ? Yiw7x6 : Riw7x6);
assign Hpjov6 = (Fjw7x6 & Osv7x6);
assign Osv7x6 = (~(Mjw7x6 & Tjw7x6));
assign Mjw7x6 = (~(Iniov6 | Vas7x6));
assign Fjw7x6 = (~(Akw7x6 & Hkw7x6));
assign Hkw7x6 = (~(Trv7x6 & Hsv7x6));
assign Akw7x6 = (Okw7x6 & Vsv7x6);
assign Vsv7x6 = (~(Vkw7x6 & Clw7x6));
assign Vkw7x6 = (~(Ckiov6 | T9s7x6));
assign Okw7x6 = (~(Jlw7x6 & Qlw7x6));
assign Qlw7x6 = (Hsv7x6 | Trv7x6);
assign Trv7x6 = (Wniov6 ? Emw7x6 : Xlw7x6);
assign Hsv7x6 = (Zmw7x6 ? Smw7x6 : Lmw7x6);
assign Jlw7x6 = (~(Gnw7x6 & Nnw7x6));
assign Nnw7x6 = (~(Unw7x6 & Yiw7x6));
assign Gnw7x6 = (~(Bow7x6 & Ipv7x6));
assign Ipv7x6 = (Wniov6 ? Pow7x6 : Iow7x6);
assign Bow7x6 = (~(Bpv7x6 | Wow7x6));
assign Wow7x6 = (~(Yiw7x6 | Unw7x6));
assign Unw7x6 = (!Riw7x6);
assign Bpv7x6 = (Zmw7x6 ? Kpw7x6 : Dpw7x6);
assign Kpw7x6 = (Ckiov6 ? Rpw7x6 : O78iw6);
assign Yiw7x6 = (Wniov6 ? Fqw7x6 : Ypw7x6);
assign Wniov6 = (~(Tjw7x6 | Mqw7x6));
assign Mqw7x6 = (Tqw7x6 & Arw7x6);
assign Arw7x6 = (Iniov6 | Vas7x6);
assign Tqw7x6 = (Hrw7x6 & Orw7x6);
assign Orw7x6 = (~(Vrw7x6 & Csw7x6));
assign Csw7x6 = (Emw7x6 | Jsw7x6);
assign Vrw7x6 = (~(Qsw7x6 & Xsw7x6));
assign Xsw7x6 = (Etw7x6 | Iow7x6);
assign Iow7x6 = (Iniov6 ? Ltw7x6 : M68iw6);
assign Etw7x6 = (~(Pow7x6 & Stw7x6));
assign Stw7x6 = (Ztw7x6 | Fqw7x6);
assign Pow7x6 = (Pniov6 ? Nuw7x6 : Guw7x6);
assign Qsw7x6 = (~(Fqw7x6 & Ztw7x6));
assign Ztw7x6 = (!Ypw7x6);
assign Hrw7x6 = (~(Jsw7x6 & Emw7x6));
assign Emw7x6 = (Ivw7x6 ? Bvw7x6 : Uuw7x6);
assign Jsw7x6 = (!Xlw7x6);
assign Xlw7x6 = (Iniov6 ? Pvw7x6 : Ub7iw6);
assign Tjw7x6 = (~(M9s7x6 | Pniov6));
assign Fqw7x6 = (Ivw7x6 ? Dww7x6 : Wvw7x6);
assign Ivw7x6 = (!Pniov6);
assign Pniov6 = (Kww7x6 & Rww7x6);
assign Rww7x6 = (Yww7x6 & Pes7x6);
assign Yww7x6 = (~(M9s7x6 & Fxw7x6));
assign M9s7x6 = (Mxw7x6 & M6j7z6[46]);
assign Mxw7x6 = (Ohj7z6[46] & Pes7x6);
assign Kww7x6 = (M6j7z6[47] & Ohj7z6[47]);
assign Ypw7x6 = (Iniov6 ? Txw7x6 : Yr7iw6);
assign Iniov6 = (Ayw7x6 & Hyw7x6);
assign Hyw7x6 = (Oyw7x6 & Pes7x6);
assign Oyw7x6 = (~(Vas7x6 & Vyw7x6));
assign Vas7x6 = (Czw7x6 & M6j7z6[44]);
assign Czw7x6 = (Ohj7z6[44] & Pes7x6);
assign Ayw7x6 = (M6j7z6[45] & Ohj7z6[45]);
assign Riw7x6 = (Zmw7x6 ? Qzw7x6 : Jzw7x6);
assign Zmw7x6 = (!Qkiov6);
assign Qkiov6 = (~(Xzw7x6 | Clw7x6));
assign Clw7x6 = (~(R8s7x6 | Jkiov6));
assign Xzw7x6 = (E0x7x6 & L0x7x6);
assign L0x7x6 = (Ckiov6 | T9s7x6);
assign E0x7x6 = (S0x7x6 & Z0x7x6);
assign Z0x7x6 = (~(G1x7x6 & N1x7x6));
assign N1x7x6 = (U1x7x6 | Smw7x6);
assign G1x7x6 = (~(B2x7x6 & I2x7x6));
assign I2x7x6 = (~(P2x7x6 & W2x7x6));
assign W2x7x6 = (Ckiov6 ? Lgj7z6[123] : Lgj7z6[120]);
assign P2x7x6 = (Dpw7x6 & D3x7x6);
assign D3x7x6 = (K3x7x6 | Jzw7x6);
assign Dpw7x6 = (F4x7x6 ? Y3x7x6 : R3x7x6);
assign B2x7x6 = (~(Jzw7x6 & K3x7x6));
assign K3x7x6 = (!Qzw7x6);
assign S0x7x6 = (~(Smw7x6 & U1x7x6));
assign U1x7x6 = (!Lmw7x6);
assign Lmw7x6 = (Jkiov6 ? Lgj7z6[131] : Lgj7z6[128]);
assign Jkiov6 = (!F4x7x6);
assign Smw7x6 = (Ckiov6 ? Lgj7z6[125] : Lgj7z6[122]);
assign Qzw7x6 = (Ckiov6 ? M4x7x6 : Ts7iw6);
assign Ckiov6 = (T4x7x6 & A5x7x6);
assign A5x7x6 = (H5x7x6 & Pes7x6);
assign H5x7x6 = (~(T9s7x6 & O5x7x6));
assign T9s7x6 = (V5x7x6 & M6j7z6[40]);
assign V5x7x6 = (Ohj7z6[40] & Pes7x6);
assign T4x7x6 = (M6j7z6[41] & Ohj7z6[41]);
assign Jzw7x6 = (F4x7x6 ? J6x7x6 : C6x7x6);
assign F4x7x6 = (~(Q6x7x6 & X6x7x6));
assign X6x7x6 = (E7x7x6 & Pes7x6);
assign E7x7x6 = (~(R8s7x6 & L7x7x6));
assign R8s7x6 = (S7x7x6 & M6j7z6[42]);
assign S7x7x6 = (Ohj7z6[42] & Pes7x6);
assign Q6x7x6 = (M6j7z6[43] & Ohj7z6[43]);
assign Dcv7x6 = (!Wiv7x6);
assign Wiv7x6 = (Knr7x6 ? G8x7x6 : Z7x7x6);
assign Knr7x6 = (!Jjjov6);
assign Jjjov6 = (~(N8x7x6 & Ghv7x6));
assign Ghv7x6 = (U8x7x6 | B9x7x6);
assign N8x7x6 = (~(I9x7x6 & P9x7x6));
assign P9x7x6 = (W9x7x6 & Dax7x6);
assign Dax7x6 = (~(Kax7x6 & Rax7x6));
assign Rax7x6 = (Yax7x6 & Fbx7x6);
assign Yax7x6 = (Mbx7x6 | Z7x7x6);
assign Kax7x6 = (Tbx7x6 & Rjv7x6);
assign Rjv7x6 = (Gtiov6 ? Hcx7x6 : Acx7x6);
assign Tbx7x6 = (!Kjv7x6);
assign Kjv7x6 = (Qjjov6 ? Vcx7x6 : Ocx7x6);
assign W9x7x6 = (~(Cdx7x6 & Z7x7x6));
assign Cdx7x6 = (Mbx7x6 & Fbx7x6);
assign Fbx7x6 = (Uhv7x6 | Jdx7x6);
assign Mbx7x6 = (!G8x7x6);
assign I9x7x6 = (Qdx7x6 & Xdx7x6);
assign Xdx7x6 = (~(Jdx7x6 & Uhv7x6));
assign Uhv7x6 = (Qjjov6 ? Lex7x6 : Eex7x6);
assign Eex7x6 = (!Sex7x6);
assign Jdx7x6 = (!Biv7x6);
assign Biv7x6 = (Gtiov6 ? Gfx7x6 : Zex7x6);
assign Qdx7x6 = (~(Sgv7x6 & Qjjov6));
assign G8x7x6 = (Gtiov6 ? Ufx7x6 : Nfx7x6);
assign Gtiov6 = (Bgx7x6 & B9x7x6);
assign B9x7x6 = (~(Igx7x6 & Pgx7x6));
assign Igx7x6 = (~(Ntiov6 | G6s7x6));
assign Bgx7x6 = (~(Wgx7x6 & Dhx7x6));
assign Dhx7x6 = (Gfx7x6 | Khx7x6);
assign Wgx7x6 = (Rhx7x6 & U8x7x6);
assign U8x7x6 = (~(Yhx7x6 & Fix7x6));
assign Yhx7x6 = (~(Iuiov6 | S5s7x6));
assign Rhx7x6 = (~(Mix7x6 & Tix7x6));
assign Tix7x6 = (~(Khx7x6 & Gfx7x6));
assign Gfx7x6 = (Ojx7x6 ? Hjx7x6 : Ajx7x6);
assign Khx7x6 = (!Zex7x6);
assign Zex7x6 = (Jkx7x6 ? Ckx7x6 : Vjx7x6);
assign Mix7x6 = (~(Qkx7x6 & Xkx7x6));
assign Xkx7x6 = (Elx7x6 | Ufx7x6);
assign Qkx7x6 = (~(Llx7x6 & Hcx7x6));
assign Hcx7x6 = (Ojx7x6 ? Zlx7x6 : Slx7x6);
assign Llx7x6 = (~(Acx7x6 | Gmx7x6));
assign Gmx7x6 = (Ufx7x6 & Elx7x6);
assign Acx7x6 = (Jkx7x6 ? Umx7x6 : Nmx7x6);
assign Umx7x6 = (Iuiov6 ? Inx7x6 : Bnx7x6);
assign Ufx7x6 = (Ojx7x6 ? Wnx7x6 : Pnx7x6);
assign Ojx7x6 = (!Buiov6);
assign Buiov6 = (~(Dox7x6 | Pgx7x6));
assign Pgx7x6 = (~(N6s7x6 | Utiov6));
assign Dox7x6 = (Kox7x6 & Rox7x6);
assign Rox7x6 = (Ntiov6 | G6s7x6);
assign Kox7x6 = (Yox7x6 & Fpx7x6);
assign Fpx7x6 = (~(Mpx7x6 & Tpx7x6));
assign Tpx7x6 = (Aqx7x6 | Hjx7x6);
assign Mpx7x6 = (~(Hqx7x6 & Oqx7x6));
assign Oqx7x6 = (Vqx7x6 | Zlx7x6);
assign Zlx7x6 = (Ntiov6 ? Gq6iw6 : Crx7x6);
assign Vqx7x6 = (~(Slx7x6 & Jrx7x6));
assign Jrx7x6 = (Wnx7x6 | Qrx7x6);
assign Slx7x6 = (Utiov6 ? Esx7x6 : Xrx7x6);
assign Hqx7x6 = (~(Qrx7x6 & Wnx7x6));
assign Qrx7x6 = (!Pnx7x6);
assign Yox7x6 = (~(Hjx7x6 & Aqx7x6));
assign Aqx7x6 = (!Ajx7x6);
assign Ajx7x6 = (Utiov6 ? Lgj7z6[95] : Lgj7z6[92]);
assign Hjx7x6 = (Lsx7x6 ? Lgj7z6[86] : Lgj7z6[89]);
assign Wnx7x6 = (Lsx7x6 ? Lgj7z6[85] : Lgj7z6[88]);
assign Lsx7x6 = (!Ntiov6);
assign Ntiov6 = (Ssx7x6 & Zsx7x6);
assign Zsx7x6 = (Gtx7x6 & Pes7x6);
assign Gtx7x6 = (~(G6s7x6 & Ntx7x6));
assign G6s7x6 = (Utx7x6 & M6j7z6[28]);
assign Utx7x6 = (Ohj7z6[28] & Pes7x6);
assign Ssx7x6 = (M6j7z6[29] & Ohj7z6[29]);
assign Pnx7x6 = (Utiov6 ? Lgj7z6[94] : Lgj7z6[91]);
assign Utiov6 = (Bux7x6 & Iux7x6);
assign Iux7x6 = (Pux7x6 & Pes7x6);
assign Pux7x6 = (~(N6s7x6 & Wux7x6));
assign N6s7x6 = (Dvx7x6 & M6j7z6[30]);
assign Dvx7x6 = (Ohj7z6[30] & Pes7x6);
assign Bux7x6 = (M6j7z6[31] & Ohj7z6[31]);
assign Nfx7x6 = (!Elx7x6);
assign Elx7x6 = (Jkx7x6 ? Rvx7x6 : Kvx7x6);
assign Jkx7x6 = (!Wuiov6);
assign Wuiov6 = (~(Yvx7x6 | Fix7x6));
assign Fix7x6 = (~(Z5s7x6 | Puiov6));
assign Yvx7x6 = (Fwx7x6 & Mwx7x6);
assign Mwx7x6 = (Iuiov6 | S5s7x6);
assign Fwx7x6 = (Twx7x6 & Axx7x6);
assign Axx7x6 = (~(Hxx7x6 & Oxx7x6));
assign Oxx7x6 = (Vxx7x6 | Ckx7x6);
assign Hxx7x6 = (~(Cyx7x6 & Jyx7x6));
assign Jyx7x6 = (~(Qyx7x6 & Xyx7x6));
assign Xyx7x6 = (Iuiov6 ? Lgj7z6[75] : Lgj7z6[72]);
assign Qyx7x6 = (Nmx7x6 & Ezx7x6);
assign Ezx7x6 = (Lzx7x6 | Kvx7x6);
assign Nmx7x6 = (G0y7x6 ? Zzx7x6 : Szx7x6);
assign Cyx7x6 = (~(Kvx7x6 & Lzx7x6));
assign Lzx7x6 = (!Rvx7x6);
assign Twx7x6 = (~(Ckx7x6 & Vxx7x6));
assign Vxx7x6 = (!Vjx7x6);
assign Vjx7x6 = (Puiov6 ? Lgj7z6[83] : Lgj7z6[80]);
assign Ckx7x6 = (Iuiov6 ? Lgj7z6[77] : Lgj7z6[74]);
assign Rvx7x6 = (Iuiov6 ? U0y7x6 : N0y7x6);
assign Iuiov6 = (B1y7x6 & I1y7x6);
assign I1y7x6 = (P1y7x6 & Pes7x6);
assign P1y7x6 = (~(S5s7x6 & W1y7x6));
assign S5s7x6 = (D2y7x6 & M6j7z6[24]);
assign D2y7x6 = (Ohj7z6[24] & Pes7x6);
assign B1y7x6 = (M6j7z6[25] & Ohj7z6[25]);
assign Kvx7x6 = (G0y7x6 ? R2y7x6 : K2y7x6);
assign G0y7x6 = (!Puiov6);
assign Puiov6 = (Y2y7x6 & F3y7x6);
assign F3y7x6 = (M3y7x6 & Pes7x6);
assign M3y7x6 = (~(Z5s7x6 & T3y7x6));
assign Z5s7x6 = (A4y7x6 & M6j7z6[26]);
assign A4y7x6 = (Ohj7z6[26] & Pes7x6);
assign Y2y7x6 = (M6j7z6[27] & Ohj7z6[27]);
assign Z7x7x6 = (Qjjov6 ? O4y7x6 : H4y7x6);
assign Qjjov6 = (~(V4y7x6 & Zgv7x6));
assign Zgv7x6 = (~(C5y7x6 & J5y7x6));
assign C5y7x6 = (~(Zliov6 | Y8s7x6));
assign V4y7x6 = (~(Q5y7x6 & X5y7x6));
assign X5y7x6 = (~(Sex7x6 & E6y7x6));
assign Q5y7x6 = (~(L6y7x6 | Sgv7x6));
assign Sgv7x6 = (S6y7x6 & Sxs7x6);
assign Sxs7x6 = (Z6y7x6 & G7y7x6);
assign G7y7x6 = (~(N7y7x6 & Pes7x6));
assign S6y7x6 = (U7y7x6 & B8y7x6);
assign L6y7x6 = (Lex7x6 & I8y7x6);
assign I8y7x6 = (E6y7x6 | Sex7x6);
assign Sex7x6 = (Nmiov6 ? W8y7x6 : P8y7x6);
assign E6y7x6 = (~(D9y7x6 & K9y7x6));
assign K9y7x6 = (~(R9y7x6 & Ocx7x6));
assign Ocx7x6 = (Nmiov6 ? Fay7x6 : Y9y7x6);
assign Fay7x6 = (Gmiov6 ? Tay7x6 : May7x6);
assign R9y7x6 = (~(Vcx7x6 | Aby7x6));
assign Aby7x6 = (Hby7x6 & H4y7x6);
assign Vcx7x6 = (Hjiov6 ? Vby7x6 : Oby7x6);
assign Oby7x6 = (U7y7x6 ? Jcy7x6 : Ccy7x6);
assign D9y7x6 = (H4y7x6 | Hby7x6);
assign Lex7x6 = (Hjiov6 ? Xcy7x6 : Qcy7x6);
assign O4y7x6 = (!Hby7x6);
assign Hby7x6 = (Hjiov6 ? Ldy7x6 : Edy7x6);
assign Hjiov6 = (Sdy7x6 & Zdy7x6);
assign Zdy7x6 = (~(Gey7x6 & Ney7x6));
assign Ney7x6 = (Uey7x6 & Bfy7x6);
assign Bfy7x6 = (~(Ify7x6 & Pfy7x6));
assign Pfy7x6 = (Wfy7x6 & Dgy7x6);
assign Wfy7x6 = (Kgy7x6 | Ldy7x6);
assign Ify7x6 = (Rgy7x6 & Vby7x6);
assign Vby7x6 = (B8y7x6 ? Fhy7x6 : Ygy7x6);
assign Rgy7x6 = (U7y7x6 ? Lgj7z6[48] : Lgj7z6[51]);
assign Uey7x6 = (~(Mhy7x6 & Ldy7x6));
assign Mhy7x6 = (Kgy7x6 & Dgy7x6);
assign Dgy7x6 = (Thy7x6 | Qcy7x6);
assign Kgy7x6 = (!Edy7x6);
assign Gey7x6 = (Aiy7x6 & Hiy7x6);
assign Hiy7x6 = (N7y7x6 | Tiiov6);
assign Aiy7x6 = (~(Qcy7x6 & Thy7x6));
assign Thy7x6 = (!Xcy7x6);
assign Xcy7x6 = (Ajiov6 ? Lgj7z6[59] : Lgj7z6[56]);
assign Ajiov6 = (!B8y7x6);
assign Qcy7x6 = (U7y7x6 ? Lgj7z6[50] : Lgj7z6[53]);
assign Sdy7x6 = (~(Z6y7x6 & B8y7x6));
assign Ldy7x6 = (B8y7x6 ? Viy7x6 : Oiy7x6);
assign B8y7x6 = (~(Cjy7x6 & Jjy7x6));
assign Jjy7x6 = (Qjy7x6 & Pes7x6);
assign Qjy7x6 = (Z6y7x6 | Xjy7x6);
assign Z6y7x6 = (~(Eky7x6 & M6j7z6[18]));
assign Eky7x6 = (Ohj7z6[18] & Pes7x6);
assign Cjy7x6 = (M6j7z6[19] & Ohj7z6[19]);
assign Edy7x6 = (Tiiov6 ? Sky7x6 : Lky7x6);
assign Tiiov6 = (!U7y7x6);
assign U7y7x6 = (~(Zky7x6 & Gly7x6));
assign Gly7x6 = (Nly7x6 & Pes7x6);
assign Nly7x6 = (~(Uly7x6 & N7y7x6));
assign N7y7x6 = (M6j7z6[16] & Ohj7z6[16]);
assign Zky7x6 = (M6j7z6[17] & Ohj7z6[17]);
assign H4y7x6 = (Nmiov6 ? Imy7x6 : Bmy7x6);
assign Nmiov6 = (~(Pmy7x6 | J5y7x6));
assign J5y7x6 = (~(F9s7x6 | Gmiov6));
assign Pmy7x6 = (Wmy7x6 & Dny7x6);
assign Dny7x6 = (Zliov6 | Y8s7x6);
assign Wmy7x6 = (Kny7x6 & Rny7x6);
assign Rny7x6 = (~(Yny7x6 & Foy7x6));
assign Foy7x6 = (W8y7x6 | Moy7x6);
assign Yny7x6 = (~(Toy7x6 & Apy7x6));
assign Apy7x6 = (~(Hpy7x6 & Opy7x6));
assign Opy7x6 = (Vpy7x6 ? May7x6 : Tay7x6);
assign Hpy7x6 = (~(Y9y7x6 | Cqy7x6));
assign Cqy7x6 = (~(Bmy7x6 | Jqy7x6));
assign Y9y7x6 = (Zliov6 ? Qqy7x6 : Ae8iw6);
assign Toy7x6 = (~(Jqy7x6 & Bmy7x6));
assign Jqy7x6 = (!Imy7x6);
assign Kny7x6 = (~(Moy7x6 & W8y7x6));
assign W8y7x6 = (Vpy7x6 ? Ery7x6 : Xqy7x6);
assign Vpy7x6 = (!Gmiov6);
assign Moy7x6 = (!P8y7x6);
assign P8y7x6 = (Zliov6 ? Lry7x6 : Sh7iw6);
assign Imy7x6 = (Gmiov6 ? Lgj7z6[70] : Lgj7z6[67]);
assign Gmiov6 = (Sry7x6 & Zry7x6);
assign Zry7x6 = (Gsy7x6 & Pes7x6);
assign Gsy7x6 = (~(F9s7x6 & Nsy7x6));
assign F9s7x6 = (Usy7x6 & M6j7z6[22]);
assign Usy7x6 = (Ohj7z6[22] & Pes7x6);
assign Sry7x6 = (M6j7z6[23] & Ohj7z6[23]);
assign Bmy7x6 = (Bty7x6 ? Lgj7z6[61] : Lgj7z6[64]);
assign Bty7x6 = (!Zliov6);
assign Zliov6 = (Ity7x6 & Pty7x6);
assign Pty7x6 = (Wty7x6 & Pes7x6);
assign Wty7x6 = (~(Y8s7x6 & Duy7x6));
assign Y8s7x6 = (Kuy7x6 & M6j7z6[20]);
assign Kuy7x6 = (Ohj7z6[20] & Pes7x6);
assign Ity7x6 = (M6j7z6[21] & Ohj7z6[21]);
assign I4v7x6 = (!T6v7x6);
assign T6v7x6 = (Itjov6 ? Yuy7x6 : Ruy7x6);
assign Itjov6 = (!Lrr7x6);
assign Lrr7x6 = (~(Fvy7x6 & Mvy7x6));
assign Mvy7x6 = (~(Tvy7x6 & Awy7x6));
assign Awy7x6 = (~(Hwy7x6 | Owy7x6));
assign Tvy7x6 = (~(Vwy7x6 | Cxy7x6));
assign Fvy7x6 = (~(Jxy7x6 & Qxy7x6));
assign Qxy7x6 = (~(Xxy7x6 | Fft7x6));
assign Fft7x6 = (Eyy7x6 & Lyy7x6);
assign Lyy7x6 = (Syy7x6 & Gsjov6);
assign Eyy7x6 = (~(Zyy7x6 | A4jov6));
assign Xxy7x6 = (Gzy7x6 & Nzy7x6);
assign Nzy7x6 = (Uzy7x6 & B0z7x6);
assign B0z7x6 = (I0z7x6 | Ruy7x6);
assign Gzy7x6 = (P0z7x6 & S9v7x6);
assign S9v7x6 = (Zrr7x6 ? D1z7x6 : W0z7x6);
assign P0z7x6 = (!L9v7x6);
assign L9v7x6 = (~(K1z7x6 & R1z7x6));
assign R1z7x6 = (~(Y1z7x6 & Kujov6));
assign K1z7x6 = (Cqr7x6 ? M2z7x6 : F2z7x6);
assign M2z7x6 = (~(Ptjov6 & T2z7x6));
assign F2z7x6 = (Kujov6 | A3z7x6);
assign Jxy7x6 = (H3z7x6 & O3z7x6);
assign O3z7x6 = (~(V3z7x6 & Ruy7x6));
assign V3z7x6 = (I0z7x6 & Uzy7x6);
assign Uzy7x6 = (C4z7x6 | Gav7x6);
assign H3z7x6 = (~(Gav7x6 & C4z7x6));
assign C4z7x6 = (!Z9v7x6);
assign Z9v7x6 = (Zrr7x6 ? Q4z7x6 : J4z7x6);
assign Gav7x6 = (Ptjov6 ? E5z7x6 : X4z7x6);
assign Yuy7x6 = (!I0z7x6);
assign I0z7x6 = (Ptjov6 ? S5z7x6 : L5z7x6);
assign Ptjov6 = (!Kujov6);
assign Kujov6 = (~(Z5z7x6 & Cxy7x6));
assign Cxy7x6 = (~(G6z7x6 & N6z7x6));
assign N6z7x6 = (U6z7x6 & V3s7x6);
assign G6z7x6 = (~(B7z7x6 | I7z7x6));
assign Z5z7x6 = (~(P7z7x6 & W7z7x6));
assign W7z7x6 = (D8z7x6 & K8z7x6);
assign K8z7x6 = (~(R8z7x6 & Y8z7x6));
assign Y8z7x6 = (F9z7x6 & M9z7x6);
assign F9z7x6 = (~(T9z7x6 & L5z7x6));
assign R8z7x6 = (Aaz7x6 & Y1z7x6);
assign Y1z7x6 = (Rujov6 ? Oaz7x6 : Haz7x6);
assign Aaz7x6 = (Wtjov6 ? A3z7x6 : Vaz7x6);
assign D8z7x6 = (Cbz7x6 | Vwy7x6);
assign Cbz7x6 = (Owy7x6 | Qqr7x6);
assign P7z7x6 = (Jbz7x6 & Qbz7x6);
assign Qbz7x6 = (Xbz7x6 | L5z7x6);
assign Xbz7x6 = (~(S5z7x6 & M9z7x6));
assign M9z7x6 = (~(X4z7x6 & Ecz7x6));
assign Jbz7x6 = (Ecz7x6 | X4z7x6);
assign X4z7x6 = (Qqr7x6 ? Scz7x6 : Lcz7x6);
assign Lcz7x6 = (!Zcz7x6);
assign Ecz7x6 = (!E5z7x6);
assign E5z7x6 = (Cqr7x6 ? Ndz7x6 : Gdz7x6);
assign S5z7x6 = (!T9z7x6);
assign T9z7x6 = (Cqr7x6 ? Bez7x6 : Udz7x6);
assign Cqr7x6 = (!Wtjov6);
assign Wtjov6 = (~(Iez7x6 & B7z7x6));
assign B7z7x6 = (~(Pez7x6 & Wez7x6));
assign Pez7x6 = (~(J5jov6 | Q4s7x6));
assign Iez7x6 = (~(Dfz7x6 & Kfz7x6));
assign Kfz7x6 = (~(Ndz7x6 & Rfz7x6));
assign Ndz7x6 = (!Yfz7x6);
assign Dfz7x6 = (Fgz7x6 & Mgz7x6);
assign Mgz7x6 = (Tgz7x6 | I7z7x6);
assign Fgz7x6 = (~(Ahz7x6 & Hhz7x6));
assign Hhz7x6 = (~(Ohz7x6 & Vhz7x6));
assign Vhz7x6 = (Bez7x6 | Ciz7x6);
assign Ohz7x6 = (~(Jiz7x6 & Vaz7x6));
assign Vaz7x6 = (!T2z7x6);
assign T2z7x6 = (X5jov6 ? Xiz7x6 : Qiz7x6);
assign Jiz7x6 = (~(A3z7x6 | Ejz7x6));
assign Ejz7x6 = (Ciz7x6 & Bez7x6);
assign A3z7x6 = (Zjz7x6 ? Sjz7x6 : Ljz7x6);
assign Sjz7x6 = (U6z7x6 ? Eg8iw6 : Gkz7x6);
assign Ahz7x6 = (~(Gdz7x6 & Yfz7x6));
assign Yfz7x6 = (X5jov6 ? Ukz7x6 : Nkz7x6);
assign Gdz7x6 = (!Rfz7x6);
assign Rfz7x6 = (Zjz7x6 ? Ilz7x6 : Blz7x6);
assign Bez7x6 = (X5jov6 ? Wlz7x6 : Plz7x6);
assign X5jov6 = (~(Dmz7x6 | Wez7x6));
assign Wez7x6 = (~(X4s7x6 | Q5jov6));
assign Dmz7x6 = (Kmz7x6 & Rmz7x6);
assign Rmz7x6 = (J5jov6 | Q4s7x6);
assign Kmz7x6 = (Ymz7x6 & Fnz7x6);
assign Fnz7x6 = (~(Mnz7x6 & Tnz7x6));
assign Tnz7x6 = (Aoz7x6 | Nkz7x6);
assign Mnz7x6 = (~(Hoz7x6 & Ooz7x6));
assign Ooz7x6 = (~(Voz7x6 & Qiz7x6));
assign Qiz7x6 = (J5jov6 ? Lgj7z6[39] : Lgj7z6[36]);
assign Voz7x6 = (~(Xiz7x6 | Cpz7x6));
assign Cpz7x6 = (~(Plz7x6 | Jpz7x6));
assign Xiz7x6 = (Q5jov6 ? Lgj7z6[45] : Lgj7z6[42]);
assign Hoz7x6 = (~(Jpz7x6 & Plz7x6));
assign Ymz7x6 = (~(Nkz7x6 & Aoz7x6));
assign Aoz7x6 = (!Ukz7x6);
assign Ukz7x6 = (Q5jov6 ? Lgj7z6[47] : Lgj7z6[44]);
assign Nkz7x6 = (J5jov6 ? Lgj7z6[41] : Lgj7z6[38]);
assign Wlz7x6 = (!Jpz7x6);
assign Jpz7x6 = (Eqz7x6 ? Xpz7x6 : Qpz7x6);
assign Eqz7x6 = (!Q5jov6);
assign Q5jov6 = (Lqz7x6 & Sqz7x6);
assign Sqz7x6 = (Zqz7x6 & Pes7x6);
assign Zqz7x6 = (~(X4s7x6 & Grz7x6));
assign X4s7x6 = (Nrz7x6 & M6j7z6[14]);
assign Nrz7x6 = (Ohj7z6[14] & Pes7x6);
assign Lqz7x6 = (M6j7z6[15] & Ohj7z6[15]);
assign Plz7x6 = (J5jov6 ? Lgj7z6[40] : Lgj7z6[37]);
assign J5jov6 = (Urz7x6 & Bsz7x6);
assign Bsz7x6 = (Isz7x6 & Pes7x6);
assign Isz7x6 = (~(Q4s7x6 & Psz7x6));
assign Q4s7x6 = (Wsz7x6 & M6j7z6[12]);
assign Wsz7x6 = (Ohj7z6[12] & Pes7x6);
assign Urz7x6 = (M6j7z6[13] & Ohj7z6[13]);
assign Udz7x6 = (!Ciz7x6);
assign Ciz7x6 = (Zjz7x6 ? Ktz7x6 : Dtz7x6);
assign Zjz7x6 = (!Zziov6);
assign Zziov6 = (Rtz7x6 & I7z7x6);
assign I7z7x6 = (C4s7x6 | Sziov6);
assign Rtz7x6 = (~(Ytz7x6 & Tgz7x6));
assign Tgz7x6 = (~(U6z7x6 & V3s7x6));
assign Ytz7x6 = (Fuz7x6 & Muz7x6);
assign Muz7x6 = (~(Tuz7x6 & Avz7x6));
assign Avz7x6 = (Hvz7x6 | Ilz7x6);
assign Tuz7x6 = (~(Ovz7x6 & Vvz7x6));
assign Vvz7x6 = (~(Cwz7x6 & Jwz7x6));
assign Jwz7x6 = (U6z7x6 ? Lgj7z6[24] : Lgj7z6[27]);
assign Cwz7x6 = (Ljz7x6 & Qwz7x6);
assign Qwz7x6 = (Xwz7x6 | Dtz7x6);
assign Ljz7x6 = (Sxz7x6 ? Lxz7x6 : Exz7x6);
assign Ovz7x6 = (~(Dtz7x6 & Xwz7x6));
assign Xwz7x6 = (!Ktz7x6);
assign Fuz7x6 = (~(Ilz7x6 & Hvz7x6));
assign Hvz7x6 = (!Blz7x6);
assign Blz7x6 = (Sziov6 ? Lgj7z6[35] : Lgj7z6[32]);
assign Ilz7x6 = (U6z7x6 ? Lgj7z6[26] : Lgj7z6[29]);
assign Ktz7x6 = (Lziov6 ? Zxz7x6 : Dy7iw6);
assign Lziov6 = (!U6z7x6);
assign U6z7x6 = (~(Gyz7x6 & Nyz7x6));
assign Nyz7x6 = (Uyz7x6 & Pes7x6);
assign Uyz7x6 = (V3s7x6 | Bzz7x6);
assign V3s7x6 = (~(Izz7x6 & M6j7z6[8]));
assign Izz7x6 = (Ohj7z6[8] & Pes7x6);
assign Gyz7x6 = (M6j7z6[9] & Ohj7z6[9]);
assign Dtz7x6 = (Sxz7x6 ? Wzz7x6 : Pzz7x6);
assign Sxz7x6 = (!Sziov6);
assign Sziov6 = (D008x6 & K008x6);
assign K008x6 = (R008x6 & Pes7x6);
assign R008x6 = (~(C4s7x6 & Y008x6));
assign C4s7x6 = (F108x6 & M6j7z6[10]);
assign F108x6 = (Ohj7z6[10] & Pes7x6);
assign D008x6 = (M6j7z6[11] & Ohj7z6[11]);
assign L5z7x6 = (Qqr7x6 ? T108x6 : M108x6);
assign Qqr7x6 = (!Rujov6);
assign Rujov6 = (~(A208x6 & Hwy7x6));
assign Hwy7x6 = (~(H208x6 & O208x6));
assign H208x6 = (~(R2jov6 | F2s7x6));
assign A208x6 = (~(V208x6 & C308x6));
assign C308x6 = (Vwy7x6 | Owy7x6);
assign V208x6 = (J308x6 & Q308x6);
assign Q308x6 = (~(Zcz7x6 & X308x6));
assign X308x6 = (E408x6 | Scz7x6);
assign Zcz7x6 = (Z408x6 ? S408x6 : L408x6);
assign S408x6 = (!G508x6);
assign J308x6 = (~(Scz7x6 & E408x6));
assign E408x6 = (~(N508x6 & U508x6));
assign U508x6 = (B608x6 | Haz7x6);
assign Haz7x6 = (F3jov6 ? P608x6 : I608x6);
assign I608x6 = (W608x6 ? Lgj7z6[12] : Lgj7z6[15]);
assign B608x6 = (~(Oaz7x6 & D708x6));
assign D708x6 = (~(M108x6 & K708x6));
assign Oaz7x6 = (!R708x6);
assign R708x6 = (Z408x6 ? F808x6 : Y708x6);
assign F808x6 = (I1jov6 ? T808x6 : M808x6);
assign N508x6 = (K708x6 | M108x6);
assign Scz7x6 = (F3jov6 ? H908x6 : A908x6);
assign T108x6 = (!K708x6);
assign K708x6 = (F3jov6 ? V908x6 : O908x6);
assign F3jov6 = (~(Ca08x6 | O208x6));
assign O208x6 = (~(Gds7x6 | Y2jov6));
assign Ca08x6 = (Ja08x6 & Qa08x6);
assign Qa08x6 = (Xa08x6 & Eb08x6);
assign Eb08x6 = (~(Lb08x6 & Sb08x6));
assign Sb08x6 = (Zb08x6 & Gc08x6);
assign Zb08x6 = (Nc08x6 | O908x6);
assign Lb08x6 = (~(Uc08x6 | P608x6));
assign P608x6 = (Y2jov6 ? Lgj7z6[21] : Lgj7z6[18]);
assign Uc08x6 = (R2jov6 ? Bd08x6 : Zg8iw6);
assign Xa08x6 = (~(Id08x6 & O908x6));
assign Id08x6 = (Nc08x6 & Gc08x6);
assign Gc08x6 = (H908x6 | Pd08x6);
assign Nc08x6 = (!V908x6);
assign Ja08x6 = (Wd08x6 & De08x6);
assign De08x6 = (~(Pd08x6 & H908x6));
assign H908x6 = (Ye08x6 ? Re08x6 : Ke08x6);
assign Pd08x6 = (!A908x6);
assign A908x6 = (R2jov6 ? Ff08x6 : Ml7iw6);
assign Wd08x6 = (R2jov6 | F2s7x6);
assign V908x6 = (Y2jov6 ? Lgj7z6[22] : Lgj7z6[19]);
assign Y2jov6 = (!Ye08x6);
assign Ye08x6 = (~(Mf08x6 & Tf08x6));
assign Tf08x6 = (Ag08x6 & Pes7x6);
assign Ag08x6 = (~(Gds7x6 & Hg08x6));
assign Gds7x6 = (Og08x6 & M6j7z6[6]);
assign Og08x6 = (Ohj7z6[6] & Pes7x6);
assign Mf08x6 = (M6j7z6[7] & Ohj7z6[7]);
assign O908x6 = (W608x6 ? Lgj7z6[13] : Lgj7z6[16]);
assign W608x6 = (!R2jov6);
assign R2jov6 = (Vg08x6 & Ch08x6);
assign Ch08x6 = (Jh08x6 & Pes7x6);
assign Jh08x6 = (~(F2s7x6 & Qh08x6));
assign F2s7x6 = (Xh08x6 & M6j7z6[4]);
assign Xh08x6 = (Ohj7z6[4] & Pes7x6);
assign Vg08x6 = (M6j7z6[5] & Ohj7z6[5]);
assign M108x6 = (Z408x6 ? Li08x6 : Ei08x6);
assign Z408x6 = (!W1jov6);
assign W1jov6 = (Si08x6 & Owy7x6);
assign Owy7x6 = (J4s7x6 | P1jov6);
assign Si08x6 = (~(Zi08x6 & Gj08x6));
assign Gj08x6 = (Nj08x6 & Vwy7x6);
assign Vwy7x6 = (Y1s7x6 | I1jov6);
assign Nj08x6 = (~(Uj08x6 & Ei08x6));
assign Uj08x6 = (Bk08x6 & Ik08x6);
assign Zi08x6 = (Pk08x6 & Wk08x6);
assign Wk08x6 = (~(Dl08x6 & Kl08x6));
assign Kl08x6 = (Rl08x6 & Ik08x6);
assign Ik08x6 = (~(L408x6 & G508x6));
assign Rl08x6 = (Bk08x6 | Ei08x6);
assign Bk08x6 = (!Li08x6);
assign Dl08x6 = (Yl08x6 & Y708x6);
assign Y708x6 = (Tm08x6 ? Mm08x6 : Fm08x6);
assign Yl08x6 = (An08x6 ? Lgj7z6[0] : Lgj7z6[3]);
assign An08x6 = (!I1jov6);
assign Pk08x6 = (G508x6 | L408x6);
assign L408x6 = (P1jov6 ? Lgj7z6[11] : Lgj7z6[8]);
assign G508x6 = (I1jov6 ? On08x6 : Hn08x6);
assign Li08x6 = (I1jov6 ? Co08x6 : Vn08x6);
assign I1jov6 = (Jo08x6 & Qo08x6);
assign Qo08x6 = (Xo08x6 & Pes7x6);
assign Xo08x6 = (~(Y1s7x6 & Ep08x6));
assign Y1s7x6 = (Lp08x6 & M6j7z6[0]);
assign Lp08x6 = (Ohj7z6[0] & Pes7x6);
assign Jo08x6 = (M6j7z6[1] & Ohj7z6[1]);
assign Ei08x6 = (Tm08x6 ? Zp08x6 : Sp08x6);
assign Tm08x6 = (!P1jov6);
assign P1jov6 = (Gq08x6 & Nq08x6);
assign Nq08x6 = (Uq08x6 & Pes7x6);
assign Uq08x6 = (~(J4s7x6 & Br08x6));
assign J4s7x6 = (Ir08x6 & M6j7z6[2]);
assign Ir08x6 = (Ohj7z6[2] & Pes7x6);
assign Gq08x6 = (M6j7z6[3] & Ohj7z6[3]);
assign Ruy7x6 = (Zrr7x6 ? Wr08x6 : Pr08x6);
assign Zrr7x6 = (!Srr7x6);
assign Srr7x6 = (~(Ds08x6 & Zyy7x6));
assign Zyy7x6 = (~(Ks08x6 & Rs08x6));
assign Ks08x6 = (Srjov6 & Yseov6);
assign Yseov6 = (!Z3j7z6[15]);
assign Ds08x6 = (~(Ys08x6 & Ft08x6));
assign Ft08x6 = (~(Fvjov6 & Mt08x6));
assign Ys08x6 = (Tt08x6 & Au08x6);
assign Au08x6 = (~(Q4z7x6 & Hu08x6));
assign Hu08x6 = (Ou08x6 | Vu08x6);
assign Q4z7x6 = (S6jov6 ? Jv08x6 : Cv08x6);
assign Tt08x6 = (~(Vu08x6 & Ou08x6));
assign Ou08x6 = (!J4z7x6);
assign J4z7x6 = (Qv08x6 & Xv08x6);
assign Xv08x6 = (~(Jyiov6 & Ew08x6));
assign Qv08x6 = (Err7x6 ? Sw08x6 : Lw08x6);
assign Sw08x6 = (Gsjov6 | Zw08x6);
assign Lw08x6 = (~(Fvjov6 & Gx08x6));
assign Vu08x6 = (~(Nx08x6 & Ux08x6));
assign Ux08x6 = (By08x6 | D1z7x6);
assign D1z7x6 = (S6jov6 ? Iy08x6 : Gaj7z6[0]);
assign By08x6 = (~(Py08x6 & W0z7x6));
assign W0z7x6 = (~(Wy08x6 & Dz08x6));
assign Dz08x6 = (~(Kz08x6 & Jyiov6));
assign Jyiov6 = (Err7x6 & Gsjov6);
assign Wy08x6 = (Err7x6 ? Yz08x6 : Rz08x6);
assign Yz08x6 = (Gsjov6 | F018x6);
assign Rz08x6 = (~(Fvjov6 & M018x6));
assign Py08x6 = (~(T018x6 & Wr08x6));
assign Nx08x6 = (Wr08x6 | T018x6);
assign Wr08x6 = (S6jov6 ? A118x6 : Gaj7z6[1]);
assign S6jov6 = (H118x6 & O118x6);
assign O118x6 = (~(V118x6 & Z3j7z6[15]));
assign V118x6 = (C218x6 & J218x6);
assign J218x6 = (~(Jv08x6 & Q218x6));
assign Q218x6 = (~(X218x6 & E318x6));
assign X218x6 = (L318x6 & Cv08x6);
assign Jv08x6 = (Srjov6 ? Z318x6 : S318x6);
assign C218x6 = (~(Gaj7z6[2] & G418x6));
assign G418x6 = (~(L318x6 & E318x6));
assign E318x6 = (A118x6 | N418x6);
assign L318x6 = (U418x6 | Iy08x6);
assign Iy08x6 = (G7jov6 ? B518x6 : Nbj7z6[0]);
assign U418x6 = (~(Gaj7z6[0] & I518x6));
assign I518x6 = (~(A118x6 & N418x6));
assign H118x6 = (~(Srjov6 & Rs08x6));
assign Rs08x6 = (Vueov6 | Oreet6);
assign Vueov6 = (!Oecet6);
assign A118x6 = (G7jov6 ? P518x6 : Nbj7z6[1]);
assign G7jov6 = (!Srjov6);
assign Srjov6 = (~(W518x6 & D618x6));
assign D618x6 = (~(K618x6 & R618x6));
assign R618x6 = (Y618x6 & F718x6);
assign F718x6 = (~(M718x6 & T718x6));
assign T718x6 = (A818x6 & H818x6);
assign A818x6 = (O818x6 | Nbj7z6[1]);
assign M718x6 = (~(B518x6 | Cehov6));
assign B518x6 = (V818x6 ? Z8j7z6[0] : T7j7z6[0]);
assign Y618x6 = (~(C918x6 & Nbj7z6[1]));
assign C918x6 = (O818x6 & H818x6);
assign H818x6 = (S318x6 | Nbj7z6[2]);
assign O818x6 = (!P518x6);
assign K618x6 = (Oecet6 & J918x6);
assign J918x6 = (~(S318x6 & Nbj7z6[2]));
assign S318x6 = (N7jov6 ? X918x6 : Q918x6);
assign W518x6 = (Ea18x6 & Pes7x6);
assign Pes7x6 = (!Oreet6);
assign Ea18x6 = (~(G5eov6 & V818x6));
assign G5eov6 = (!Fhcet6);
assign P518x6 = (N7jov6 ? T7j7z6[1] : Z8j7z6[1]);
assign N7jov6 = (!V818x6);
assign V818x6 = (~(Zfcet6 & La18x6));
assign La18x6 = (~(Fhcet6 & Sa18x6));
assign Pr08x6 = (!T018x6);
assign T018x6 = (Err7x6 ? Gb18x6 : Za18x6);
assign Err7x6 = (!Mt08x6);
assign Mt08x6 = (~(Fvjov6 & Nb18x6));
assign Nb18x6 = (~(Syy7x6 & Gsjov6));
assign Syy7x6 = (~(Qyiov6 | K1s7x6));
assign Gb18x6 = (Gsjov6 ? Bc18x6 : Ub18x6);
assign Gsjov6 = (~(Ic18x6 & Micet6));
assign Ic18x6 = (Z3j7z6[12] & Pc18x6);
assign Pc18x6 = (~(Wc18x6 & Dd18x6));
assign Dd18x6 = (Kd18x6 & Rd18x6);
assign Rd18x6 = (~(Yd18x6 & Fe18x6));
assign Fe18x6 = (Me18x6 & F018x6);
assign Yd18x6 = (Kz08x6 & Te18x6);
assign Te18x6 = (Af18x6 | Ub18x6);
assign Kz08x6 = (Qyiov6 ? Zdj7z6[0] : Ffj7z6[0]);
assign Kd18x6 = (~(Hf18x6 & Af18x6));
assign Hf18x6 = (Me18x6 & Ub18x6);
assign Me18x6 = (Ew08x6 | Zw08x6);
assign Wc18x6 = (Of18x6 & Vf18x6);
assign Vf18x6 = (~(Ew08x6 & Zw08x6));
assign Ew08x6 = (Qyiov6 ? Zdj7z6[2] : Ffj7z6[2]);
assign Of18x6 = (Qyiov6 | K1s7x6);
assign Bc18x6 = (!Af18x6);
assign Af18x6 = (Qyiov6 ? Zdj7z6[1] : Ffj7z6[1]);
assign Qyiov6 = (Cg18x6 & Z3j7z6[14]);
assign Cg18x6 = (Sjcet6 & Jg18x6);
assign Jg18x6 = (~(K1s7x6 & Qg18x6));
assign K1s7x6 = (Z3j7z6[13] & Ykcet6);
assign Za18x6 = (A4jov6 | Xg18x6);
assign A4jov6 = (!Fvjov6);
assign Fvjov6 = (Nxeov6 & Uxeov6);
assign Uxeov6 = (!V5get6);
assign Nxeov6 = (!Hdcet6);
assign Pzs7x6 = (Izs7x6 | Inadt6);
assign K9r7x6 = (Eh18x6 & Iwa7x6);
assign Iwa7x6 = (!Lh18x6);
assign Eh18x6 = (~(Bxi7z6[1] & Sh18x6));
assign Sh18x6 = (~(O8fov6 & B52nv6));
assign O8fov6 = (Yhc7x6 & Zh18x6);
assign Yhc7x6 = (Eec7x6 & Pb8iw6);
assign V3w7v6 = (~(Gi18x6 & Ni18x6));
assign Ni18x6 = (~(Fjb7z6[2] & Lriiw6));
assign Gi18x6 = (~(Ui18x6 & Bj18x6));
assign Bj18x6 = (Ij18x6 & Pj18x6);
assign Pj18x6 = (Wj18x6 | Te2nv6);
assign Wj18x6 = (Dk18x6 & Kk18x6);
assign Ij18x6 = (~(Yd2nv6 | A0fet6));
assign Ui18x6 = (Rk18x6 & Sriiw6);
assign Rk18x6 = (E1cet6 & Yk18x6);
assign Yk18x6 = (~(Lunov6 & Nmadt6));
assign O3w7v6 = (~(Fl18x6 & Ml18x6));
assign Ml18x6 = (~(Nxm7x6 & Tteov6));
assign Fl18x6 = (Tl18x6 & Am18x6);
assign Am18x6 = (~(Ohj7z6[0] & Hm18x6));
assign Hm18x6 = (~(Om18x6 & Vm18x6));
assign Vm18x6 = (Cn18x6 & Jn18x6);
assign Cn18x6 = (~(Qn18x6 & Xn18x6));
assign Xn18x6 = (Eo18x6 & M808x6);
assign Eo18x6 = (~(Lgj7z6[2] & Lo18x6));
assign Qn18x6 = (So18x6 & Zo18x6);
assign Zo18x6 = (~(Gp18x6 & Lgj7z6[1]));
assign Om18x6 = (Np18x6 & Up18x6);
assign Up18x6 = (~(Bq18x6 & Vn08x6));
assign Bq18x6 = (~(Iq18x6 & Pq18x6));
assign Pq18x6 = (~(Wq18x6 & Hn08x6));
assign Hn08x6 = (!Lgj7z6[2]);
assign Np18x6 = (Dr18x6 | Lgj7z6[2]);
assign Tl18x6 = (~(Fjb7z6[3] & Lriiw6));
assign H3w7v6 = (~(Kr18x6 & Rr18x6));
assign Rr18x6 = (~(Nxm7x6 & Cheov6));
assign Kr18x6 = (Yr18x6 & Fs18x6);
assign Fs18x6 = (~(Ohj7z6[1] & Ms18x6));
assign Ms18x6 = (~(Ts18x6 & At18x6));
assign At18x6 = (Ht18x6 & Jn18x6);
assign Ht18x6 = (~(Ot18x6 & Vt18x6));
assign Vt18x6 = (Cu18x6 & T808x6);
assign Cu18x6 = (~(Lgj7z6[5] & Lo18x6));
assign Ot18x6 = (So18x6 & Ju18x6);
assign Ju18x6 = (~(Gp18x6 & Lgj7z6[4]));
assign Ts18x6 = (Qu18x6 & Xu18x6);
assign Xu18x6 = (~(Ev18x6 & On08x6));
assign Ev18x6 = (~(Dr18x6 & Lv18x6));
assign Lv18x6 = (~(Wq18x6 & Co08x6));
assign Qu18x6 = (Iq18x6 | Lgj7z6[4]);
assign Yr18x6 = (~(Fjb7z6[4] & Lriiw6));
assign A3w7v6 = (~(Sv18x6 & Zv18x6));
assign Zv18x6 = (~(Nxm7x6 & Breov6));
assign Sv18x6 = (Gw18x6 & Nw18x6);
assign Nw18x6 = (~(Ohj7z6[2] & Uw18x6));
assign Uw18x6 = (~(Bx18x6 & Ix18x6));
assign Ix18x6 = (Px18x6 & Jn18x6);
assign Px18x6 = (~(Wx18x6 & Dy18x6));
assign Dy18x6 = (Ky18x6 & Mm08x6);
assign Ky18x6 = (~(Lgj7z6[8] & Lo18x6));
assign Wx18x6 = (So18x6 & Ry18x6);
assign Ry18x6 = (~(Gp18x6 & Lgj7z6[7]));
assign Bx18x6 = (Yy18x6 & Fz18x6);
assign Fz18x6 = (~(Mz18x6 & Zp08x6));
assign Mz18x6 = (~(Iq18x6 & Tz18x6));
assign Tz18x6 = (~(Wq18x6 & A028x6));
assign Yy18x6 = (Dr18x6 | Lgj7z6[8]);
assign Gw18x6 = (~(Fjb7z6[5] & Lriiw6));
assign T2w7v6 = (~(H028x6 & O028x6));
assign O028x6 = (~(Nxm7x6 & Vgeov6));
assign H028x6 = (V028x6 & C128x6);
assign C128x6 = (~(Ohj7z6[3] & J128x6));
assign J128x6 = (~(Q128x6 & X128x6));
assign X128x6 = (E228x6 & Jn18x6);
assign E228x6 = (~(L228x6 & S228x6));
assign S228x6 = (Z228x6 & Fm08x6);
assign Z228x6 = (~(Lgj7z6[11] & Lo18x6));
assign L228x6 = (So18x6 & G328x6);
assign G328x6 = (~(Gp18x6 & Lgj7z6[10]));
assign Q128x6 = (N328x6 & U328x6);
assign U328x6 = (~(B428x6 & I428x6));
assign B428x6 = (~(Dr18x6 & P428x6));
assign P428x6 = (~(Wq18x6 & Sp08x6));
assign N328x6 = (Iq18x6 | Lgj7z6[10]);
assign V028x6 = (~(Fjb7z6[6] & Lriiw6));
assign M2w7v6 = (~(W428x6 & D528x6));
assign D528x6 = (~(Nxm7x6 & Uqeov6));
assign W428x6 = (K528x6 & R528x6);
assign R528x6 = (~(Ohj7z6[4] & Y528x6));
assign Y528x6 = (~(F628x6 & M628x6));
assign M628x6 = (T628x6 & Jn18x6);
assign T628x6 = (~(A728x6 & H728x6));
assign H728x6 = (O728x6 & Zg8iw6);
assign O728x6 = (~(Lgj7z6[14] & Lo18x6));
assign A728x6 = (So18x6 & V728x6);
assign V728x6 = (~(Gp18x6 & Lgj7z6[13]));
assign F628x6 = (C828x6 & J828x6);
assign J828x6 = (~(Q828x6 & Yy7iw6));
assign Q828x6 = (~(Iq18x6 & X828x6));
assign X828x6 = (~(Wq18x6 & Ml7iw6));
assign Ml7iw6 = (!Lgj7z6[14]);
assign C828x6 = (Dr18x6 | Lgj7z6[14]);
assign K528x6 = (~(Fjb7z6[7] & Lriiw6));
assign F2w7v6 = (~(E928x6 & L928x6));
assign L928x6 = (~(Nxm7x6 & Yeeov6));
assign E928x6 = (S928x6 & Z928x6);
assign Z928x6 = (~(Ohj7z6[5] & Ga28x6));
assign Ga28x6 = (~(Na28x6 & Ua28x6));
assign Ua28x6 = (Bb28x6 & Jn18x6);
assign Bb28x6 = (~(Ib28x6 & Pb28x6));
assign Pb28x6 = (Wb28x6 & Bd08x6);
assign Wb28x6 = (~(Lgj7z6[17] & Lo18x6));
assign Ib28x6 = (So18x6 & Dc28x6);
assign Dc28x6 = (~(Gp18x6 & Lgj7z6[16]));
assign Na28x6 = (Kc28x6 & Rc28x6);
assign Rc28x6 = (~(Yc28x6 & Ff08x6));
assign Yc28x6 = (~(Dr18x6 & Fd28x6));
assign Fd28x6 = (~(Wq18x6 & Md28x6));
assign Kc28x6 = (Iq18x6 | Lgj7z6[16]);
assign S928x6 = (~(Fjb7z6[8] & Lriiw6));
assign Y1w7v6 = (~(Td28x6 & Ae28x6));
assign Ae28x6 = (~(Nxm7x6 & Zpeov6));
assign Td28x6 = (He28x6 & Oe28x6);
assign Oe28x6 = (~(Ohj7z6[6] & Ve28x6));
assign Ve28x6 = (~(Cf28x6 & Jf28x6));
assign Jf28x6 = (Qf28x6 & Jn18x6);
assign Qf28x6 = (~(Xf28x6 & Eg28x6));
assign Eg28x6 = (Lg28x6 & Sg28x6);
assign Lg28x6 = (~(Lgj7z6[20] & Lo18x6));
assign Xf28x6 = (So18x6 & Zg28x6);
assign Zg28x6 = (~(Gp18x6 & Lgj7z6[19]));
assign Cf28x6 = (Gh28x6 & Nh28x6);
assign Nh28x6 = (~(Uh28x6 & Bi28x6));
assign Uh28x6 = (~(Iq18x6 & Ii28x6));
assign Ii28x6 = (~(Wq18x6 & Re08x6));
assign Re08x6 = (!Lgj7z6[20]);
assign Gh28x6 = (Dr18x6 | Lgj7z6[20]);
assign He28x6 = (~(Fjb7z6[9] & Lriiw6));
assign R1w7v6 = (~(Pi28x6 & Wi28x6));
assign Wi28x6 = (~(Nxm7x6 & Ageov6));
assign Pi28x6 = (Dj28x6 & Kj28x6);
assign Kj28x6 = (~(Ohj7z6[7] & Rj28x6));
assign Rj28x6 = (~(Yj28x6 & Fk28x6));
assign Fk28x6 = (Mk28x6 & Jn18x6);
assign Mk28x6 = (~(Tk28x6 & Al28x6));
assign Al28x6 = (Hl28x6 & Ol28x6);
assign Hl28x6 = (~(Lgj7z6[23] & Lo18x6));
assign Tk28x6 = (So18x6 & Vl28x6);
assign Vl28x6 = (~(Gp18x6 & Lgj7z6[22]));
assign Yj28x6 = (Cm28x6 & Jm28x6);
assign Jm28x6 = (~(Qm28x6 & Ke08x6));
assign Qm28x6 = (~(Dr18x6 & Xm28x6));
assign Xm28x6 = (~(Wq18x6 & En28x6));
assign Cm28x6 = (Iq18x6 | Lgj7z6[22]);
assign Dj28x6 = (~(Fjb7z6[10] & Lriiw6));
assign K1w7v6 = (~(Ln28x6 & Sn28x6));
assign Sn28x6 = (~(Nxm7x6 & E4eov6));
assign Ln28x6 = (Zn28x6 & Go28x6);
assign Go28x6 = (~(Ohj7z6[8] & No28x6));
assign No28x6 = (~(Uo28x6 & Bp28x6));
assign Bp28x6 = (Ip28x6 & Jn18x6);
assign Ip28x6 = (~(Pp28x6 & Wp28x6));
assign Wp28x6 = (Dq28x6 & Eg8iw6);
assign Dq28x6 = (~(Lgj7z6[26] & Lo18x6));
assign Pp28x6 = (So18x6 & Kq28x6);
assign Kq28x6 = (~(Gp18x6 & Lgj7z6[25]));
assign Uo28x6 = (Rq28x6 & Yq28x6);
assign Yq28x6 = (~(Fr28x6 & Dy7iw6));
assign Fr28x6 = (~(Iq18x6 & Mr28x6));
assign Mr28x6 = (~(Wq18x6 & Kk7iw6));
assign Rq28x6 = (Dr18x6 | Lgj7z6[26]);
assign Zn28x6 = (~(Fjb7z6[11] & Lriiw6));
assign D1w7v6 = (~(Tr28x6 & As28x6));
assign As28x6 = (~(Nxm7x6 & X3eov6));
assign Tr28x6 = (Hs28x6 & Os28x6);
assign Os28x6 = (~(Ohj7z6[9] & Vs28x6));
assign Vs28x6 = (~(Ct28x6 & Jt28x6));
assign Jt28x6 = (Qt28x6 & Jn18x6);
assign Qt28x6 = (~(Xt28x6 & Eu28x6));
assign Eu28x6 = (Lu28x6 & Gkz7x6);
assign Lu28x6 = (~(Lgj7z6[29] & Lo18x6));
assign Xt28x6 = (So18x6 & Su28x6);
assign Su28x6 = (~(Gp18x6 & Lgj7z6[28]));
assign Ct28x6 = (Zu28x6 & Gv28x6);
assign Gv28x6 = (~(Nv28x6 & Uv28x6));
assign Nv28x6 = (~(Dr18x6 & Bw28x6));
assign Bw28x6 = (~(Wq18x6 & Zxz7x6));
assign Zu28x6 = (Iq18x6 | Lgj7z6[28]);
assign Hs28x6 = (~(Fjb7z6[12] & Lriiw6));
assign W0w7v6 = (~(Iw28x6 & Pw28x6));
assign Pw28x6 = (~(Nxm7x6 & O2eov6));
assign Iw28x6 = (Ww28x6 & Dx28x6);
assign Dx28x6 = (~(Ohj7z6[10] & Kx28x6));
assign Kx28x6 = (~(Rx28x6 & Yx28x6));
assign Yx28x6 = (Fy28x6 & Jn18x6);
assign Fy28x6 = (~(My28x6 & Ty28x6));
assign Ty28x6 = (Az28x6 & Lxz7x6);
assign Az28x6 = (~(Lgj7z6[32] & Lo18x6));
assign My28x6 = (So18x6 & Hz28x6);
assign Hz28x6 = (~(Gp18x6 & Lgj7z6[31]));
assign Rx28x6 = (Oz28x6 & Vz28x6);
assign Vz28x6 = (~(C038x6 & Wzz7x6));
assign C038x6 = (~(Iq18x6 & J038x6));
assign J038x6 = (~(Wq18x6 & Q038x6));
assign Oz28x6 = (Dr18x6 | Lgj7z6[32]);
assign Ww28x6 = (~(Fjb7z6[13] & Lriiw6));
assign P0w7v6 = (~(X038x6 & E138x6));
assign E138x6 = (~(Nxm7x6 & H2eov6));
assign X038x6 = (L138x6 & S138x6);
assign S138x6 = (~(Ohj7z6[11] & Z138x6));
assign Z138x6 = (~(G238x6 & N238x6));
assign N238x6 = (U238x6 & Jn18x6);
assign U238x6 = (~(B338x6 & I338x6));
assign I338x6 = (P338x6 & Exz7x6);
assign P338x6 = (~(Lgj7z6[35] & Lo18x6));
assign B338x6 = (So18x6 & W338x6);
assign W338x6 = (~(Gp18x6 & Lgj7z6[34]));
assign G238x6 = (D438x6 & K438x6);
assign K438x6 = (~(R438x6 & Y438x6));
assign R438x6 = (~(Dr18x6 & F538x6));
assign F538x6 = (~(Wq18x6 & Pzz7x6));
assign D438x6 = (Iq18x6 | Lgj7z6[34]);
assign L138x6 = (~(Fjb7z6[14] & Lriiw6));
assign I0w7v6 = (~(M538x6 & T538x6));
assign T538x6 = (~(Nxm7x6 & K0eov6));
assign M538x6 = (A638x6 & H638x6);
assign H638x6 = (~(Ohj7z6[12] & O638x6));
assign O638x6 = (~(V638x6 & C738x6));
assign C738x6 = (J738x6 & Jn18x6);
assign J738x6 = (~(Q738x6 & X738x6));
assign X738x6 = (~(E838x6 | Lgj7z6[36]));
assign E838x6 = (Lgj7z6[38] & Lo18x6);
assign Q738x6 = (So18x6 & L838x6);
assign L838x6 = (~(Gp18x6 & Lgj7z6[37]));
assign V638x6 = (S838x6 & Z838x6);
assign Z838x6 = (~(G938x6 & N938x6));
assign G938x6 = (~(Iq18x6 & U938x6));
assign U938x6 = (Ba38x6 | Lgj7z6[38]);
assign S838x6 = (Dr18x6 | Lgj7z6[38]);
assign A638x6 = (~(Fjb7z6[15] & Lriiw6));
assign B0w7v6 = (~(Ia38x6 & Pa38x6));
assign Pa38x6 = (~(Nxm7x6 & M1eov6));
assign Ia38x6 = (Wa38x6 & Db38x6);
assign Db38x6 = (~(Ohj7z6[13] & Kb38x6));
assign Kb38x6 = (~(Rb38x6 & Yb38x6));
assign Yb38x6 = (Fc38x6 & Jn18x6);
assign Fc38x6 = (~(Mc38x6 & Tc38x6));
assign Tc38x6 = (Ad38x6 & Hd38x6);
assign Ad38x6 = (~(Lgj7z6[41] & Lo18x6));
assign Mc38x6 = (So18x6 & Od38x6);
assign Od38x6 = (~(Gp18x6 & Lgj7z6[40]));
assign Rb38x6 = (Vd38x6 & Ce38x6);
assign Ce38x6 = (~(Je38x6 & Qe38x6));
assign Je38x6 = (~(Dr18x6 & Xe38x6));
assign Xe38x6 = (~(Wq18x6 & Ef38x6));
assign Vd38x6 = (Iq18x6 | Lgj7z6[40]);
assign Wa38x6 = (~(Fjb7z6[16] & Lriiw6));
assign Uzv7v6 = (~(Lf38x6 & Sf38x6));
assign Sf38x6 = (~(Nxm7x6 & F1eov6));
assign Lf38x6 = (Zf38x6 & Gg38x6);
assign Gg38x6 = (~(Ohj7z6[14] & Ng38x6));
assign Ng38x6 = (~(Ug38x6 & Bh38x6));
assign Bh38x6 = (Ih38x6 & Jn18x6);
assign Ih38x6 = (~(Ph38x6 & Wh38x6));
assign Wh38x6 = (Di38x6 & Ki38x6);
assign Di38x6 = (~(Lgj7z6[44] & Lo18x6));
assign Ph38x6 = (So18x6 & Ri38x6);
assign Ri38x6 = (~(Gp18x6 & Lgj7z6[43]));
assign Ug38x6 = (Yi38x6 & Fj38x6);
assign Fj38x6 = (~(Mj38x6 & Xpz7x6));
assign Mj38x6 = (~(Iq18x6 & Tj38x6));
assign Tj38x6 = (~(Wq18x6 & Ak38x6));
assign Yi38x6 = (Dr18x6 | Lgj7z6[44]);
assign Zf38x6 = (~(Fjb7z6[17] & Lriiw6));
assign Nzv7v6 = (~(Hk38x6 & Ok38x6));
assign Ok38x6 = (~(Nxm7x6 & Nydov6));
assign Hk38x6 = (Vk38x6 & Cl38x6);
assign Cl38x6 = (~(Ohj7z6[15] & Jl38x6));
assign Jl38x6 = (~(Ql38x6 & Xl38x6));
assign Xl38x6 = (Em38x6 & Jn18x6);
assign Em38x6 = (~(Lm38x6 & Sm38x6));
assign Sm38x6 = (Zm38x6 & Gn38x6);
assign Zm38x6 = (~(Lgj7z6[47] & Lo18x6));
assign Lm38x6 = (So18x6 & Nn38x6);
assign Nn38x6 = (~(Gp18x6 & Lgj7z6[46]));
assign Ql38x6 = (Un38x6 & Bo38x6);
assign Bo38x6 = (~(Io38x6 & Po38x6));
assign Io38x6 = (~(Dr18x6 & Wo38x6));
assign Wo38x6 = (~(Wq18x6 & Qpz7x6));
assign Un38x6 = (Iq18x6 | Lgj7z6[46]);
assign Vk38x6 = (~(Fjb7z6[18] & Lriiw6));
assign Gzv7v6 = (~(Dp38x6 & Kp38x6));
assign Kp38x6 = (~(Nxm7x6 & Speov6));
assign Dp38x6 = (Rp38x6 & Yp38x6);
assign Yp38x6 = (~(Ohj7z6[16] & Fq38x6));
assign Fq38x6 = (~(Mq38x6 & Tq38x6));
assign Tq38x6 = (Ar38x6 & Jn18x6);
assign Ar38x6 = (~(Hr38x6 & Or38x6));
assign Or38x6 = (Vr38x6 & Jcy7x6);
assign Vr38x6 = (~(Lgj7z6[50] & Lo18x6));
assign Hr38x6 = (So18x6 & Cs38x6);
assign Cs38x6 = (~(Gp18x6 & Lgj7z6[49]));
assign Mq38x6 = (Js38x6 & Qs38x6);
assign Qs38x6 = (~(Xs38x6 & Lky7x6));
assign Xs38x6 = (~(Iq18x6 & Et38x6));
assign Et38x6 = (Ba38x6 | Lgj7z6[50]);
assign Js38x6 = (Dr18x6 | Lgj7z6[50]);
assign Rp38x6 = (~(Fjb7z6[19] & Lriiw6));
assign Zyv7v6 = (~(Lt38x6 & St38x6));
assign St38x6 = (~(Nxm7x6 & Tfeov6));
assign Lt38x6 = (Zt38x6 & Gu38x6);
assign Gu38x6 = (~(Ohj7z6[17] & Nu38x6));
assign Nu38x6 = (~(Uu38x6 & Bv38x6));
assign Bv38x6 = (Iv38x6 & Jn18x6);
assign Iv38x6 = (~(Pv38x6 & Wv38x6));
assign Wv38x6 = (Dw38x6 & Ccy7x6);
assign Dw38x6 = (~(Lgj7z6[53] & Lo18x6));
assign Pv38x6 = (So18x6 & Kw38x6);
assign Kw38x6 = (~(Gp18x6 & Lgj7z6[52]));
assign Uu38x6 = (Rw38x6 & Yw38x6);
assign Yw38x6 = (~(Fx38x6 & Mx38x6));
assign Fx38x6 = (~(Dr18x6 & Tx38x6));
assign Tx38x6 = (Ba38x6 | Lgj7z6[52]);
assign Rw38x6 = (Iq18x6 | Lgj7z6[52]);
assign Zt38x6 = (~(Fjb7z6[20] & Lriiw6));
assign Syv7v6 = (~(Ay38x6 & Hy38x6));
assign Hy38x6 = (~(Nxm7x6 & Joeov6));
assign Ay38x6 = (Oy38x6 & Vy38x6);
assign Vy38x6 = (~(Ohj7z6[18] & Cz38x6));
assign Cz38x6 = (~(Jz38x6 & Qz38x6));
assign Qz38x6 = (Xz38x6 & Jn18x6);
assign Xz38x6 = (~(E048x6 & L048x6));
assign L048x6 = (S048x6 & Fhy7x6);
assign S048x6 = (~(Lgj7z6[56] & Lo18x6));
assign E048x6 = (So18x6 & Z048x6);
assign Z048x6 = (~(Gp18x6 & Lgj7z6[55]));
assign Jz38x6 = (G148x6 & N148x6);
assign N148x6 = (~(U148x6 & Viy7x6));
assign U148x6 = (~(Iq18x6 & B248x6));
assign B248x6 = (Ba38x6 | Lgj7z6[56]);
assign G148x6 = (Dr18x6 | Lgj7z6[56]);
assign Oy38x6 = (~(Fjb7z6[21] & Lriiw6));
assign Lyv7v6 = (~(I248x6 & P248x6));
assign P248x6 = (~(Nxm7x6 & Bdeov6));
assign I248x6 = (W248x6 & D348x6);
assign D348x6 = (~(Ohj7z6[19] & K348x6));
assign K348x6 = (~(R348x6 & Y348x6));
assign Y348x6 = (F448x6 & Jn18x6);
assign F448x6 = (~(M448x6 & T448x6));
assign T448x6 = (A548x6 & Ygy7x6);
assign A548x6 = (~(Lgj7z6[59] & Lo18x6));
assign M448x6 = (So18x6 & H548x6);
assign H548x6 = (~(Gp18x6 & Lgj7z6[58]));
assign R348x6 = (O548x6 & V548x6);
assign V548x6 = (~(C648x6 & J648x6));
assign C648x6 = (~(Dr18x6 & Q648x6));
assign Q648x6 = (Ba38x6 | Lgj7z6[58]);
assign O548x6 = (Iq18x6 | Lgj7z6[58]);
assign W248x6 = (~(Fjb7z6[22] & Lriiw6));
assign Eyv7v6 = (~(X648x6 & E748x6));
assign E748x6 = (~(Nxm7x6 & Coeov6));
assign X648x6 = (L748x6 & S748x6);
assign S748x6 = (~(Ohj7z6[20] & Z748x6));
assign Z748x6 = (~(G848x6 & N848x6));
assign N848x6 = (U848x6 & Jn18x6);
assign U848x6 = (~(B948x6 & I948x6));
assign I948x6 = (P948x6 & Ae8iw6);
assign Ae8iw6 = (!Lgj7z6[60]);
assign P948x6 = (~(Lgj7z6[62] & Lo18x6));
assign B948x6 = (So18x6 & W948x6);
assign W948x6 = (~(Gp18x6 & Lgj7z6[61]));
assign G848x6 = (Da48x6 & Ka48x6);
assign Ka48x6 = (~(Ra48x6 & Gw7iw6));
assign Ra48x6 = (~(Iq18x6 & Ya48x6));
assign Ya48x6 = (Ba38x6 | Lgj7z6[62]);
assign Da48x6 = (Dr18x6 | Lgj7z6[62]);
assign L748x6 = (~(Fjb7z6[23] & Lriiw6));
assign Xxv7v6 = (~(Fb48x6 & Mb48x6));
assign Mb48x6 = (~(Nxm7x6 & Uceov6));
assign Fb48x6 = (Tb48x6 & Ac48x6);
assign Ac48x6 = (~(Ohj7z6[21] & Hc48x6));
assign Hc48x6 = (~(Oc48x6 & Vc48x6));
assign Vc48x6 = (Cd48x6 & Jn18x6);
assign Cd48x6 = (~(Jd48x6 & Qd48x6));
assign Qd48x6 = (Xd48x6 & Qqy7x6);
assign Qqy7x6 = (!Lgj7z6[63]);
assign Xd48x6 = (~(Lgj7z6[65] & Lo18x6));
assign Jd48x6 = (So18x6 & Ee48x6);
assign Ee48x6 = (~(Gp18x6 & Lgj7z6[64]));
assign Oc48x6 = (Le48x6 & Se48x6);
assign Se48x6 = (~(Ze48x6 & Lry7x6));
assign Ze48x6 = (~(Dr18x6 & Gf48x6));
assign Gf48x6 = (Ba38x6 | Lgj7z6[64]);
assign Le48x6 = (Iq18x6 | Lgj7z6[64]);
assign Tb48x6 = (~(Fjb7z6[24] & Lriiw6));
assign Qxv7v6 = (~(Nf48x6 & Uf48x6));
assign Uf48x6 = (~(Nxm7x6 & Fmeov6));
assign Nf48x6 = (Bg48x6 & Ig48x6);
assign Ig48x6 = (~(Ohj7z6[22] & Pg48x6));
assign Pg48x6 = (~(Wg48x6 & Dh48x6));
assign Dh48x6 = (Kh48x6 & Jn18x6);
assign Kh48x6 = (~(Rh48x6 & Yh48x6));
assign Yh48x6 = (Fi48x6 & May7x6);
assign Fi48x6 = (~(Lgj7z6[68] & Lo18x6));
assign Rh48x6 = (So18x6 & Mi48x6);
assign Mi48x6 = (~(Gp18x6 & Lgj7z6[67]));
assign Wg48x6 = (Ti48x6 & Aj48x6);
assign Aj48x6 = (~(Hj48x6 & Oj48x6));
assign Hj48x6 = (~(Iq18x6 & Vj48x6));
assign Vj48x6 = (Ba38x6 | Lgj7z6[68]);
assign Ti48x6 = (Dr18x6 | Lgj7z6[68]);
assign Bg48x6 = (~(Fjb7z6[25] & Lriiw6));
assign Jxv7v6 = (~(Ck48x6 & Jk48x6));
assign Jk48x6 = (~(Nxm7x6 & Zbeov6));
assign Ck48x6 = (Qk48x6 & Xk48x6);
assign Xk48x6 = (~(Ohj7z6[23] & El48x6));
assign El48x6 = (~(Ll48x6 & Sl48x6));
assign Sl48x6 = (Zl48x6 & Jn18x6);
assign Zl48x6 = (~(Gm48x6 & Nm48x6));
assign Nm48x6 = (Um48x6 & Tay7x6);
assign Um48x6 = (~(Lgj7z6[71] & Lo18x6));
assign Gm48x6 = (So18x6 & Bn48x6);
assign Bn48x6 = (~(Gp18x6 & Lgj7z6[70]));
assign Ll48x6 = (In48x6 & Pn48x6);
assign Pn48x6 = (~(Wn48x6 & Xqy7x6));
assign Wn48x6 = (~(Dr18x6 & Do48x6));
assign Do48x6 = (Ba38x6 | Lgj7z6[70]);
assign In48x6 = (Iq18x6 | Lgj7z6[70]);
assign Qk48x6 = (~(Fjb7z6[26] & Lriiw6));
assign Cxv7v6 = (~(Ko48x6 & Ro48x6));
assign Ro48x6 = (~(Nxm7x6 & Gydov6));
assign Ko48x6 = (Yo48x6 & Fp48x6);
assign Fp48x6 = (~(Ohj7z6[24] & Mp48x6));
assign Mp48x6 = (~(Tp48x6 & Aq48x6));
assign Aq48x6 = (Hq48x6 & Jn18x6);
assign Hq48x6 = (~(Oq48x6 & Vq48x6));
assign Vq48x6 = (Cr48x6 & Bnx7x6);
assign Cr48x6 = (~(Lgj7z6[74] & Lo18x6));
assign Oq48x6 = (So18x6 & Jr48x6);
assign Jr48x6 = (~(Gp18x6 & Lgj7z6[73]));
assign Tp48x6 = (Qr48x6 & Xr48x6);
assign Xr48x6 = (~(Es48x6 & N0y7x6));
assign Es48x6 = (~(Iq18x6 & Ls48x6));
assign Ls48x6 = (Ba38x6 | Lgj7z6[74]);
assign Qr48x6 = (Dr18x6 | Lgj7z6[74]);
assign Yo48x6 = (~(Fjb7z6[27] & Lriiw6));
assign Vwv7v6 = (~(Ss48x6 & Zs48x6));
assign Zs48x6 = (~(Nxm7x6 & Lxdov6));
assign Ss48x6 = (Gt48x6 & Nt48x6);
assign Nt48x6 = (~(Ohj7z6[25] & Ut48x6));
assign Ut48x6 = (~(Bu48x6 & Iu48x6));
assign Iu48x6 = (Pu48x6 & Jn18x6);
assign Pu48x6 = (~(Wu48x6 & Dv48x6));
assign Dv48x6 = (Kv48x6 & Inx7x6);
assign Kv48x6 = (~(Lgj7z6[77] & Lo18x6));
assign Wu48x6 = (So18x6 & Rv48x6);
assign Rv48x6 = (~(Gp18x6 & Lgj7z6[76]));
assign Bu48x6 = (Yv48x6 & Fw48x6);
assign Fw48x6 = (~(Mw48x6 & Tw48x6));
assign Mw48x6 = (~(Dr18x6 & Ax48x6));
assign Ax48x6 = (Ba38x6 | Lgj7z6[76]);
assign Yv48x6 = (Iq18x6 | Lgj7z6[76]);
assign Gt48x6 = (~(Fjb7z6[28] & Lriiw6));
assign Owv7v6 = (~(Hx48x6 & Ox48x6));
assign Ox48x6 = (~(Nxm7x6 & Exdov6));
assign Hx48x6 = (Vx48x6 & Cy48x6);
assign Cy48x6 = (~(Ohj7z6[26] & Jy48x6));
assign Jy48x6 = (~(Qy48x6 & Xy48x6));
assign Xy48x6 = (Ez48x6 & Jn18x6);
assign Ez48x6 = (~(Lz48x6 & Sz48x6));
assign Sz48x6 = (Zz48x6 & Zzx7x6);
assign Zz48x6 = (~(Lgj7z6[80] & Lo18x6));
assign Lz48x6 = (So18x6 & G058x6);
assign G058x6 = (~(Gp18x6 & Lgj7z6[79]));
assign Qy48x6 = (N058x6 & U058x6);
assign U058x6 = (~(B158x6 & R2y7x6));
assign B158x6 = (~(Iq18x6 & I158x6));
assign I158x6 = (Ba38x6 | Lgj7z6[80]);
assign N058x6 = (Dr18x6 | Lgj7z6[80]);
assign Vx48x6 = (~(Fjb7z6[29] & Lriiw6));
assign Hwv7v6 = (~(P158x6 & W158x6));
assign W158x6 = (~(Nxm7x6 & Vvdov6));
assign P158x6 = (D258x6 & K258x6);
assign K258x6 = (~(Ohj7z6[27] & R258x6));
assign R258x6 = (~(Y258x6 & F358x6));
assign F358x6 = (M358x6 & Jn18x6);
assign M358x6 = (~(T358x6 & A458x6));
assign A458x6 = (H458x6 & Szx7x6);
assign H458x6 = (~(Lgj7z6[83] & Lo18x6));
assign T358x6 = (So18x6 & O458x6);
assign O458x6 = (~(Gp18x6 & Lgj7z6[82]));
assign Y258x6 = (V458x6 & C558x6);
assign C558x6 = (~(J558x6 & Q558x6));
assign J558x6 = (~(Dr18x6 & X558x6));
assign X558x6 = (Ba38x6 | Lgj7z6[82]);
assign V458x6 = (Iq18x6 | Lgj7z6[82]);
assign D258x6 = (~(Fjb7z6[30] & Lriiw6));
assign Awv7v6 = (~(E658x6 & L658x6));
assign L658x6 = (~(Nxm7x6 & Ovdov6));
assign E658x6 = (S658x6 & Z658x6);
assign Z658x6 = (~(Ohj7z6[28] & G758x6));
assign G758x6 = (~(N758x6 & U758x6));
assign U758x6 = (B858x6 & Jn18x6);
assign B858x6 = (~(I858x6 & P858x6));
assign P858x6 = (W858x6 & Crx7x6);
assign Crx7x6 = (!Lgj7z6[84]);
assign W858x6 = (~(Lgj7z6[86] & Lo18x6));
assign I858x6 = (So18x6 & D958x6);
assign D958x6 = (~(Gp18x6 & Lgj7z6[85]));
assign N758x6 = (K958x6 & R958x6);
assign R958x6 = (~(Y958x6 & Fa58x6));
assign Y958x6 = (~(Iq18x6 & Ma58x6));
assign Ma58x6 = (Ba38x6 | Lgj7z6[86]);
assign K958x6 = (Dr18x6 | Lgj7z6[86]);
assign S658x6 = (~(Fjb7z6[31] & Lriiw6));
assign Tvv7v6 = (~(Ta58x6 & Ab58x6));
assign Ab58x6 = (~(Nxm7x6 & Rtdov6));
assign Ta58x6 = (Hb58x6 & Ob58x6);
assign Ob58x6 = (~(Ohj7z6[29] & Vb58x6));
assign Vb58x6 = (~(Cc58x6 & Jc58x6));
assign Jc58x6 = (Qc58x6 & Jn18x6);
assign Qc58x6 = (~(Xc58x6 & Ed58x6));
assign Ed58x6 = (Ld58x6 & Gq6iw6);
assign Ld58x6 = (~(Lgj7z6[89] & Lo18x6));
assign Xc58x6 = (So18x6 & Sd58x6);
assign Sd58x6 = (~(Gp18x6 & Lgj7z6[88]));
assign Cc58x6 = (Zd58x6 & Ge58x6);
assign Ge58x6 = (~(Ne58x6 & T16iw6));
assign Ne58x6 = (~(Dr18x6 & Ue58x6));
assign Ue58x6 = (Ba38x6 | Lgj7z6[88]);
assign Zd58x6 = (Iq18x6 | Lgj7z6[88]);
assign Hb58x6 = (~(Fjb7z6[32] & Lriiw6));
assign Mvv7v6 = (~(Bf58x6 & If58x6));
assign If58x6 = (~(Nxm7x6 & Tudov6));
assign Bf58x6 = (Pf58x6 & Wf58x6);
assign Wf58x6 = (~(Ohj7z6[30] & Dg58x6));
assign Dg58x6 = (~(Kg58x6 & Rg58x6));
assign Rg58x6 = (Yg58x6 & Jn18x6);
assign Yg58x6 = (~(Fh58x6 & Mh58x6));
assign Mh58x6 = (Th58x6 & Xrx7x6);
assign Th58x6 = (~(Lgj7z6[92] & Lo18x6));
assign Fh58x6 = (So18x6 & Ai58x6);
assign Ai58x6 = (~(Gp18x6 & Lgj7z6[91]));
assign Kg58x6 = (Hi58x6 & Oi58x6);
assign Oi58x6 = (~(Vi58x6 & Cj58x6));
assign Vi58x6 = (~(Iq18x6 & Jj58x6));
assign Jj58x6 = (Ba38x6 | Lgj7z6[92]);
assign Hi58x6 = (Dr18x6 | Lgj7z6[92]);
assign Pf58x6 = (~(Fjb7z6[33] & Lriiw6));
assign Fvv7v6 = (~(Qj58x6 & Xj58x6));
assign Xj58x6 = (~(Nxm7x6 & Mudov6));
assign Qj58x6 = (Ek58x6 & Lk58x6);
assign Lk58x6 = (~(Ohj7z6[31] & Sk58x6));
assign Sk58x6 = (~(Zk58x6 & Gl58x6));
assign Gl58x6 = (Nl58x6 & Jn18x6);
assign Nl58x6 = (~(Ul58x6 & Bm58x6));
assign Bm58x6 = (Im58x6 & Esx7x6);
assign Im58x6 = (~(Lgj7z6[95] & Lo18x6));
assign Ul58x6 = (So18x6 & Pm58x6);
assign Pm58x6 = (~(Gp18x6 & Lgj7z6[94]));
assign Zk58x6 = (Wm58x6 & Dn58x6);
assign Dn58x6 = (~(Kn58x6 & Rn58x6));
assign Kn58x6 = (~(Dr18x6 & Yn58x6));
assign Yn58x6 = (Ba38x6 | Lgj7z6[94]);
assign Wm58x6 = (Iq18x6 | Lgj7z6[94]);
assign Ek58x6 = (~(Fjb7z6[34] & Lriiw6));
assign Yuv7v6 = (~(Fo58x6 & Mo58x6));
assign Mo58x6 = (~(Nxm7x6 & Hneov6));
assign Fo58x6 = (To58x6 & Ap58x6);
assign Ap58x6 = (~(Ohj7z6[32] & Hp58x6));
assign Hp58x6 = (~(Op58x6 & Vp58x6));
assign Vp58x6 = (Cq58x6 & Jn18x6);
assign Cq58x6 = (~(Jq58x6 & Qq58x6));
assign Qq58x6 = (Xq58x6 & Ua8iw6);
assign Xq58x6 = (~(Lgj7z6[98] & Lo18x6));
assign Jq58x6 = (So18x6 & Er58x6);
assign Er58x6 = (~(Gp18x6 & Lgj7z6[97]));
assign Op58x6 = (Lr58x6 & Sr58x6);
assign Sr58x6 = (~(Zr58x6 & Ju7iw6));
assign Zr58x6 = (~(Iq18x6 & Gs58x6));
assign Gs58x6 = (Ba38x6 | Lgj7z6[98]);
assign Lr58x6 = (Dr18x6 | Lgj7z6[98]);
assign To58x6 = (~(Fjb7z6[35] & Lriiw6));
assign Ruv7v6 = (~(Ns58x6 & Us58x6));
assign Us58x6 = (~(Nxm7x6 & Sbeov6));
assign Ns58x6 = (Bt58x6 & It58x6);
assign It58x6 = (~(Ohj7z6[33] & Pt58x6));
assign Pt58x6 = (~(Wt58x6 & Du58x6));
assign Du58x6 = (Ku58x6 & Jn18x6);
assign Ku58x6 = (~(Ru58x6 & Yu58x6));
assign Yu58x6 = (Fv58x6 & J0w7x6);
assign Fv58x6 = (~(Lgj7z6[101] & Lo18x6));
assign Ru58x6 = (So18x6 & Mv58x6);
assign Mv58x6 = (~(Gp18x6 & Lgj7z6[100]));
assign Wt58x6 = (Tv58x6 & Aw58x6);
assign Aw58x6 = (~(Hw58x6 & Ow58x6));
assign Hw58x6 = (~(Dr18x6 & Vw58x6));
assign Vw58x6 = (Ba38x6 | Lgj7z6[100]);
assign Tv58x6 = (Iq18x6 | Lgj7z6[100]);
assign Bt58x6 = (~(Fjb7z6[36] & Lriiw6));
assign Kuv7v6 = (~(Cx58x6 & Jx58x6));
assign Jx58x6 = (~(Nxm7x6 & Aneov6));
assign Cx58x6 = (Qx58x6 & Xx58x6);
assign Xx58x6 = (~(Ohj7z6[34] & Ey58x6));
assign Ey58x6 = (~(Ly58x6 & Sy58x6));
assign Sy58x6 = (Zy58x6 & Jn18x6);
assign Zy58x6 = (~(Gz58x6 & Nz58x6));
assign Nz58x6 = (Uz58x6 & Qew7x6);
assign Uz58x6 = (~(Lgj7z6[104] & Lo18x6));
assign Gz58x6 = (So18x6 & B068x6);
assign B068x6 = (~(Gp18x6 & Lgj7z6[103]));
assign Ly58x6 = (I068x6 & P068x6);
assign P068x6 = (~(W068x6 & Bhw7x6));
assign W068x6 = (~(Iq18x6 & D168x6));
assign D168x6 = (Ba38x6 | Lgj7z6[104]);
assign I068x6 = (Dr18x6 | Lgj7z6[104]);
assign Qx58x6 = (~(Fjb7z6[37] & Lriiw6));
assign Duv7v6 = (~(K168x6 & R168x6));
assign R168x6 = (~(Nxm7x6 & Jaeov6));
assign K168x6 = (Y168x6 & F268x6);
assign F268x6 = (~(Ohj7z6[35] & M268x6));
assign M268x6 = (~(T268x6 & A368x6));
assign A368x6 = (H368x6 & Jn18x6);
assign H368x6 = (~(O368x6 & V368x6));
assign V368x6 = (C468x6 & Jew7x6);
assign C468x6 = (~(Lgj7z6[107] & Lo18x6));
assign O368x6 = (So18x6 & J468x6);
assign J468x6 = (~(Gp18x6 & Lgj7z6[106]));
assign T268x6 = (Q468x6 & X468x6);
assign X468x6 = (~(E568x6 & L568x6));
assign E568x6 = (~(Dr18x6 & S568x6));
assign S568x6 = (Ba38x6 | Lgj7z6[106]);
assign Q468x6 = (Iq18x6 | Lgj7z6[106]);
assign Y168x6 = (~(Fjb7z6[38] & Lriiw6));
assign Wtv7v6 = (~(Z568x6 & G668x6));
assign G668x6 = (~(Nxm7x6 & Ujeov6));
assign Z568x6 = (N668x6 & U668x6);
assign U668x6 = (~(Ohj7z6[36] & B768x6));
assign B768x6 = (~(I768x6 & P768x6));
assign P768x6 = (W768x6 & Jn18x6);
assign W768x6 = (~(D868x6 & K868x6));
assign K868x6 = (R868x6 & Q88iw6);
assign R868x6 = (~(Lgj7z6[110] & Lo18x6));
assign D868x6 = (So18x6 & Y868x6);
assign Y868x6 = (~(Gp18x6 & Lgj7z6[109]));
assign I768x6 = (F968x6 & M968x6);
assign M968x6 = (~(T968x6 & Ot7iw6));
assign T968x6 = (~(Iq18x6 & Aa68x6));
assign Aa68x6 = (Ba38x6 | Lgj7z6[110]);
assign F968x6 = (Dr18x6 | Lgj7z6[110]);
assign N668x6 = (~(Fjb7z6[39] & Lriiw6));
assign Ptv7v6 = (~(Ha68x6 & Oa68x6));
assign Oa68x6 = (~(Nxm7x6 & Caeov6));
assign Ha68x6 = (Va68x6 & Cb68x6);
assign Cb68x6 = (~(Ohj7z6[37] & Jb68x6));
assign Jb68x6 = (~(Qb68x6 & Xb68x6));
assign Xb68x6 = (Ec68x6 & Jn18x6);
assign Ec68x6 = (~(Lc68x6 & Sc68x6));
assign Sc68x6 = (Zc68x6 & Myv7x6);
assign Zc68x6 = (~(Lgj7z6[113] & Lo18x6));
assign Lc68x6 = (So18x6 & Gd68x6);
assign Gd68x6 = (~(Gp18x6 & Lgj7z6[112]));
assign Qb68x6 = (Nd68x6 & Ud68x6);
assign Ud68x6 = (~(Be68x6 & V6w7x6));
assign Be68x6 = (~(Dr18x6 & Ie68x6));
assign Ie68x6 = (Ba38x6 | Lgj7z6[112]);
assign Nd68x6 = (Iq18x6 | Lgj7z6[112]);
assign Va68x6 = (~(Fjb7z6[40] & Lriiw6));
assign Itv7v6 = (~(Pe68x6 & We68x6));
assign We68x6 = (~(Nxm7x6 & Njeov6));
assign Pe68x6 = (Df68x6 & Kf68x6);
assign Kf68x6 = (~(Ohj7z6[38] & Rf68x6));
assign Rf68x6 = (~(Yf68x6 & Fg68x6));
assign Fg68x6 = (Mg68x6 & Jn18x6);
assign Mg68x6 = (~(Tg68x6 & Ah68x6));
assign Ah68x6 = (Hh68x6 & T5w7x6);
assign Hh68x6 = (~(Lgj7z6[116] & Lo18x6));
assign Tg68x6 = (So18x6 & Oh68x6);
assign Oh68x6 = (~(Gp18x6 & Lgj7z6[115]));
assign Yf68x6 = (Vh68x6 & Ci68x6);
assign Ci68x6 = (~(Ji68x6 & Qi68x6));
assign Ji68x6 = (~(Iq18x6 & Xi68x6));
assign Xi68x6 = (Ba38x6 | Lgj7z6[116]);
assign Vh68x6 = (Dr18x6 | Lgj7z6[116]);
assign Df68x6 = (~(Fjb7z6[41] & Lriiw6));
assign Btv7v6 = (~(Ej68x6 & Lj68x6));
assign Lj68x6 = (~(Nxm7x6 & F8eov6));
assign Ej68x6 = (Sj68x6 & Zj68x6);
assign Zj68x6 = (~(Ohj7z6[39] & Gk68x6));
assign Gk68x6 = (~(Nk68x6 & Uk68x6));
assign Uk68x6 = (Bl68x6 & Jn18x6);
assign Bl68x6 = (~(Il68x6 & Pl68x6));
assign Pl68x6 = (Wl68x6 & A6w7x6);
assign Wl68x6 = (~(Lgj7z6[119] & Lo18x6));
assign Il68x6 = (So18x6 & Dm68x6);
assign Dm68x6 = (~(Gp18x6 & Lgj7z6[118]));
assign Nk68x6 = (Km68x6 & Rm68x6);
assign Rm68x6 = (~(Ym68x6 & O6w7x6));
assign Ym68x6 = (~(Dr18x6 & Fn68x6));
assign Fn68x6 = (Ba38x6 | Lgj7z6[118]);
assign Km68x6 = (Iq18x6 | Lgj7z6[118]);
assign Sj68x6 = (~(Fjb7z6[42] & Lriiw6));
assign Usv7v6 = (~(Mn68x6 & Tn68x6));
assign Tn68x6 = (~(Nxm7x6 & Grdov6));
assign Mn68x6 = (Ao68x6 & Ho68x6);
assign Ho68x6 = (~(Ohj7z6[40] & Oo68x6));
assign Oo68x6 = (~(Vo68x6 & Cp68x6));
assign Cp68x6 = (Jp68x6 & Jn18x6);
assign Jp68x6 = (~(Qp68x6 & Xp68x6));
assign Xp68x6 = (Eq68x6 & O78iw6);
assign Eq68x6 = (~(Lgj7z6[122] & Lo18x6));
assign Qp68x6 = (So18x6 & Lq68x6);
assign Lq68x6 = (~(Gp18x6 & Lgj7z6[121]));
assign Vo68x6 = (Sq68x6 & Zq68x6);
assign Zq68x6 = (~(Gr68x6 & Ts7iw6));
assign Gr68x6 = (~(Iq18x6 & Nr68x6));
assign Nr68x6 = (Ba38x6 | Lgj7z6[122]);
assign Sq68x6 = (Dr18x6 | Lgj7z6[122]);
assign Ao68x6 = (~(Fjb7z6[43] & Lriiw6));
assign Nsv7v6 = (~(Ur68x6 & Bs68x6));
assign Bs68x6 = (~(Nxm7x6 & Zqdov6));
assign Ur68x6 = (Is68x6 & Ps68x6);
assign Ps68x6 = (~(Ohj7z6[41] & Ws68x6));
assign Ws68x6 = (~(Dt68x6 & Kt68x6));
assign Kt68x6 = (Rt68x6 & Jn18x6);
assign Rt68x6 = (~(Yt68x6 & Fu68x6));
assign Fu68x6 = (Mu68x6 & Rpw7x6);
assign Mu68x6 = (~(Lgj7z6[125] & Lo18x6));
assign Yt68x6 = (So18x6 & Tu68x6);
assign Tu68x6 = (~(Gp18x6 & Lgj7z6[124]));
assign Dt68x6 = (Av68x6 & Hv68x6);
assign Hv68x6 = (~(Ov68x6 & Vv68x6));
assign Ov68x6 = (~(Dr18x6 & Cw68x6));
assign Cw68x6 = (Ba38x6 | Lgj7z6[124]);
assign Av68x6 = (Iq18x6 | Lgj7z6[124]);
assign Is68x6 = (~(Fjb7z6[44] & Lriiw6));
assign Gsv7v6 = (~(Jw68x6 & Qw68x6));
assign Qw68x6 = (~(Nxm7x6 & Eqdov6));
assign Jw68x6 = (Xw68x6 & Ex68x6);
assign Ex68x6 = (~(Ohj7z6[42] & Lx68x6));
assign Lx68x6 = (~(Sx68x6 & Zx68x6));
assign Zx68x6 = (Gy68x6 & Jn18x6);
assign Gy68x6 = (~(Ny68x6 & Uy68x6));
assign Uy68x6 = (Bz68x6 & Y3x7x6);
assign Bz68x6 = (~(Lgj7z6[128] & Lo18x6));
assign Ny68x6 = (So18x6 & Iz68x6);
assign Iz68x6 = (~(Gp18x6 & Lgj7z6[127]));
assign Sx68x6 = (Pz68x6 & Wz68x6);
assign Wz68x6 = (~(D078x6 & J6x7x6));
assign D078x6 = (~(Iq18x6 & K078x6));
assign K078x6 = (Ba38x6 | Lgj7z6[128]);
assign Pz68x6 = (Dr18x6 | Lgj7z6[128]);
assign Xw68x6 = (~(Fjb7z6[45] & Lriiw6));
assign Zrv7v6 = (~(R078x6 & Y078x6));
assign Y078x6 = (~(Nxm7x6 & Xpdov6));
assign R078x6 = (F178x6 & M178x6);
assign M178x6 = (~(Ohj7z6[43] & T178x6));
assign T178x6 = (~(A278x6 & H278x6));
assign H278x6 = (O278x6 & Jn18x6);
assign O278x6 = (~(V278x6 & C378x6));
assign C378x6 = (J378x6 & R3x7x6);
assign J378x6 = (~(Lgj7z6[131] & Lo18x6));
assign V278x6 = (So18x6 & Q378x6);
assign Q378x6 = (~(Gp18x6 & Lgj7z6[130]));
assign A278x6 = (X378x6 & E478x6);
assign E478x6 = (~(L478x6 & S478x6));
assign L478x6 = (~(Dr18x6 & Z478x6));
assign Z478x6 = (Ba38x6 | Lgj7z6[130]);
assign X378x6 = (Iq18x6 | Lgj7z6[130]);
assign F178x6 = (~(Fjb7z6[46] & Lriiw6));
assign Srv7v6 = (~(G578x6 & N578x6));
assign N578x6 = (~(Nxm7x6 & Oodov6));
assign G578x6 = (U578x6 & B678x6);
assign B678x6 = (~(Ohj7z6[44] & I678x6));
assign I678x6 = (~(P678x6 & W678x6));
assign W678x6 = (D778x6 & Jn18x6);
assign D778x6 = (~(K778x6 & R778x6));
assign R778x6 = (Y778x6 & M68iw6);
assign M68iw6 = (!Lgj7z6[132]);
assign Y778x6 = (~(Lgj7z6[134] & Lo18x6));
assign K778x6 = (So18x6 & F878x6);
assign F878x6 = (~(Gp18x6 & Lgj7z6[133]));
assign P678x6 = (M878x6 & T878x6);
assign T878x6 = (~(A978x6 & Yr7iw6));
assign A978x6 = (~(Iq18x6 & H978x6));
assign H978x6 = (Ba38x6 | Lgj7z6[134]);
assign M878x6 = (Dr18x6 | Lgj7z6[134]);
assign U578x6 = (~(Fjb7z6[47] & Lriiw6));
assign Lrv7v6 = (~(O978x6 & V978x6));
assign V978x6 = (~(Nxm7x6 & Hodov6));
assign O978x6 = (Ca78x6 & Ja78x6);
assign Ja78x6 = (~(Ohj7z6[45] & Qa78x6));
assign Qa78x6 = (~(Xa78x6 & Eb78x6));
assign Eb78x6 = (Lb78x6 & Jn18x6);
assign Lb78x6 = (~(Sb78x6 & Zb78x6));
assign Zb78x6 = (Gc78x6 & Ltw7x6);
assign Gc78x6 = (~(Lgj7z6[137] & Lo18x6));
assign Sb78x6 = (So18x6 & Nc78x6);
assign Nc78x6 = (~(Gp18x6 & Lgj7z6[136]));
assign Xa78x6 = (Uc78x6 & Bd78x6);
assign Bd78x6 = (~(Id78x6 & Pvw7x6));
assign Id78x6 = (~(Dr18x6 & Pd78x6));
assign Pd78x6 = (Ba38x6 | Lgj7z6[136]);
assign Uc78x6 = (Iq18x6 | Lgj7z6[136]);
assign Ca78x6 = (~(Fjb7z6[48] & Lriiw6));
assign Erv7v6 = (~(Wd78x6 & De78x6));
assign De78x6 = (~(Nxm7x6 & Kmdov6));
assign Wd78x6 = (Ke78x6 & Re78x6);
assign Re78x6 = (~(Ohj7z6[46] & Ye78x6));
assign Ye78x6 = (~(Ff78x6 & Mf78x6));
assign Mf78x6 = (Tf78x6 & Jn18x6);
assign Tf78x6 = (~(Ag78x6 & Hg78x6));
assign Hg78x6 = (Og78x6 & Guw7x6);
assign Og78x6 = (~(Lgj7z6[140] & Lo18x6));
assign Ag78x6 = (So18x6 & Vg78x6);
assign Vg78x6 = (~(Gp18x6 & Lgj7z6[139]));
assign Ff78x6 = (Ch78x6 & Jh78x6);
assign Jh78x6 = (~(Qh78x6 & Dww7x6));
assign Qh78x6 = (~(Iq18x6 & Xh78x6));
assign Xh78x6 = (Ba38x6 | Lgj7z6[140]);
assign Ch78x6 = (Dr18x6 | Lgj7z6[140]);
assign Ke78x6 = (~(Fjb7z6[49] & Lriiw6));
assign Xqv7v6 = (~(Ei78x6 & Li78x6));
assign Li78x6 = (~(Nxm7x6 & Aueov6));
assign Ei78x6 = (Si78x6 & Zi78x6);
assign Zi78x6 = (~(Ohj7z6[47] & Gj78x6));
assign Gj78x6 = (~(Nj78x6 & Uj78x6));
assign Uj78x6 = (Bk78x6 & Jn18x6);
assign Bk78x6 = (~(Ik78x6 & Pk78x6));
assign Pk78x6 = (Wk78x6 & Nuw7x6);
assign Wk78x6 = (~(Lgj7z6[143] & Lo18x6));
assign Ik78x6 = (So18x6 & Dl78x6);
assign Dl78x6 = (~(Gp18x6 & Lgj7z6[142]));
assign Nj78x6 = (Kl78x6 & Rl78x6);
assign Rl78x6 = (~(Yl78x6 & Uuw7x6));
assign Yl78x6 = (~(Dr18x6 & Fm78x6));
assign Fm78x6 = (Ba38x6 | Lgj7z6[142]);
assign Kl78x6 = (Iq18x6 | Lgj7z6[142]);
assign Si78x6 = (~(Fjb7z6[50] & Lriiw6));
assign Qqv7v6 = (~(Mm78x6 & Tm78x6));
assign Tm78x6 = (~(Nxm7x6 & Sieov6));
assign Mm78x6 = (An78x6 & Hn78x6);
assign Hn78x6 = (~(Ohj7z6[48] & On78x6));
assign On78x6 = (~(Vn78x6 & Co78x6));
assign Co78x6 = (Jo78x6 & Jn18x6);
assign Jo78x6 = (~(Qo78x6 & Xo78x6));
assign Xo78x6 = (Ep78x6 & Xvt7x6);
assign Ep78x6 = (~(Lgj7z6[146] & Lo18x6));
assign Qo78x6 = (So18x6 & Lp78x6);
assign Lp78x6 = (~(Gp18x6 & Lgj7z6[145]));
assign Vn78x6 = (Sp78x6 & Zp78x6);
assign Zp78x6 = (~(Gq78x6 & Wcu7x6));
assign Gq78x6 = (~(Iq18x6 & Nq78x6));
assign Nq78x6 = (Ba38x6 | Lgj7z6[146]);
assign Sp78x6 = (Dr18x6 | Lgj7z6[146]);
assign An78x6 = (~(Fjb7z6[51] & Lriiw6));
assign Jqv7v6 = (~(Uq78x6 & Br78x6));
assign Br78x6 = (~(Nxm7x6 & H9eov6));
assign Uq78x6 = (Ir78x6 & Pr78x6);
assign Pr78x6 = (~(Ohj7z6[49] & Wr78x6));
assign Wr78x6 = (~(Ds78x6 & Ks78x6));
assign Ks78x6 = (Rs78x6 & Jn18x6);
assign Rs78x6 = (~(Ys78x6 & Ft78x6));
assign Ft78x6 = (Mt78x6 & Qvt7x6);
assign Mt78x6 = (~(Lgj7z6[149] & Lo18x6));
assign Ys78x6 = (So18x6 & Tt78x6);
assign Tt78x6 = (~(Gp18x6 & Lgj7z6[148]));
assign Ds78x6 = (Au78x6 & Hu78x6);
assign Hu78x6 = (~(Ou78x6 & Vu78x6));
assign Ou78x6 = (~(Dr18x6 & Cv78x6));
assign Cv78x6 = (Ba38x6 | Lgj7z6[148]);
assign Au78x6 = (Iq18x6 | Lgj7z6[148]);
assign Ir78x6 = (~(Fjb7z6[52] & Lriiw6));
assign Cqv7v6 = (~(Jv78x6 & Qv78x6));
assign Qv78x6 = (~(Nxm7x6 & Lieov6));
assign Jv78x6 = (Xv78x6 & Ew78x6);
assign Ew78x6 = (~(Ohj7z6[50] & Lw78x6));
assign Lw78x6 = (~(Sw78x6 & Zw78x6));
assign Zw78x6 = (Gx78x6 & Jn18x6);
assign Gx78x6 = (~(Nx78x6 & Ux78x6));
assign Ux78x6 = (By78x6 & J9u7x6);
assign By78x6 = (~(Lgj7z6[152] & Lo18x6));
assign Nx78x6 = (So18x6 & Iy78x6);
assign Iy78x6 = (~(Gp18x6 & Lgj7z6[151]));
assign Sw78x6 = (Py78x6 & Wy78x6);
assign Wy78x6 = (~(Dz78x6 & Gbu7x6));
assign Dz78x6 = (~(Iq18x6 & Kz78x6));
assign Kz78x6 = (Ba38x6 | Lgj7z6[152]);
assign Py78x6 = (Dr18x6 | Lgj7z6[152]);
assign Xv78x6 = (~(Fjb7z6[53] & Lriiw6));
assign Vpv7v6 = (~(Rz78x6 & Yz78x6));
assign Yz78x6 = (~(Nxm7x6 & A9eov6));
assign Rz78x6 = (F088x6 & M088x6);
assign M088x6 = (~(Ohj7z6[51] & T088x6));
assign T088x6 = (~(A188x6 & H188x6));
assign H188x6 = (O188x6 & Jn18x6);
assign O188x6 = (~(V188x6 & C288x6));
assign C288x6 = (J288x6 & C9u7x6);
assign J288x6 = (~(Lgj7z6[155] & Lo18x6));
assign V188x6 = (So18x6 & Q288x6);
assign Q288x6 = (~(Gp18x6 & Lgj7z6[154]));
assign A188x6 = (X288x6 & E388x6);
assign E388x6 = (~(L388x6 & S388x6));
assign L388x6 = (~(Dr18x6 & Z388x6));
assign Z388x6 = (Ba38x6 | Lgj7z6[154]);
assign X288x6 = (Iq18x6 | Lgj7z6[154]);
assign F088x6 = (~(Fjb7z6[54] & Lriiw6));
assign Opv7v6 = (~(G488x6 & N488x6));
assign N488x6 = (~(Nxm7x6 & Jidov6));
assign G488x6 = (U488x6 & B588x6);
assign B588x6 = (~(Ohj7z6[52] & I588x6));
assign I588x6 = (~(P588x6 & W588x6));
assign W588x6 = (D688x6 & Jn18x6);
assign D688x6 = (~(K688x6 & R688x6));
assign R688x6 = (Y688x6 & F0u7x6);
assign Y688x6 = (~(Lgj7z6[158] & Lo18x6));
assign K688x6 = (So18x6 & F788x6);
assign F788x6 = (~(Gp18x6 & Lgj7z6[157]));
assign P588x6 = (M788x6 & T788x6);
assign T788x6 = (~(A888x6 & H888x6));
assign A888x6 = (~(Iq18x6 & O888x6));
assign O888x6 = (Ba38x6 | Lgj7z6[158]);
assign M788x6 = (Dr18x6 | Lgj7z6[158]);
assign U488x6 = (~(Fjb7z6[55] & Lriiw6));
assign Hpv7v6 = (~(V888x6 & C988x6));
assign C988x6 = (~(Nxm7x6 & Ljdov6));
assign V888x6 = (J988x6 & Q988x6);
assign Q988x6 = (~(Ohj7z6[53] & X988x6));
assign X988x6 = (~(Ea88x6 & La88x6));
assign La88x6 = (Sa88x6 & Jn18x6);
assign Sa88x6 = (~(Za88x6 & Gb88x6));
assign Gb88x6 = (Nb88x6 & M0u7x6);
assign Nb88x6 = (~(Lgj7z6[161] & Lo18x6));
assign Za88x6 = (So18x6 & Ub88x6);
assign Ub88x6 = (~(Gp18x6 & Lgj7z6[160]));
assign Ea88x6 = (Bc88x6 & Ic88x6);
assign Ic88x6 = (~(Pc88x6 & V1u7x6));
assign Pc88x6 = (~(Dr18x6 & Wc88x6));
assign Wc88x6 = (Ba38x6 | Lgj7z6[160]);
assign Bc88x6 = (Iq18x6 | Lgj7z6[160]);
assign J988x6 = (~(Fjb7z6[56] & Lriiw6));
assign Apv7v6 = (~(Dd88x6 & Kd88x6));
assign Kd88x6 = (~(Nxm7x6 & Ejdov6));
assign Dd88x6 = (Rd88x6 & Yd88x6);
assign Yd88x6 = (~(Ohj7z6[54] & Fe88x6));
assign Fe88x6 = (~(Me88x6 & Te88x6));
assign Te88x6 = (Af88x6 & Jn18x6);
assign Af88x6 = (~(Hf88x6 & Of88x6));
assign Of88x6 = (Vf88x6 & Cg88x6);
assign Vf88x6 = (~(Lgj7z6[164] & Lo18x6));
assign Hf88x6 = (So18x6 & Jg88x6);
assign Jg88x6 = (~(Gp18x6 & Lgj7z6[163]));
assign Me88x6 = (Qg88x6 & Xg88x6);
assign Xg88x6 = (~(Eh88x6 & C2u7x6));
assign Eh88x6 = (~(Iq18x6 & Lh88x6));
assign Lh88x6 = (Ba38x6 | Lgj7z6[164]);
assign Qg88x6 = (Dr18x6 | Lgj7z6[164]);
assign Rd88x6 = (~(Fjb7z6[57] & Lriiw6));
assign Tov7v6 = (~(Sh88x6 & Zh88x6));
assign Zh88x6 = (~(Nxm7x6 & Ahdov6));
assign Sh88x6 = (Gi88x6 & Ni88x6);
assign Ni88x6 = (~(Ohj7z6[55] & Ui88x6));
assign Ui88x6 = (~(Bj88x6 & Ij88x6));
assign Ij88x6 = (Pj88x6 & Jn18x6);
assign Pj88x6 = (~(Wj88x6 & Dk88x6));
assign Dk88x6 = (Kk88x6 & Rk88x6);
assign Kk88x6 = (~(Lgj7z6[167] & Lo18x6));
assign Wj88x6 = (So18x6 & Yk88x6);
assign Yk88x6 = (~(Gp18x6 & Lgj7z6[166]));
assign Bj88x6 = (Fl88x6 & Ml88x6);
assign Ml88x6 = (~(Tl88x6 & Am88x6));
assign Tl88x6 = (~(Dr18x6 & Hm88x6));
assign Hm88x6 = (Ba38x6 | Lgj7z6[166]);
assign Fl88x6 = (Iq18x6 | Lgj7z6[166]);
assign Gi88x6 = (~(Fjb7z6[58] & Lriiw6));
assign Mov7v6 = (~(Om88x6 & Vm88x6));
assign Vm88x6 = (~(Nxm7x6 & Mndov6));
assign Om88x6 = (Cn88x6 & Jn88x6);
assign Jn88x6 = (~(Ohj7z6[56] & Qn88x6));
assign Qn88x6 = (~(Xn88x6 & Eo88x6));
assign Eo88x6 = (Lo88x6 & Jn18x6);
assign Lo88x6 = (~(So88x6 & Zo88x6));
assign Zo88x6 = (Gp88x6 & Cnu7x6);
assign Gp88x6 = (~(Lgj7z6[170] & Lo18x6));
assign So88x6 = (So18x6 & Np88x6);
assign Np88x6 = (~(Gp18x6 & Lgj7z6[169]));
assign Xn88x6 = (Up88x6 & Bq88x6);
assign Bq88x6 = (~(Iq88x6 & Pq88x6));
assign Iq88x6 = (~(Iq18x6 & Wq88x6));
assign Wq88x6 = (Ba38x6 | Lgj7z6[170]);
assign Up88x6 = (Dr18x6 | Lgj7z6[170]);
assign Cn88x6 = (~(Fjb7z6[59] & Lriiw6));
assign Fov7v6 = (~(Dr88x6 & Kr88x6));
assign Kr88x6 = (~(Nxm7x6 & Fndov6));
assign Dr88x6 = (Rr88x6 & Yr88x6);
assign Yr88x6 = (~(Ohj7z6[57] & Fs88x6));
assign Fs88x6 = (~(Ms88x6 & Ts88x6));
assign Ts88x6 = (At88x6 & Jn18x6);
assign At88x6 = (~(Ht88x6 & Ot88x6));
assign Ot88x6 = (Vt88x6 & Vmu7x6);
assign Vt88x6 = (~(Lgj7z6[173] & Lo18x6));
assign Ht88x6 = (So18x6 & Cu88x6);
assign Cu88x6 = (~(Gp18x6 & Lgj7z6[172]));
assign Ms88x6 = (Ju88x6 & Qu88x6);
assign Qu88x6 = (~(Xu88x6 & J1v7x6));
assign Xu88x6 = (~(Dr18x6 & Ev88x6));
assign Ev88x6 = (Ba38x6 | Lgj7z6[172]);
assign Ju88x6 = (Iq18x6 | Lgj7z6[172]);
assign Rr88x6 = (~(Fjb7z6[60] & Lriiw6));
assign Ynv7v6 = (~(Lv88x6 & Sv88x6));
assign Sv88x6 = (~(Nxm7x6 & Nkdov6));
assign Lv88x6 = (Zv88x6 & Gw88x6);
assign Gw88x6 = (~(Ohj7z6[58] & Nw88x6));
assign Nw88x6 = (~(Uw88x6 & Bx88x6));
assign Bx88x6 = (Ix88x6 & Jn18x6);
assign Ix88x6 = (~(Px88x6 & Wx88x6));
assign Wx88x6 = (Dy88x6 & A0v7x6);
assign Dy88x6 = (~(Lgj7z6[176] & Lo18x6));
assign Px88x6 = (So18x6 & Ky88x6);
assign Ky88x6 = (~(Gp18x6 & Lgj7z6[175]));
assign Uw88x6 = (Ry88x6 & Yy88x6);
assign Yy88x6 = (~(Fz88x6 & Mz88x6));
assign Fz88x6 = (~(Iq18x6 & Tz88x6));
assign Tz88x6 = (Ba38x6 | Lgj7z6[176]);
assign Ry88x6 = (Dr18x6 | Lgj7z6[176]);
assign Zv88x6 = (~(Fjb7z6[61] & Lriiw6));
assign Rnv7v6 = (~(A098x6 & H098x6));
assign H098x6 = (~(Nxm7x6 & Gkdov6));
assign A098x6 = (O098x6 & V098x6);
assign V098x6 = (~(Ohj7z6[59] & C198x6));
assign C198x6 = (~(J198x6 & Q198x6));
assign Q198x6 = (X198x6 & Jn18x6);
assign X198x6 = (~(E298x6 & L298x6));
assign L298x6 = (S298x6 & H0v7x6);
assign S298x6 = (~(Lgj7z6[179] & Lo18x6));
assign E298x6 = (So18x6 & Z298x6);
assign Z298x6 = (~(Gp18x6 & Lgj7z6[178]));
assign J198x6 = (G398x6 & N398x6);
assign N398x6 = (~(U398x6 & O0v7x6));
assign U398x6 = (~(Dr18x6 & B498x6));
assign B498x6 = (Ba38x6 | Lgj7z6[178]);
assign G398x6 = (Iq18x6 | Lgj7z6[178]);
assign O098x6 = (~(Fjb7z6[62] & Lriiw6));
assign Knv7v6 = (~(I498x6 & P498x6));
assign P498x6 = (~(Nxm7x6 & Tgdov6));
assign I498x6 = (W498x6 & D598x6);
assign D598x6 = (~(Ohj7z6[60] & K598x6));
assign K598x6 = (~(R598x6 & Y598x6));
assign Y598x6 = (F698x6 & Jn18x6);
assign F698x6 = (~(M698x6 & T698x6));
assign T698x6 = (A798x6 & H798x6);
assign A798x6 = (~(Lgj7z6[182] & Lo18x6));
assign M698x6 = (So18x6 & O798x6);
assign O798x6 = (~(Gp18x6 & Lgj7z6[181]));
assign R598x6 = (V798x6 & C898x6);
assign C898x6 = (~(J898x6 & Q898x6));
assign J898x6 = (~(Iq18x6 & X898x6));
assign X898x6 = (Ba38x6 | Lgj7z6[182]);
assign V798x6 = (Dr18x6 | Lgj7z6[182]);
assign W498x6 = (~(Fjb7z6[63] & Lriiw6));
assign Dnv7v6 = (~(E998x6 & L998x6));
assign L998x6 = (~(Nxm7x6 & Wedov6));
assign E998x6 = (S998x6 & Z998x6);
assign Z998x6 = (~(Ohj7z6[61] & Ga98x6));
assign Ga98x6 = (~(Na98x6 & Ua98x6));
assign Ua98x6 = (Bb98x6 & Jn18x6);
assign Bb98x6 = (~(Ib98x6 & Pb98x6));
assign Pb98x6 = (Wb98x6 & Dc98x6);
assign Wb98x6 = (~(Lgj7z6[185] & Lo18x6));
assign Ib98x6 = (So18x6 & Kc98x6);
assign Kc98x6 = (~(Gp18x6 & Lgj7z6[184]));
assign So18x6 = (Rc98x6 & Yc98x6);
assign Na98x6 = (Fd98x6 & Md98x6);
assign Md98x6 = (~(Td98x6 & Ae98x6));
assign Td98x6 = (~(Dr18x6 & He98x6));
assign He98x6 = (Ba38x6 | Lgj7z6[184]);
assign Fd98x6 = (Iq18x6 | Lgj7z6[184]);
assign S998x6 = (~(Fjb7z6[64] & Lriiw6));
assign Wmv7v6 = (~(Oe98x6 & Ve98x6));
assign Ve98x6 = (~(Nxm7x6 & Rfdov6));
assign Oe98x6 = (Cf98x6 & Jf98x6);
assign Jf98x6 = (~(Ohj7z6[62] & Qf98x6));
assign Qf98x6 = (~(Xf98x6 & Eg98x6));
assign Eg98x6 = (Lg98x6 & Jn18x6);
assign Lg98x6 = (~(Sg98x6 & Zg98x6));
assign Sg98x6 = (~(Iq18x6 & Gh98x6));
assign Gh98x6 = (Ba38x6 | Lgj7z6[188]);
assign Xf98x6 = (Nh98x6 & Uh98x6);
assign Uh98x6 = (Dr18x6 | Lgj7z6[188]);
assign Nh98x6 = (~(Bi98x6 & Ii98x6));
assign Ii98x6 = (Pi98x6 & Yru7x6);
assign Pi98x6 = (~(Wi98x6 & Lo18x6));
assign Wi98x6 = (~(Rc98x6 & Dj98x6));
assign Bi98x6 = (Yc98x6 & Kj98x6);
assign Kj98x6 = (~(Gp18x6 & Lgj7z6[187]));
assign Cf98x6 = (~(Fjb7z6[65] & Lriiw6));
assign Pmv7v6 = (~(Rj98x6 & Yj98x6));
assign Yj98x6 = (~(Nxm7x6 & Sweov6));
assign Nxm7x6 = (Fk98x6 & Sriiw6);
assign Fk98x6 = (Zriiw6 & L2cet6);
assign Rj98x6 = (Mk98x6 & Tk98x6);
assign Tk98x6 = (~(Ohj7z6[63] & Al98x6));
assign Al98x6 = (~(Hl98x6 & Ol98x6));
assign Ol98x6 = (Vl98x6 & Jn18x6);
assign Jn18x6 = (~(Cm98x6 & Yc98x6));
assign Cm98x6 = (Jm98x6 & Qm98x6);
assign Qm98x6 = (~(Za2nv6 & Pym7x6));
assign Vl98x6 = (~(Xm98x6 & En98x6));
assign Xm98x6 = (~(Dr18x6 & Ln98x6));
assign Ln98x6 = (Ba38x6 | Lgj7z6[190]);
assign Ba38x6 = (!Wq18x6);
assign Dr18x6 = (Sn98x6 | Zn98x6);
assign Hl98x6 = (Go98x6 & No98x6);
assign No98x6 = (Iq18x6 | Lgj7z6[190]);
assign Iq18x6 = (~(Wq18x6 & Uo98x6));
assign Wq18x6 = (~(Zn98x6 | Bp98x6));
assign Zn98x6 = (!Yc98x6);
assign Go98x6 = (~(Ip98x6 & Pp98x6));
assign Pp98x6 = (Wp98x6 & Rru7x6);
assign Wp98x6 = (~(Dq98x6 & Lo18x6));
assign Lo18x6 = (~(Rc98x6 & Uo98x6));
assign Uo98x6 = (~(H1m8v6 & Sn98x6));
assign Sn98x6 = (~(Kq98x6 & H1m8v6));
assign Kq98x6 = (Pym7x6 ? CURRPRI[7] : Ppb7z6[7]);
assign Dq98x6 = (~(Rc98x6 & En98x6));
assign Rc98x6 = (Rq98x6 & Rwl8v6);
assign Rq98x6 = (Pym7x6 ? CURRPRI[5] : Ppb7z6[5]);
assign Pym7x6 = (!Dk18x6);
assign Ip98x6 = (Yc98x6 & Yq98x6);
assign Yq98x6 = (~(Gp18x6 & Lgj7z6[190]));
assign Gp18x6 = (Bp98x6 & Zyl8v6);
assign Bp98x6 = (Dk18x6 ? Fr98x6 : Bfr7x6);
assign Dk18x6 = (Sugov6 & Ea2nv6);
assign Fr98x6 = (~(Zyl8v6 & Ppb7z6[6]));
assign Yc98x6 = (Mr98x6 & Sriiw6);
assign Sriiw6 = (!Gsiiw6);
assign Mr98x6 = (Kk18x6 & Tr98x6);
assign Tr98x6 = (~(As98x6 & Zriiw6));
assign As98x6 = (~(Hs98x6 | L2cet6));
assign Kk18x6 = (~(Inadt6 & Offov6));
assign Offov6 = (~(Os98x6 & Sugov6));
assign Os98x6 = (Inadt6 & Vs98x6);
assign Mk98x6 = (~(Fjb7z6[66] & Lriiw6));
assign Lriiw6 = (Gsiiw6 & Usiiw6);
assign Usiiw6 = (!M6bdt6);
assign Gsiiw6 = (~(Ct98x6 & Dzeov6));
assign Dzeov6 = (Hcget6 & U3cet6);
assign Ct98x6 = (Jd47v6 & Jt98x6);
assign Jt98x6 = (!Byeov6);
assign Byeov6 = (~(Qt98x6 & Pyeov6));
assign Qt98x6 = (~(Lunov6 & Sunov6));
assign Lunov6 = (Xt98x6 & Eu98x6);
assign Imv7v6 = (~(Lu98x6 & Su98x6));
assign Su98x6 = (~(L8wnv6 & Itb7z6[26]));
assign Lu98x6 = (Zu98x6 & Gv98x6);
assign Gv98x6 = (~(G9wnv6 & Nv98x6));
assign Nv98x6 = (~(Uv98x6 & Bw98x6));
assign Bw98x6 = (Iw98x6 & Pw98x6);
assign Pw98x6 = (Wawnv6 | Ww98x6);
assign Iw98x6 = (~(Dtm7z6[3] & Dx98x6));
assign Uv98x6 = (Kx98x6 & Rx98x6);
assign Rx98x6 = (~(Dtm7z6[0] & HRDATAD[26]));
assign Kx98x6 = (~(Dtm7z6[1] & HRDATAS[26]));
assign Zu98x6 = (~(Fcwnv6 & Voyhw6));
assign Voyhw6 = (JTAGNSW ? Aixmz6[26] : Ulxmz6[26]);
assign Bmv7v6 = (K94iw6 ? Mi5ft6 : Yx98x6);
assign Ulv7v6 = (~(Fy98x6 & My98x6));
assign My98x6 = (Ty98x6 & Az98x6);
assign Ty98x6 = (~(X9fov6 | Xle8v6));
assign Xle8v6 = (Hz98x6 & Oz98x6);
assign Oz98x6 = (V0fiw6 & Vz98x6);
assign Hz98x6 = (Hyp7z6[3] & HTMDHBURST[0]);
assign Fy98x6 = (C0a8x6 & U0r7x6);
assign C0a8x6 = (~(Eo2ft6 & J0a8x6));
assign J0a8x6 = (~(Na9ov6 & Q0a8x6));
assign Nlv7v6 = (~(X0a8x6 & E1a8x6));
assign E1a8x6 = (L1a8x6 & S1a8x6);
assign L1a8x6 = (~(Eafov6 | Yfw7v6));
assign Yfw7v6 = (Z1a8x6 & G2a8x6);
assign G2a8x6 = (~(N2a8x6 | Hmp7z6[2]));
assign Z1a8x6 = (Hmp7z6[3] & HTMDHBURST[0]);
assign X0a8x6 = (U2a8x6 & B3a8x6);
assign B3a8x6 = (~(Fk2ft6 & I3a8x6));
assign I3a8x6 = (~(Na9ov6 & P3a8x6));
assign Na9ov6 = (Aj4ft6 & M297z6);
assign U2a8x6 = (~(M55ft6 & Bb9ov6));
assign Glv7v6 = (~(W3a8x6 & D4a8x6));
assign D4a8x6 = (~(K4a8x6 & Xy5ft6));
assign Zkv7v6 = (~(R4a8x6 & Y4a8x6));
assign Y4a8x6 = (~(F5a8x6 & Q8o7x6));
assign F5a8x6 = (~(Az98x6 & M5a8x6));
assign M5a8x6 = (~(T5a8x6 & S1a8x6));
assign R4a8x6 = (~(Jhr7z6[0] & K4a8x6));
assign Skv7v6 = (T5a8x6 ? A6a8x6 : Jhr7z6[1]);
assign A6a8x6 = (Q8o7x6 & Az98x6);
assign Lkv7v6 = (~(H6a8x6 & O6a8x6));
assign O6a8x6 = (~(V6a8x6 & U42nv6));
assign H6a8x6 = (Pdq7z6[0] ? J7a8x6 : C7a8x6);
assign Ekv7v6 = (~(Q7a8x6 & X7a8x6));
assign X7a8x6 = (~(V6a8x6 & B52nv6));
assign Q7a8x6 = (Pdq7z6[1] ? L8a8x6 : E8a8x6);
assign E8a8x6 = (~(S8a8x6 & Pdq7z6[0]));
assign Xjv7v6 = (~(Z8a8x6 & G9a8x6));
assign G9a8x6 = (~(V6a8x6 & I52nv6));
assign Z8a8x6 = (Pdq7z6[2] ? U9a8x6 : N9a8x6);
assign U9a8x6 = (L8a8x6 & Baa8x6);
assign Baa8x6 = (C7a8x6 | Pdq7z6[1]);
assign L8a8x6 = (J7a8x6 & Iaa8x6);
assign Iaa8x6 = (C7a8x6 | Pdq7z6[0]);
assign N9a8x6 = (~(Paa8x6 & S8a8x6));
assign Qjv7v6 = (~(Waa8x6 & Dba8x6));
assign Dba8x6 = (~(V6a8x6 & P52nv6));
assign Waa8x6 = (Pdq7z6[3] ? Rba8x6 : Kba8x6);
assign Kba8x6 = (~(Yba8x6 & S8a8x6));
assign Jjv7v6 = (~(Fca8x6 & Mca8x6));
assign Mca8x6 = (~(V6a8x6 & W52nv6));
assign Fca8x6 = (Pdq7z6[4] ? Ada8x6 : Tca8x6);
assign Ada8x6 = (Rba8x6 & Hda8x6);
assign Hda8x6 = (C7a8x6 | Pdq7z6[3]);
assign Rba8x6 = (J7a8x6 & Oda8x6);
assign Oda8x6 = (C7a8x6 | Yba8x6);
assign Tca8x6 = (~(Vda8x6 & Yba8x6));
assign Vda8x6 = (S8a8x6 & Pdq7z6[3]);
assign Cjv7v6 = (~(Cea8x6 & Jea8x6));
assign Jea8x6 = (~(V6a8x6 & D62nv6));
assign Cea8x6 = (Pdq7z6[5] ? Xea8x6 : Qea8x6);
assign Qea8x6 = (~(Efa8x6 & S8a8x6));
assign Viv7v6 = (~(Lfa8x6 & Sfa8x6));
assign Sfa8x6 = (~(V6a8x6 & K62nv6));
assign Lfa8x6 = (Pdq7z6[6] ? Gga8x6 : Zfa8x6);
assign Oiv7v6 = (~(Nga8x6 & Uga8x6));
assign Uga8x6 = (~(V6a8x6 & R62nv6));
assign Nga8x6 = (Pdq7z6[7] ? Iha8x6 : Bha8x6);
assign Iha8x6 = (Gga8x6 & Pha8x6);
assign Pha8x6 = (~(S8a8x6 & Wha8x6));
assign Gga8x6 = (Xea8x6 & Dia8x6);
assign Dia8x6 = (C7a8x6 | Pdq7z6[5]);
assign Xea8x6 = (J7a8x6 & Kia8x6);
assign Kia8x6 = (C7a8x6 | Efa8x6);
assign J7a8x6 = (!Ria8x6);
assign Bha8x6 = (Zfa8x6 | Wha8x6);
assign Wha8x6 = (!Pdq7z6[6]);
assign Zfa8x6 = (~(Yia8x6 & Efa8x6));
assign Yia8x6 = (S8a8x6 & Pdq7z6[5]);
assign S8a8x6 = (!C7a8x6);
assign C7a8x6 = (Fja8x6 | Ria8x6);
assign Ria8x6 = (~(Fja8x6 | Mja8x6));
assign Fja8x6 = (V6a8x6 | Tja8x6);
assign Tja8x6 = (Aka8x6 & Etgiw6);
assign Aka8x6 = (~(Hka8x6 | Kxfiw6));
assign V6a8x6 = (Jsgiw6 & Oka8x6);
assign Hiv7v6 = (~(Vka8x6 & Cla8x6));
assign Cla8x6 = (~(Jla8x6 & U42nv6));
assign Vka8x6 = (Cjq7z6[0] ? Xla8x6 : Qla8x6);
assign Aiv7v6 = (~(Ema8x6 & Lma8x6));
assign Lma8x6 = (~(Jla8x6 & B52nv6));
assign Ema8x6 = (Cjq7z6[1] ? Zma8x6 : Sma8x6);
assign Sma8x6 = (~(Gna8x6 & Cjq7z6[0]));
assign Thv7v6 = (~(Nna8x6 & Una8x6));
assign Una8x6 = (~(Jla8x6 & I52nv6));
assign Nna8x6 = (Cjq7z6[2] ? Ioa8x6 : Boa8x6);
assign Ioa8x6 = (Zma8x6 & Poa8x6);
assign Poa8x6 = (Qla8x6 | Cjq7z6[1]);
assign Zma8x6 = (Xla8x6 & Woa8x6);
assign Woa8x6 = (Qla8x6 | Cjq7z6[0]);
assign Boa8x6 = (~(Dpa8x6 & Gna8x6));
assign Mhv7v6 = (~(Kpa8x6 & Rpa8x6));
assign Rpa8x6 = (~(Jla8x6 & P52nv6));
assign Kpa8x6 = (Cjq7z6[3] ? Fqa8x6 : Ypa8x6);
assign Ypa8x6 = (~(Mqa8x6 & Gna8x6));
assign Fhv7v6 = (~(Tqa8x6 & Ara8x6));
assign Ara8x6 = (~(Jla8x6 & W52nv6));
assign Tqa8x6 = (Cjq7z6[4] ? Ora8x6 : Hra8x6);
assign Ora8x6 = (Fqa8x6 & Vra8x6);
assign Vra8x6 = (Qla8x6 | Cjq7z6[3]);
assign Fqa8x6 = (Xla8x6 & Csa8x6);
assign Csa8x6 = (Qla8x6 | Mqa8x6);
assign Hra8x6 = (~(Jsa8x6 & Mqa8x6));
assign Jsa8x6 = (Gna8x6 & Cjq7z6[3]);
assign Ygv7v6 = (~(Qsa8x6 & Xsa8x6));
assign Xsa8x6 = (~(Jla8x6 & D62nv6));
assign Qsa8x6 = (Cjq7z6[5] ? Lta8x6 : Eta8x6);
assign Eta8x6 = (~(Sta8x6 & Gna8x6));
assign Rgv7v6 = (~(Zta8x6 & Gua8x6));
assign Gua8x6 = (~(Jla8x6 & K62nv6));
assign Zta8x6 = (Cjq7z6[6] ? Uua8x6 : Nua8x6);
assign Kgv7v6 = (~(Bva8x6 & Iva8x6));
assign Iva8x6 = (~(Jla8x6 & R62nv6));
assign Bva8x6 = (Cjq7z6[7] ? Wva8x6 : Pva8x6);
assign Wva8x6 = (Uua8x6 & Dwa8x6);
assign Dwa8x6 = (~(Gna8x6 & Kwa8x6));
assign Uua8x6 = (Lta8x6 & Rwa8x6);
assign Rwa8x6 = (Qla8x6 | Cjq7z6[5]);
assign Lta8x6 = (Xla8x6 & Ywa8x6);
assign Ywa8x6 = (Qla8x6 | Sta8x6);
assign Xla8x6 = (!Fxa8x6);
assign Pva8x6 = (Nua8x6 | Kwa8x6);
assign Kwa8x6 = (!Cjq7z6[6]);
assign Nua8x6 = (~(Mxa8x6 & Sta8x6));
assign Mxa8x6 = (Gna8x6 & Cjq7z6[5]);
assign Gna8x6 = (!Qla8x6);
assign Qla8x6 = (Txa8x6 | Fxa8x6);
assign Fxa8x6 = (~(Txa8x6 | Aya8x6));
assign Txa8x6 = (Jla8x6 | Hya8x6);
assign Hya8x6 = (Oya8x6 & Etgiw6);
assign Oya8x6 = (~(Vya8x6 | Oyhov6));
assign Jla8x6 = (Jsgiw6 & Cza8x6);
assign Dgv7v6 = (~(Jza8x6 & Qza8x6));
assign Qza8x6 = (~(Gqr7z6[1] & Inhiw6));
assign Jza8x6 = (Xza8x6 & E0b8x6);
assign E0b8x6 = (~(L0b8x6 & Aw77z6));
assign Xza8x6 = (~(Rzr7z6[1] & S0b8x6));
assign Wfv7v6 = (~(Z0b8x6 & G1b8x6));
assign G1b8x6 = (~(Gqr7z6[2] & Inhiw6));
assign Z0b8x6 = (N1b8x6 & U1b8x6);
assign U1b8x6 = (~(L0b8x6 & Sv77z6));
assign N1b8x6 = (~(Rzr7z6[2] & S0b8x6));
assign Pfv7v6 = (~(B2b8x6 & I2b8x6));
assign I2b8x6 = (~(Gqr7z6[3] & Inhiw6));
assign B2b8x6 = (P2b8x6 & W2b8x6);
assign W2b8x6 = (~(L0b8x6 & Kv77z6));
assign P2b8x6 = (~(Rzr7z6[3] & S0b8x6));
assign Ifv7v6 = (~(D3b8x6 & K3b8x6));
assign K3b8x6 = (~(Gqr7z6[4] & Inhiw6));
assign D3b8x6 = (R3b8x6 & Y3b8x6);
assign Y3b8x6 = (~(L0b8x6 & Cv77z6));
assign R3b8x6 = (~(Rzr7z6[4] & S0b8x6));
assign Bfv7v6 = (~(F4b8x6 & M4b8x6));
assign M4b8x6 = (~(Gqr7z6[5] & Inhiw6));
assign F4b8x6 = (T4b8x6 & A5b8x6);
assign A5b8x6 = (~(L0b8x6 & Uu77z6));
assign T4b8x6 = (~(Rzr7z6[5] & S0b8x6));
assign Uev7v6 = (~(H5b8x6 & O5b8x6));
assign O5b8x6 = (~(Gqr7z6[6] & Inhiw6));
assign H5b8x6 = (V5b8x6 & C6b8x6);
assign C6b8x6 = (~(L0b8x6 & Mu77z6));
assign V5b8x6 = (~(Rzr7z6[6] & S0b8x6));
assign Nev7v6 = (~(J6b8x6 & Q6b8x6));
assign Q6b8x6 = (~(Gqr7z6[7] & Inhiw6));
assign J6b8x6 = (X6b8x6 & E7b8x6);
assign E7b8x6 = (~(L0b8x6 & Eu77z6));
assign X6b8x6 = (~(Rzr7z6[7] & S0b8x6));
assign Gev7v6 = (~(L7b8x6 & S7b8x6));
assign S7b8x6 = (~(Gqr7z6[8] & Inhiw6));
assign L7b8x6 = (Z7b8x6 & G8b8x6);
assign G8b8x6 = (~(L0b8x6 & Wt77z6));
assign Z7b8x6 = (~(Rzr7z6[8] & S0b8x6));
assign Zdv7v6 = (~(N8b8x6 & U8b8x6));
assign U8b8x6 = (~(Gqr7z6[9] & Inhiw6));
assign N8b8x6 = (B9b8x6 & I9b8x6);
assign I9b8x6 = (~(L0b8x6 & Ot77z6));
assign B9b8x6 = (~(Rzr7z6[9] & S0b8x6));
assign Sdv7v6 = (~(P9b8x6 & W9b8x6));
assign W9b8x6 = (~(Gqr7z6[10] & Inhiw6));
assign P9b8x6 = (Dab8x6 & Kab8x6);
assign Kab8x6 = (~(L0b8x6 & Gt77z6));
assign Dab8x6 = (~(Rzr7z6[10] & S0b8x6));
assign Ldv7v6 = (~(Rab8x6 & Yab8x6));
assign Yab8x6 = (~(Gqr7z6[11] & Inhiw6));
assign Rab8x6 = (Fbb8x6 & Mbb8x6);
assign Mbb8x6 = (~(L0b8x6 & Ys77z6));
assign Fbb8x6 = (~(Rzr7z6[11] & S0b8x6));
assign Edv7v6 = (~(Tbb8x6 & Acb8x6));
assign Acb8x6 = (~(Gqr7z6[12] & Inhiw6));
assign Tbb8x6 = (Hcb8x6 & Ocb8x6);
assign Ocb8x6 = (~(L0b8x6 & Qs77z6));
assign Hcb8x6 = (~(Rzr7z6[12] & S0b8x6));
assign Xcv7v6 = (~(Vcb8x6 & Cdb8x6));
assign Cdb8x6 = (~(Gqr7z6[13] & Inhiw6));
assign Vcb8x6 = (Jdb8x6 & Qdb8x6);
assign Qdb8x6 = (~(L0b8x6 & Is77z6));
assign Jdb8x6 = (~(Rzr7z6[13] & S0b8x6));
assign Qcv7v6 = (~(Xdb8x6 & Eeb8x6));
assign Eeb8x6 = (~(Gqr7z6[14] & Inhiw6));
assign Xdb8x6 = (Leb8x6 & Seb8x6);
assign Seb8x6 = (~(L0b8x6 & As77z6));
assign Leb8x6 = (~(Rzr7z6[14] & S0b8x6));
assign Jcv7v6 = (~(Zeb8x6 & Gfb8x6));
assign Gfb8x6 = (~(Gqr7z6[15] & Inhiw6));
assign Zeb8x6 = (Nfb8x6 & Ufb8x6);
assign Ufb8x6 = (~(L0b8x6 & Sr77z6));
assign Nfb8x6 = (~(Rzr7z6[15] & S0b8x6));
assign Ccv7v6 = (~(Bgb8x6 & Igb8x6));
assign Igb8x6 = (~(Gqr7z6[16] & Inhiw6));
assign Bgb8x6 = (Pgb8x6 & Wgb8x6);
assign Wgb8x6 = (~(L0b8x6 & Kr77z6));
assign Pgb8x6 = (~(Rzr7z6[16] & S0b8x6));
assign Vbv7v6 = (~(Dhb8x6 & Khb8x6));
assign Khb8x6 = (~(Gqr7z6[17] & Inhiw6));
assign Dhb8x6 = (Rhb8x6 & Yhb8x6);
assign Yhb8x6 = (~(L0b8x6 & Cr77z6));
assign Rhb8x6 = (~(Rzr7z6[17] & S0b8x6));
assign Obv7v6 = (~(Fib8x6 & Mib8x6));
assign Mib8x6 = (~(Gqr7z6[18] & Inhiw6));
assign Fib8x6 = (Tib8x6 & Ajb8x6);
assign Ajb8x6 = (~(L0b8x6 & Uq77z6));
assign Tib8x6 = (~(Rzr7z6[18] & S0b8x6));
assign Hbv7v6 = (~(Hjb8x6 & Ojb8x6));
assign Ojb8x6 = (~(Gqr7z6[19] & Inhiw6));
assign Hjb8x6 = (Vjb8x6 & Ckb8x6);
assign Ckb8x6 = (~(L0b8x6 & Mq77z6));
assign Vjb8x6 = (~(Rzr7z6[19] & S0b8x6));
assign Abv7v6 = (~(Jkb8x6 & Qkb8x6));
assign Qkb8x6 = (~(Gqr7z6[20] & Inhiw6));
assign Jkb8x6 = (Xkb8x6 & Elb8x6);
assign Elb8x6 = (~(L0b8x6 & Eq77z6));
assign Xkb8x6 = (~(Rzr7z6[20] & S0b8x6));
assign Tav7v6 = (~(Llb8x6 & Slb8x6));
assign Slb8x6 = (~(Gqr7z6[21] & Inhiw6));
assign Llb8x6 = (Zlb8x6 & Gmb8x6);
assign Gmb8x6 = (~(L0b8x6 & Wp77z6));
assign Zlb8x6 = (~(Rzr7z6[21] & S0b8x6));
assign Mav7v6 = (~(Nmb8x6 & Umb8x6));
assign Umb8x6 = (~(Gqr7z6[22] & Inhiw6));
assign Nmb8x6 = (Bnb8x6 & Inb8x6);
assign Inb8x6 = (~(L0b8x6 & Op77z6));
assign Bnb8x6 = (~(Rzr7z6[22] & S0b8x6));
assign Fav7v6 = (~(Pnb8x6 & Wnb8x6));
assign Wnb8x6 = (~(Gqr7z6[23] & Inhiw6));
assign Pnb8x6 = (Dob8x6 & Kob8x6);
assign Kob8x6 = (~(L0b8x6 & Gp77z6));
assign Dob8x6 = (~(Rzr7z6[23] & S0b8x6));
assign Y9v7v6 = (~(Rob8x6 & Yob8x6));
assign Yob8x6 = (~(Gqr7z6[24] & Inhiw6));
assign Rob8x6 = (Fpb8x6 & Mpb8x6);
assign Mpb8x6 = (~(L0b8x6 & Yo77z6));
assign Fpb8x6 = (~(Rzr7z6[24] & S0b8x6));
assign R9v7v6 = (~(Tpb8x6 & Aqb8x6));
assign Aqb8x6 = (~(Gqr7z6[25] & Inhiw6));
assign Tpb8x6 = (Hqb8x6 & Oqb8x6);
assign Oqb8x6 = (~(L0b8x6 & Qo77z6));
assign Hqb8x6 = (~(Rzr7z6[25] & S0b8x6));
assign K9v7v6 = (~(Vqb8x6 & Crb8x6));
assign Crb8x6 = (~(Gqr7z6[26] & Inhiw6));
assign Vqb8x6 = (Jrb8x6 & Qrb8x6);
assign Qrb8x6 = (~(L0b8x6 & Io77z6));
assign Jrb8x6 = (~(Rzr7z6[26] & S0b8x6));
assign D9v7v6 = (~(Xrb8x6 & Esb8x6));
assign Esb8x6 = (~(Gqr7z6[27] & Inhiw6));
assign Xrb8x6 = (Lsb8x6 & Ssb8x6);
assign Ssb8x6 = (~(L0b8x6 & Ao77z6));
assign Lsb8x6 = (~(Rzr7z6[27] & S0b8x6));
assign W8v7v6 = (~(Zsb8x6 & Gtb8x6));
assign Gtb8x6 = (~(Gqr7z6[28] & Inhiw6));
assign Zsb8x6 = (Ntb8x6 & Utb8x6);
assign Utb8x6 = (~(L0b8x6 & Sn77z6));
assign Ntb8x6 = (~(Rzr7z6[28] & S0b8x6));
assign P8v7v6 = (~(Bub8x6 & Iub8x6));
assign Iub8x6 = (~(Gqr7z6[29] & Inhiw6));
assign Bub8x6 = (Pub8x6 & Wub8x6);
assign Wub8x6 = (~(L0b8x6 & Kn77z6));
assign Pub8x6 = (~(Rzr7z6[29] & S0b8x6));
assign I8v7v6 = (~(Dvb8x6 & Kvb8x6));
assign Kvb8x6 = (~(Gqr7z6[30] & Inhiw6));
assign Dvb8x6 = (Rvb8x6 & Yvb8x6);
assign Yvb8x6 = (~(L0b8x6 & Cn77z6));
assign Rvb8x6 = (~(Rzr7z6[30] & S0b8x6));
assign B8v7v6 = (~(Fwb8x6 & Mwb8x6));
assign Mwb8x6 = (~(Gqr7z6[31] & Inhiw6));
assign Fwb8x6 = (Twb8x6 & Axb8x6);
assign Axb8x6 = (~(L0b8x6 & Um77z6));
assign L0b8x6 = (~(Inhiw6 | Wfo7v6));
assign Twb8x6 = (~(Rzr7z6[31] & S0b8x6));
assign S0b8x6 = (~(Inhiw6 | Wdtnv6));
assign U7v7v6 = (~(Hxb8x6 & Oxb8x6));
assign Oxb8x6 = (~(Z3gnv6 & Vxb8x6));
assign Z3gnv6 = (HTMDHBURST[0] & Cmm7z6[0]);
assign Hxb8x6 = (~(Cor7z6[0] & K4a8x6));
assign N7v7v6 = (~(Cyb8x6 & Jyb8x6));
assign Jyb8x6 = (Qyb8x6 & Xyb8x6);
assign Xyb8x6 = (~(Gxfnv6 & Vxb8x6));
assign Gxfnv6 = (HTMDHBURST[0] & Cmm7z6[1]);
assign Qyb8x6 = (~(Ezb8x6 & Aw77z6));
assign Cyb8x6 = (Lzb8x6 & Szb8x6);
assign Szb8x6 = (~(Zzb8x6 & Rzr7z6[1]));
assign Lzb8x6 = (~(Cor7z6[1] & K4a8x6));
assign G7v7v6 = (~(G0c8x6 & N0c8x6));
assign N0c8x6 = (U0c8x6 & B1c8x6);
assign B1c8x6 = (~(Qvfnv6 & Vxb8x6));
assign Qvfnv6 = (~(I1c8x6 | Kygnv6));
assign U0c8x6 = (~(Ezb8x6 & Sv77z6));
assign G0c8x6 = (P1c8x6 & W1c8x6);
assign W1c8x6 = (~(Zzb8x6 & Rzr7z6[2]));
assign P1c8x6 = (~(Cor7z6[2] & K4a8x6));
assign Z6v7v6 = (~(D2c8x6 & K2c8x6));
assign K2c8x6 = (R2c8x6 & Y2c8x6);
assign Y2c8x6 = (~(Jvfnv6 & Vxb8x6));
assign Jvfnv6 = (~(F3c8x6 | Kygnv6));
assign F3c8x6 = (!Cmm7z6[3]);
assign R2c8x6 = (~(Ezb8x6 & Kv77z6));
assign D2c8x6 = (M3c8x6 & T3c8x6);
assign T3c8x6 = (~(Zzb8x6 & Rzr7z6[3]));
assign M3c8x6 = (~(Cor7z6[3] & K4a8x6));
assign S6v7v6 = (~(A4c8x6 & H4c8x6));
assign H4c8x6 = (O4c8x6 & V4c8x6);
assign V4c8x6 = (~(Hufnv6 & Vxb8x6));
assign Hufnv6 = (~(C5c8x6 | Kygnv6));
assign C5c8x6 = (!Cmm7z6[4]);
assign O4c8x6 = (~(Ezb8x6 & Cv77z6));
assign A4c8x6 = (J5c8x6 & Q5c8x6);
assign Q5c8x6 = (~(Zzb8x6 & Rzr7z6[4]));
assign J5c8x6 = (~(Cor7z6[4] & K4a8x6));
assign L6v7v6 = (~(X5c8x6 & E6c8x6));
assign E6c8x6 = (L6c8x6 & S6c8x6);
assign S6c8x6 = (~(Ttfnv6 & Vxb8x6));
assign Ttfnv6 = (~(Z6c8x6 | Kygnv6));
assign Z6c8x6 = (!Cmm7z6[5]);
assign L6c8x6 = (~(Ezb8x6 & Uu77z6));
assign X5c8x6 = (G7c8x6 & N7c8x6);
assign N7c8x6 = (~(Zzb8x6 & Rzr7z6[5]));
assign G7c8x6 = (~(Cor7z6[5] & K4a8x6));
assign E6v7v6 = (~(U7c8x6 & B8c8x6));
assign B8c8x6 = (I8c8x6 & P8c8x6);
assign P8c8x6 = (~(Ysfnv6 & Vxb8x6));
assign Ysfnv6 = (~(Kygnv6 | W8c8x6));
assign W8c8x6 = (!Cmm7z6[6]);
assign I8c8x6 = (~(Ezb8x6 & Mu77z6));
assign U7c8x6 = (D9c8x6 & K9c8x6);
assign K9c8x6 = (~(Zzb8x6 & Rzr7z6[6]));
assign D9c8x6 = (~(Cor7z6[6] & K4a8x6));
assign X5v7v6 = (~(R9c8x6 & Y9c8x6));
assign Y9c8x6 = (Fac8x6 & Mac8x6);
assign Mac8x6 = (~(Rsfnv6 & Vxb8x6));
assign Rsfnv6 = (~(Kygnv6 | Tac8x6));
assign Tac8x6 = (!Cmm7z6[7]);
assign Fac8x6 = (~(Ezb8x6 & Eu77z6));
assign R9c8x6 = (Abc8x6 & Hbc8x6);
assign Hbc8x6 = (~(Zzb8x6 & Rzr7z6[7]));
assign Abc8x6 = (~(K4a8x6 & Cor7z6[7]));
assign Q5v7v6 = (~(Obc8x6 & Vbc8x6));
assign Vbc8x6 = (Ccc8x6 & Jcc8x6);
assign Jcc8x6 = (~(Ksfnv6 & Vxb8x6));
assign Ksfnv6 = (~(Kygnv6 | Qcc8x6));
assign Qcc8x6 = (!Cmm7z6[8]);
assign Ccc8x6 = (~(Ezb8x6 & Wt77z6));
assign Obc8x6 = (Xcc8x6 & Edc8x6);
assign Edc8x6 = (~(Zzb8x6 & Rzr7z6[8]));
assign Xcc8x6 = (~(Cor7z6[8] & K4a8x6));
assign J5v7v6 = (~(Ldc8x6 & Sdc8x6));
assign Sdc8x6 = (Zdc8x6 & Gec8x6);
assign Gec8x6 = (~(Dsfnv6 & Vxb8x6));
assign Dsfnv6 = (~(Kygnv6 | Nec8x6));
assign Nec8x6 = (!Cmm7z6[9]);
assign Zdc8x6 = (~(Ezb8x6 & Ot77z6));
assign Ldc8x6 = (Uec8x6 & Bfc8x6);
assign Bfc8x6 = (~(Zzb8x6 & Rzr7z6[9]));
assign Uec8x6 = (~(Cor7z6[9] & K4a8x6));
assign C5v7v6 = (~(Ifc8x6 & Pfc8x6));
assign Pfc8x6 = (Wfc8x6 & Dgc8x6);
assign Dgc8x6 = (~(Wyfnv6 & Vxb8x6));
assign Wyfnv6 = (~(Kygnv6 | Kgc8x6));
assign Kgc8x6 = (!Cmm7z6[10]);
assign Wfc8x6 = (~(Ezb8x6 & Gt77z6));
assign Ifc8x6 = (Rgc8x6 & Ygc8x6);
assign Ygc8x6 = (~(Zzb8x6 & Rzr7z6[10]));
assign Rgc8x6 = (~(Cor7z6[10] & K4a8x6));
assign V4v7v6 = (~(Fhc8x6 & Mhc8x6));
assign Mhc8x6 = (Thc8x6 & Aic8x6);
assign Aic8x6 = (~(Pyfnv6 & Vxb8x6));
assign Pyfnv6 = (~(Kygnv6 | Hic8x6));
assign Hic8x6 = (!Cmm7z6[11]);
assign Thc8x6 = (~(Ezb8x6 & Ys77z6));
assign Fhc8x6 = (Oic8x6 & Vic8x6);
assign Vic8x6 = (~(Zzb8x6 & Rzr7z6[11]));
assign Oic8x6 = (~(Cor7z6[11] & K4a8x6));
assign O4v7v6 = (~(Cjc8x6 & Jjc8x6));
assign Jjc8x6 = (Qjc8x6 & Xjc8x6);
assign Xjc8x6 = (~(Byfnv6 & Vxb8x6));
assign Byfnv6 = (~(Kygnv6 | Ekc8x6));
assign Ekc8x6 = (!Cmm7z6[12]);
assign Qjc8x6 = (~(Ezb8x6 & Qs77z6));
assign Cjc8x6 = (Lkc8x6 & Skc8x6);
assign Skc8x6 = (~(Zzb8x6 & Rzr7z6[12]));
assign Lkc8x6 = (~(Cor7z6[12] & K4a8x6));
assign H4v7v6 = (~(Zkc8x6 & Glc8x6));
assign Glc8x6 = (Nlc8x6 & Ulc8x6);
assign Ulc8x6 = (~(Uxfnv6 & Vxb8x6));
assign Uxfnv6 = (~(Kygnv6 | Bmc8x6));
assign Bmc8x6 = (!Cmm7z6[13]);
assign Nlc8x6 = (~(Ezb8x6 & Is77z6));
assign Zkc8x6 = (Imc8x6 & Pmc8x6);
assign Pmc8x6 = (~(Zzb8x6 & Rzr7z6[13]));
assign Imc8x6 = (~(Cor7z6[13] & K4a8x6));
assign A4v7v6 = (~(Wmc8x6 & Dnc8x6));
assign Dnc8x6 = (Knc8x6 & Rnc8x6);
assign Rnc8x6 = (~(Nxfnv6 & Vxb8x6));
assign Nxfnv6 = (~(Kygnv6 | Ync8x6));
assign Ync8x6 = (!Cmm7z6[14]);
assign Knc8x6 = (~(Ezb8x6 & As77z6));
assign Wmc8x6 = (Foc8x6 & Moc8x6);
assign Moc8x6 = (~(Zzb8x6 & Rzr7z6[14]));
assign Foc8x6 = (~(Cor7z6[14] & K4a8x6));
assign T3v7v6 = (~(Toc8x6 & Apc8x6));
assign Apc8x6 = (Hpc8x6 & Opc8x6);
assign Opc8x6 = (~(Ezb8x6 & Sr77z6));
assign Hpc8x6 = (~(Zzb8x6 & Rzr7z6[15]));
assign Toc8x6 = (Vpc8x6 & Cqc8x6);
assign Cqc8x6 = (~(Tp5ft6 & Vxb8x6));
assign Tp5ft6 = (~(Kygnv6 | Jqc8x6));
assign Jqc8x6 = (!Cmm7z6[15]);
assign Vpc8x6 = (~(K4a8x6 & Cor7z6[15]));
assign M3v7v6 = (~(Qqc8x6 & Xqc8x6));
assign Xqc8x6 = (~(Cor7z6[16] & K4a8x6));
assign Qqc8x6 = (Erc8x6 & Lrc8x6);
assign Lrc8x6 = (~(Ezb8x6 & Kr77z6));
assign Erc8x6 = (~(Zzb8x6 & Rzr7z6[16]));
assign F3v7v6 = (~(Src8x6 & Zrc8x6));
assign Zrc8x6 = (~(Cor7z6[17] & K4a8x6));
assign Src8x6 = (Gsc8x6 & Nsc8x6);
assign Nsc8x6 = (~(Ezb8x6 & Cr77z6));
assign Gsc8x6 = (~(Zzb8x6 & Rzr7z6[17]));
assign Y2v7v6 = (~(Usc8x6 & Btc8x6));
assign Btc8x6 = (~(Cor7z6[18] & K4a8x6));
assign Usc8x6 = (Itc8x6 & Ptc8x6);
assign Ptc8x6 = (~(Ezb8x6 & Uq77z6));
assign Itc8x6 = (~(Zzb8x6 & Rzr7z6[18]));
assign R2v7v6 = (~(Wtc8x6 & Duc8x6));
assign Duc8x6 = (~(Cor7z6[19] & K4a8x6));
assign Wtc8x6 = (Kuc8x6 & Ruc8x6);
assign Ruc8x6 = (~(Ezb8x6 & Mq77z6));
assign Kuc8x6 = (~(Zzb8x6 & Rzr7z6[19]));
assign K2v7v6 = (~(Yuc8x6 & Fvc8x6));
assign Fvc8x6 = (~(Cor7z6[20] & K4a8x6));
assign Yuc8x6 = (Mvc8x6 & Tvc8x6);
assign Tvc8x6 = (~(Ezb8x6 & Eq77z6));
assign Mvc8x6 = (~(Zzb8x6 & Rzr7z6[20]));
assign D2v7v6 = (~(Awc8x6 & Hwc8x6));
assign Hwc8x6 = (~(Cor7z6[21] & K4a8x6));
assign Awc8x6 = (Owc8x6 & Vwc8x6);
assign Vwc8x6 = (~(Ezb8x6 & Wp77z6));
assign Owc8x6 = (~(Zzb8x6 & Rzr7z6[21]));
assign W1v7v6 = (~(Cxc8x6 & Jxc8x6));
assign Jxc8x6 = (~(Cor7z6[22] & K4a8x6));
assign Cxc8x6 = (Qxc8x6 & Xxc8x6);
assign Xxc8x6 = (~(Ezb8x6 & Op77z6));
assign Qxc8x6 = (~(Zzb8x6 & Rzr7z6[22]));
assign P1v7v6 = (~(Eyc8x6 & Lyc8x6));
assign Lyc8x6 = (~(K4a8x6 & Cor7z6[23]));
assign Eyc8x6 = (Syc8x6 & Zyc8x6);
assign Zyc8x6 = (~(Ezb8x6 & Gp77z6));
assign Syc8x6 = (~(Zzb8x6 & Rzr7z6[23]));
assign I1v7v6 = (~(Gzc8x6 & Nzc8x6));
assign Nzc8x6 = (~(Cor7z6[24] & K4a8x6));
assign Gzc8x6 = (Uzc8x6 & B0d8x6);
assign B0d8x6 = (~(Ezb8x6 & Yo77z6));
assign Uzc8x6 = (~(Zzb8x6 & Rzr7z6[24]));
assign B1v7v6 = (~(I0d8x6 & P0d8x6));
assign P0d8x6 = (~(Cor7z6[25] & K4a8x6));
assign I0d8x6 = (W0d8x6 & D1d8x6);
assign D1d8x6 = (~(Ezb8x6 & Qo77z6));
assign W0d8x6 = (~(Zzb8x6 & Rzr7z6[25]));
assign U0v7v6 = (~(K1d8x6 & R1d8x6));
assign R1d8x6 = (~(Cor7z6[26] & K4a8x6));
assign K1d8x6 = (Y1d8x6 & F2d8x6);
assign F2d8x6 = (~(Ezb8x6 & Io77z6));
assign Y1d8x6 = (~(Zzb8x6 & Rzr7z6[26]));
assign N0v7v6 = (~(M2d8x6 & T2d8x6));
assign T2d8x6 = (~(Cor7z6[27] & K4a8x6));
assign M2d8x6 = (A3d8x6 & H3d8x6);
assign H3d8x6 = (~(Ezb8x6 & Ao77z6));
assign A3d8x6 = (~(Zzb8x6 & Rzr7z6[27]));
assign G0v7v6 = (~(O3d8x6 & V3d8x6));
assign V3d8x6 = (~(Cor7z6[28] & K4a8x6));
assign O3d8x6 = (C4d8x6 & J4d8x6);
assign J4d8x6 = (~(Ezb8x6 & Sn77z6));
assign C4d8x6 = (~(Zzb8x6 & Rzr7z6[28]));
assign Zzu7v6 = (~(Q4d8x6 & X4d8x6));
assign X4d8x6 = (~(Cor7z6[29] & K4a8x6));
assign Q4d8x6 = (E5d8x6 & L5d8x6);
assign L5d8x6 = (~(Ezb8x6 & Kn77z6));
assign E5d8x6 = (~(Zzb8x6 & Rzr7z6[29]));
assign Szu7v6 = (~(S5d8x6 & Z5d8x6));
assign Z5d8x6 = (~(Cor7z6[30] & K4a8x6));
assign S5d8x6 = (G6d8x6 & N6d8x6);
assign N6d8x6 = (~(Ezb8x6 & Cn77z6));
assign G6d8x6 = (~(Zzb8x6 & Rzr7z6[30]));
assign Lzu7v6 = (~(U6d8x6 & B7d8x6));
assign B7d8x6 = (~(K4a8x6 & Cor7z6[31]));
assign U6d8x6 = (I7d8x6 & P7d8x6);
assign P7d8x6 = (~(Ezb8x6 & Um77z6));
assign Ezb8x6 = (W7d8x6 & W3a8x6);
assign W7d8x6 = (T5a8x6 & Wdtnv6);
assign I7d8x6 = (~(Zzb8x6 & Rzr7z6[31]));
assign Zzb8x6 = (D8d8x6 & W3a8x6);
assign W3a8x6 = (!Vxb8x6);
assign Vxb8x6 = (Q8o7x6 ? K8d8x6 : M12ft6);
assign K8d8x6 = (Az98x6 ? R8d8x6 : Gs2ft6);
assign R8d8x6 = (S1a8x6 ? Y8d8x6 : Dm2ft6);
assign Y8d8x6 = (~(E99ov6 | A0fiw6));
assign A0fiw6 = (!Ei2ft6);
assign D8d8x6 = (Wfo7v6 & T5a8x6);
assign Ezu7v6 = (!F9d8x6);
assign F9d8x6 = (E1b7x6 ? M9d8x6 : I1wiw6);
assign E1b7x6 = (!Jgliw6);
assign M9d8x6 = (~(Qmbet6 & Wfo7v6));
assign Xyu7v6 = (T9d8x6 & Jgliw6);
assign T9d8x6 = (Had8x6 ? Aad8x6 : A0vnv6);
assign Aad8x6 = (~(Oad8x6 & Vad8x6));
assign Oad8x6 = (Cbd8x6 & Qv0ov6);
assign Cbd8x6 = (~(Jbd8x6 & Kvbov6));
assign A0vnv6 = (!O197z6);
assign Qyu7v6 = (Had8x6 ? Qbd8x6 : Qobet6);
assign Had8x6 = (Xbd8x6 | Ecd8x6);
assign Ecd8x6 = (Phhov6 ? Tlmov6 : Lcd8x6);
assign Lcd8x6 = (Rihov6 & Wdtnv6);
assign Xbd8x6 = (T7mov6 | Teliw6);
assign T7mov6 = (Tlmov6 & Ierov6);
assign Qbd8x6 = (Scd8x6 & Jgliw6);
assign Scd8x6 = (~(Vad8x6 & Rihov6));
assign Vad8x6 = (~(Phhov6 | Teliw6));
assign Jyu7v6 = (Ie77v6 & Zcd8x6);
assign Zcd8x6 = (!Wy67v6);
assign Cyu7v6 = (!Gdd8x6);
assign Gdd8x6 = (At67v6 ? Ndd8x6 : Jjrnv6);
assign Ndd8x6 = (Udd8x6 ? Orhov6 : Y097z6);
assign Udd8x6 = (Bed8x6 & Ied8x6);
assign Vxu7v6 = (Ped8x6 & Y9rnv6);
assign Ped8x6 = (Bj77v6 | Nernv6);
assign Oxu7v6 = (~(Wed8x6 & Dfd8x6));
assign Dfd8x6 = (~(Jdymz6[1] & Kfd8x6));
assign Kfd8x6 = (Rfd8x6 | L19iw6);
assign Wed8x6 = (~(Yfd8x6 & B52nv6));
assign Hxu7v6 = (~(Fgd8x6 & Mgd8x6));
assign Mgd8x6 = (~(Jdymz6[0] & Tgd8x6));
assign Tgd8x6 = (Rfd8x6 | Orhov6);
assign Fgd8x6 = (~(Yfd8x6 & U42nv6));
assign Axu7v6 = (~(Ahd8x6 & Hhd8x6));
assign Hhd8x6 = (~(Jdymz6[2] & Ohd8x6));
assign Ohd8x6 = (Rfd8x6 | Fhrnv6);
assign Fhrnv6 = (!I52nv6);
assign Ahd8x6 = (~(Yfd8x6 & I52nv6));
assign Twu7v6 = (~(Vhd8x6 & Cid8x6));
assign Cid8x6 = (~(Jdymz6[3] & Jid8x6));
assign Jid8x6 = (Rfd8x6 | Pohov6);
assign Vhd8x6 = (~(Yfd8x6 & P52nv6));
assign Yfd8x6 = (~(Qid8x6 | Rfd8x6));
assign Rfd8x6 = (~(Xid8x6 & Ejd8x6));
assign Ejd8x6 = (Ljd8x6 | Sjd8x6);
assign Mwu7v6 = (Mi77z6 & Jgliw6);
assign Fwu7v6 = (Pyeov6 ? Zriiw6 : Zjd8x6);
assign Pyeov6 = (~(Gkd8x6 & Nkd8x6));
assign Nkd8x6 = (Ukd8x6 & Bld8x6);
assign Bld8x6 = (~(Zjd8x6 & Ild8x6));
assign Ukd8x6 = (~(R7fet6 & Qubet6));
assign Gkd8x6 = (Pld8x6 & Eu98x6);
assign Eu98x6 = (Wld8x6 | Sh2nv6);
assign Wld8x6 = (!Aiadt6);
assign Pld8x6 = (Wyeov6 ? Kmd8x6 : Dmd8x6);
assign Wyeov6 = (!Y3fet6);
assign Kmd8x6 = (Rmd8x6 & Ymd8x6);
assign Ymd8x6 = (~(Fnd8x6 & Zriiw6));
assign Fnd8x6 = (~(Ild8x6 | T5fet6));
assign Rmd8x6 = (Xt98x6 | Qubet6);
assign Xt98x6 = (~(Qyddt6 & Mnd8x6));
assign Dmd8x6 = (Ldh7v6 & Flg7x6);
assign Zriiw6 = (!Sunov6);
assign Zjd8x6 = (!Ic77z6);
assign Yvu7v6 = (Tnd8x6 ? T5fet6 : Sunov6);
assign Tnd8x6 = (Aod8x6 & Sunov6);
assign Aod8x6 = (~(Ic77z6 & Hod8x6));
assign Hod8x6 = (~(Ood8x6 & Vod8x6));
assign Vod8x6 = (Ga3nv6 & Flg7x6);
assign Flg7x6 = (!Opeet6);
assign Ood8x6 = (~(Ild8x6 | Sugov6));
assign Sugov6 = (!Sh2nv6);
assign Sh2nv6 = (~(Cpd8x6 & Eyknv6));
assign Cpd8x6 = (O5a7z6 & M6a7x6);
assign Ild8x6 = (~(Jpd8x6 & Qpd8x6));
assign Qpd8x6 = (~(TXEV | Ei77z6));
assign Jpd8x6 = (Xpd8x6 & Eqd8x6);
assign Eqd8x6 = (~(RXEV & Lqd8x6));
assign Lqd8x6 = (!Fjb7z6[0]);
assign Xpd8x6 = (~(Itbet6 & L2cet6));
assign Sunov6 = (~(M0edt6 & Mnd8x6));
assign Mnd8x6 = (~(Sqd8x6 | Bklhw6));
assign Sqd8x6 = (~(Mrnov6 & C0wnv6));
assign Rvu7v6 = (~(Zqd8x6 & Grd8x6));
assign Grd8x6 = (~(Ruymz6[15] & Nrd8x6));
assign Zqd8x6 = (Urd8x6 & Bsd8x6);
assign Bsd8x6 = (~(Isd8x6 & Biymz6[15]));
assign Urd8x6 = (~(Ctymz6[15] & Psd8x6));
assign Kvu7v6 = (~(Wsd8x6 & Dtd8x6));
assign Dtd8x6 = (~(Ruymz6[0] & Nrd8x6));
assign Wsd8x6 = (Ktd8x6 & Rtd8x6);
assign Rtd8x6 = (~(Isd8x6 & Biymz6[0]));
assign Ktd8x6 = (~(Ctymz6[0] & Psd8x6));
assign Dvu7v6 = (~(Ytd8x6 & Fud8x6));
assign Fud8x6 = (~(Ruymz6[1] & Nrd8x6));
assign Ytd8x6 = (Mud8x6 & Tud8x6);
assign Tud8x6 = (~(Isd8x6 & Biymz6[1]));
assign Mud8x6 = (~(Ctymz6[1] & Psd8x6));
assign Wuu7v6 = (~(Avd8x6 & Hvd8x6));
assign Hvd8x6 = (~(Ruymz6[2] & Nrd8x6));
assign Avd8x6 = (Ovd8x6 & Vvd8x6);
assign Vvd8x6 = (~(Isd8x6 & Biymz6[2]));
assign Ovd8x6 = (~(Ctymz6[2] & Psd8x6));
assign Puu7v6 = (~(Cwd8x6 & Jwd8x6));
assign Jwd8x6 = (~(Ruymz6[3] & Nrd8x6));
assign Cwd8x6 = (Qwd8x6 & Xwd8x6);
assign Xwd8x6 = (~(Isd8x6 & Biymz6[3]));
assign Qwd8x6 = (~(Ctymz6[3] & Psd8x6));
assign Iuu7v6 = (~(Exd8x6 & Lxd8x6));
assign Lxd8x6 = (~(Ruymz6[4] & Nrd8x6));
assign Exd8x6 = (Sxd8x6 & Zxd8x6);
assign Zxd8x6 = (~(Isd8x6 & Biymz6[4]));
assign Sxd8x6 = (~(Ctymz6[4] & Psd8x6));
assign Buu7v6 = (~(Gyd8x6 & Nyd8x6));
assign Nyd8x6 = (~(Ruymz6[5] & Nrd8x6));
assign Gyd8x6 = (Uyd8x6 & Bzd8x6);
assign Bzd8x6 = (~(Isd8x6 & Biymz6[5]));
assign Uyd8x6 = (~(Ctymz6[5] & Psd8x6));
assign Utu7v6 = (~(Izd8x6 & Pzd8x6));
assign Pzd8x6 = (~(Ruymz6[6] & Nrd8x6));
assign Izd8x6 = (Wzd8x6 & D0e8x6);
assign D0e8x6 = (~(Isd8x6 & Biymz6[6]));
assign Wzd8x6 = (~(Ctymz6[6] & Psd8x6));
assign Ntu7v6 = (~(K0e8x6 & R0e8x6));
assign R0e8x6 = (~(Ruymz6[7] & Nrd8x6));
assign K0e8x6 = (Y0e8x6 & F1e8x6);
assign F1e8x6 = (~(Isd8x6 & Biymz6[7]));
assign Y0e8x6 = (~(Ctymz6[7] & Psd8x6));
assign Gtu7v6 = (~(M1e8x6 & T1e8x6));
assign T1e8x6 = (~(Ruymz6[8] & Nrd8x6));
assign M1e8x6 = (A2e8x6 & H2e8x6);
assign H2e8x6 = (~(Isd8x6 & Biymz6[8]));
assign A2e8x6 = (~(Ctymz6[8] & Psd8x6));
assign Zsu7v6 = (~(O2e8x6 & V2e8x6));
assign V2e8x6 = (~(Ruymz6[9] & Nrd8x6));
assign O2e8x6 = (C3e8x6 & J3e8x6);
assign J3e8x6 = (~(Isd8x6 & Biymz6[9]));
assign C3e8x6 = (~(Ctymz6[9] & Psd8x6));
assign Ssu7v6 = (~(Q3e8x6 & X3e8x6));
assign X3e8x6 = (~(Ruymz6[10] & Nrd8x6));
assign Q3e8x6 = (E4e8x6 & L4e8x6);
assign L4e8x6 = (~(Isd8x6 & Biymz6[10]));
assign E4e8x6 = (~(Ctymz6[10] & Psd8x6));
assign Lsu7v6 = (~(S4e8x6 & Z4e8x6));
assign Z4e8x6 = (~(Ruymz6[11] & Nrd8x6));
assign S4e8x6 = (G5e8x6 & N5e8x6);
assign N5e8x6 = (~(Isd8x6 & Biymz6[11]));
assign G5e8x6 = (~(Ctymz6[11] & Psd8x6));
assign Esu7v6 = (~(U5e8x6 & B6e8x6));
assign B6e8x6 = (~(Ruymz6[12] & Nrd8x6));
assign U5e8x6 = (I6e8x6 & P6e8x6);
assign P6e8x6 = (~(Isd8x6 & Biymz6[12]));
assign I6e8x6 = (~(Ctymz6[12] & Psd8x6));
assign Xru7v6 = (~(W6e8x6 & D7e8x6));
assign D7e8x6 = (~(Ruymz6[13] & Nrd8x6));
assign W6e8x6 = (K7e8x6 & R7e8x6);
assign R7e8x6 = (~(Isd8x6 & Biymz6[13]));
assign K7e8x6 = (~(Ctymz6[13] & Psd8x6));
assign Qru7v6 = (~(Y7e8x6 & F8e8x6));
assign F8e8x6 = (~(Ruymz6[14] & Nrd8x6));
assign Y7e8x6 = (M8e8x6 & T8e8x6);
assign T8e8x6 = (~(Isd8x6 & Biymz6[14]));
assign Isd8x6 = (A9e8x6 & I7dov6);
assign A9e8x6 = (Uh77v6 | Gernv6);
assign M8e8x6 = (~(Ctymz6[14] & Psd8x6));
assign Psd8x6 = (H9e8x6 & I7dov6);
assign I7dov6 = (!Nrd8x6);
assign Nrd8x6 = (~(P7snv6 | Gernv6));
assign H9e8x6 = (~(Gernv6 | Uh77v6));
assign Jru7v6 = (Gecov6 ? O9e8x6 : Ka87v6);
assign Cru7v6 = (Gecov6 ? V9e8x6 : Gnzmz6[39]);
assign Vqu7v6 = (Gecov6 ? Cae8x6 : Gnzmz6[31]);
assign Oqu7v6 = (Gecov6 ? Jae8x6 : Gnzmz6[23]);
assign Hqu7v6 = (Gecov6 ? Wfcov6 : Gnzmz6[15]);
assign Gecov6 = (~(I0snv6 & R1snv6));
assign Wfcov6 = (~(Qae8x6 & Xae8x6));
assign Xae8x6 = (Ebe8x6 & Lbe8x6);
assign Lbe8x6 = (Sbe8x6 & Zbe8x6);
assign Zbe8x6 = (~(TSVALUEB[19] ^ Gnzmz6[21]));
assign Sbe8x6 = (~(Jae8x6 | Gce8x6));
assign Gce8x6 = (Gnzmz6[15] & I0snv6);
assign Jae8x6 = (~(Nce8x6 & Uce8x6));
assign Uce8x6 = (Bde8x6 & Ide8x6);
assign Ide8x6 = (Pde8x6 & Wde8x6);
assign Wde8x6 = (~(TSVALUEB[26] ^ Gnzmz6[29]));
assign Pde8x6 = (~(Cae8x6 | Dee8x6));
assign Dee8x6 = (Gnzmz6[23] & I0snv6);
assign Cae8x6 = (~(Kee8x6 & Ree8x6));
assign Ree8x6 = (Yee8x6 & Ffe8x6);
assign Ffe8x6 = (Mfe8x6 & Tfe8x6);
assign Tfe8x6 = (~(TSVALUEB[33] ^ Gnzmz6[37]));
assign Mfe8x6 = (~(V9e8x6 | Age8x6));
assign Age8x6 = (Gnzmz6[31] & I0snv6);
assign V9e8x6 = (~(Hge8x6 & Oge8x6));
assign Oge8x6 = (Vge8x6 & Che8x6);
assign Che8x6 = (Jhe8x6 & Qhe8x6);
assign Qhe8x6 = (~(TSVALUEB[40] ^ Gnzmz6[45]));
assign Jhe8x6 = (~(O9e8x6 | Xhe8x6));
assign Xhe8x6 = (Gnzmz6[39] & I0snv6);
assign O9e8x6 = (~(Eie8x6 & Lie8x6));
assign Lie8x6 = (Sie8x6 & Zie8x6);
assign Zie8x6 = (~(Gje8x6 | Jc87v6));
assign Jc87v6 = (Xz67v6 & Nje8x6);
assign Nje8x6 = (~(Uje8x6 & F2snv6));
assign F2snv6 = (Uzrnv6 & Bke8x6);
assign Uje8x6 = (Ike8x6 & Y9rnv6);
assign Ike8x6 = (~(L587v6 & I0snv6));
assign Gje8x6 = (Ka87v6 & I0snv6);
assign Sie8x6 = (Pke8x6 & Qg3xx6);
assign Qg3xx6 = (~(TSVALUEB[46] ^ Emc7v6));
assign Pke8x6 = (~(TSVALUEB[44] ^ Qic7v6));
assign Eie8x6 = (Xg3xx6 & Eh3xx6);
assign Eh3xx6 = (Lh3xx6 & Sh3xx6);
assign Sh3xx6 = (~(TSVALUEB[42] ^ Cfc7v6));
assign Lh3xx6 = (~(TSVALUEB[43] ^ Wgc7v6));
assign Xg3xx6 = (Zh3xx6 & Gi3xx6);
assign Gi3xx6 = (~(TSVALUEB[47] ^ Ync7v6));
assign Zh3xx6 = (~(TSVALUEB[45] ^ Kkc7v6));
assign Vge8x6 = (Ni3xx6 & Ui3xx6);
assign Ui3xx6 = (~(TSVALUEB[39] ^ Gnzmz6[44]));
assign Ni3xx6 = (~(TSVALUEB[35] ^ Gnzmz6[40]));
assign Hge8x6 = (Bj3xx6 & Ij3xx6);
assign Ij3xx6 = (Pj3xx6 & Wj3xx6);
assign Wj3xx6 = (~(TSVALUEB[38] ^ Gnzmz6[43]));
assign Pj3xx6 = (~(TSVALUEB[36] ^ Gnzmz6[41]));
assign Bj3xx6 = (Dk3xx6 & Kk3xx6);
assign Kk3xx6 = (~(TSVALUEB[41] ^ Gnzmz6[46]));
assign Dk3xx6 = (~(TSVALUEB[37] ^ Gnzmz6[42]));
assign Yee8x6 = (Rk3xx6 & Yk3xx6);
assign Yk3xx6 = (~(TSVALUEB[31] ^ Gnzmz6[35]));
assign Rk3xx6 = (~(TSVALUEB[28] ^ Gnzmz6[32]));
assign Kee8x6 = (Fl3xx6 & Ml3xx6);
assign Ml3xx6 = (Tl3xx6 & Am3xx6);
assign Am3xx6 = (~(TSVALUEB[30] ^ Gnzmz6[34]));
assign Tl3xx6 = (~(TSVALUEB[29] ^ Gnzmz6[33]));
assign Fl3xx6 = (Hm3xx6 & Om3xx6);
assign Om3xx6 = (~(TSVALUEB[34] ^ Gnzmz6[38]));
assign Hm3xx6 = (~(TSVALUEB[32] ^ Gnzmz6[36]));
assign Bde8x6 = (Vm3xx6 & Cn3xx6);
assign Cn3xx6 = (~(TSVALUEB[24] ^ Gnzmz6[27]));
assign Vm3xx6 = (~(TSVALUEB[21] ^ Gnzmz6[24]));
assign Nce8x6 = (Jn3xx6 & Qn3xx6);
assign Qn3xx6 = (Xn3xx6 & Eo3xx6);
assign Eo3xx6 = (~(TSVALUEB[23] ^ Gnzmz6[26]));
assign Xn3xx6 = (~(TSVALUEB[22] ^ Gnzmz6[25]));
assign Jn3xx6 = (Lo3xx6 & So3xx6);
assign So3xx6 = (~(TSVALUEB[27] ^ Gnzmz6[30]));
assign Lo3xx6 = (~(TSVALUEB[25] ^ Gnzmz6[28]));
assign Ebe8x6 = (Zo3xx6 & Gp3xx6);
assign Gp3xx6 = (~(TSVALUEB[18] ^ Gnzmz6[20]));
assign Zo3xx6 = (~(TSVALUEB[14] ^ Gnzmz6[16]));
assign Qae8x6 = (Np3xx6 & Up3xx6);
assign Up3xx6 = (Bq3xx6 & Iq3xx6);
assign Iq3xx6 = (~(TSVALUEB[17] ^ Gnzmz6[19]));
assign Bq3xx6 = (~(TSVALUEB[15] ^ Gnzmz6[17]));
assign Np3xx6 = (Pq3xx6 & Wq3xx6);
assign Wq3xx6 = (~(TSVALUEB[20] ^ Gnzmz6[22]));
assign Pq3xx6 = (~(TSVALUEB[16] ^ Gnzmz6[18]));
assign Aqu7v6 = (Dr3xx6 ? L5zmz6[8] : P3zmz6[8]);
assign L5zmz6[8] = (Ursnv6 ? Kr3xx6 : Rjzmz6[8]);
assign Kr3xx6 = (!Kr67z6);
assign Tpu7v6 = (Dr3xx6 ? L5zmz6[9] : P3zmz6[9]);
assign L5zmz6[9] = (Ursnv6 ? Rr3xx6 : Rjzmz6[9]);
assign Rr3xx6 = (!Cr67z6);
assign Mpu7v6 = (Dr3xx6 ? L5zmz6[10] : P3zmz6[10]);
assign L5zmz6[10] = (Fs3xx6 ? Rjzmz6[10] : Yr3xx6);
assign Yr3xx6 = (!Uq67z6);
assign Fpu7v6 = (Dr3xx6 ? L5zmz6[11] : P3zmz6[11]);
assign L5zmz6[11] = (Fs3xx6 ? Rjzmz6[11] : Ms3xx6);
assign Ms3xx6 = (!Mq67z6);
assign You7v6 = (Dr3xx6 ? L5zmz6[12] : P3zmz6[12]);
assign L5zmz6[12] = (Fs3xx6 ? Rjzmz6[12] : Ts3xx6);
assign Ts3xx6 = (!Eq67z6);
assign Rou7v6 = (Dr3xx6 ? L5zmz6[13] : P3zmz6[13]);
assign L5zmz6[13] = (Ursnv6 ? At3xx6 : Rjzmz6[13]);
assign At3xx6 = (!Wp67z6);
assign Kou7v6 = (Dr3xx6 ? L5zmz6[14] : P3zmz6[14]);
assign L5zmz6[14] = (Ursnv6 ? Ht3xx6 : Rjzmz6[14]);
assign Ht3xx6 = (!Op67z6);
assign Dou7v6 = (Dr3xx6 ? L5zmz6[15] : P3zmz6[15]);
assign L5zmz6[15] = (Ursnv6 ? Ot3xx6 : Rjzmz6[15]);
assign Ot3xx6 = (!Gp67z6);
assign Wnu7v6 = (Dr3xx6 ? L5zmz6[16] : P3zmz6[16]);
assign L5zmz6[16] = (Ursnv6 ? Vt3xx6 : Rjzmz6[16]);
assign Vt3xx6 = (!Yo67z6);
assign Pnu7v6 = (Dr3xx6 ? L5zmz6[17] : P3zmz6[17]);
assign L5zmz6[17] = (Ursnv6 ? Cu3xx6 : Rjzmz6[17]);
assign Cu3xx6 = (!Qo67z6);
assign Inu7v6 = (Dr3xx6 ? L5zmz6[18] : P3zmz6[18]);
assign L5zmz6[18] = (Ursnv6 ? Ju3xx6 : Rjzmz6[18]);
assign Ju3xx6 = (!Io67z6);
assign Bnu7v6 = (Dr3xx6 ? L5zmz6[19] : P3zmz6[19]);
assign L5zmz6[19] = (Ursnv6 ? Qu3xx6 : Rjzmz6[19]);
assign Qu3xx6 = (!Ao67z6);
assign Umu7v6 = (Dr3xx6 ? Tct8v6 : P3zmz6[20]);
assign Tct8v6 = (Ursnv6 ? Slzmz6[20] : Rjzmz6[20]);
assign Nmu7v6 = (Dr3xx6 ? L5zmz6[21] : P3zmz6[21]);
assign L5zmz6[21] = (Ursnv6 ? Xu3xx6 : Rjzmz6[21]);
assign Xu3xx6 = (!Sn67z6);
assign Gmu7v6 = (Dr3xx6 ? L5zmz6[22] : P3zmz6[22]);
assign L5zmz6[22] = (Ursnv6 ? Ev3xx6 : Rjzmz6[22]);
assign Ev3xx6 = (!Kn67z6);
assign Zlu7v6 = (Dr3xx6 ? L5zmz6[23] : P3zmz6[23]);
assign L5zmz6[23] = (Ursnv6 ? Lv3xx6 : Rjzmz6[23]);
assign Lv3xx6 = (!Cn67z6);
assign Slu7v6 = (Dr3xx6 ? L5zmz6[24] : P3zmz6[24]);
assign L5zmz6[24] = (Ursnv6 ? Sv3xx6 : Rjzmz6[24]);
assign Sv3xx6 = (!Um67z6);
assign Llu7v6 = (Dr3xx6 ? L5zmz6[25] : P3zmz6[25]);
assign L5zmz6[25] = (Ursnv6 ? Zv3xx6 : Rjzmz6[25]);
assign Zv3xx6 = (!Mm67z6);
assign Elu7v6 = (Dr3xx6 ? L5zmz6[26] : P3zmz6[26]);
assign L5zmz6[26] = (Ursnv6 ? Gw3xx6 : Rjzmz6[26]);
assign Gw3xx6 = (!Em67z6);
assign Xku7v6 = (Dr3xx6 ? L5zmz6[27] : P3zmz6[27]);
assign L5zmz6[27] = (!L9vnv6);
assign L9vnv6 = (Fs3xx6 ? Nw3xx6 : Wl67z6);
assign Nw3xx6 = (!Rjzmz6[27]);
assign Qku7v6 = (Dr3xx6 ? L5zmz6[28] : P3zmz6[28]);
assign Dr3xx6 = (!Uw3xx6);
assign L5zmz6[28] = (Ursnv6 ? Bx3xx6 : Rjzmz6[28]);
assign Bx3xx6 = (!Ol67z6);
assign Jku7v6 = (Uw3xx6 ? P3zmz6[29] : L5zmz6[29]);
assign L5zmz6[29] = (Ursnv6 ? Ix3xx6 : Rjzmz6[29]);
assign Ix3xx6 = (!Gl67z6);
assign Cku7v6 = (Uw3xx6 ? P3zmz6[30] : L5zmz6[30]);
assign L5zmz6[30] = (!X8vnv6);
assign X8vnv6 = (Fs3xx6 ? Px3xx6 : Yk67z6);
assign Px3xx6 = (!Rjzmz6[30]);
assign Vju7v6 = (Uw3xx6 ? P3zmz6[31] : L5zmz6[31]);
assign L5zmz6[31] = (Ursnv6 ? Wx3xx6 : Rjzmz6[31]);
assign Wx3xx6 = (!Qk67z6);
assign Oju7v6 = (Uw3xx6 ? P3zmz6[7] : L5zmz6[7]);
assign Uw3xx6 = (~(H0vnv6 | Edo7v6));
assign H0vnv6 = (Oosnv6 | Qatnv6);
assign Qatnv6 = (Dy3xx6 & Ky3xx6);
assign Ky3xx6 = (Ry3xx6 & Yy3xx6);
assign Yy3xx6 = (~(Tkb7v6 | I9b7v6));
assign Ry3xx6 = (~(Bba7v6 | Mbc7v6));
assign Dy3xx6 = (Fz3xx6 & Mz3xx6);
assign Mz3xx6 = (Tz3xx6 & A04xx6);
assign Fz3xx6 = (~(H04xx6 | O04xx6));
assign H04xx6 = (Ro87v6 ? V04xx6 : Sqsnv6);
assign V04xx6 = (Lczmz6[1] | Gdc7v6);
assign Oosnv6 = (X4snv6 & W8zmz6[0]);
assign W8zmz6[0] = (~(C14xx6 & J14xx6));
assign J14xx6 = (~(Q14xx6 & Ymsnv6));
assign Ymsnv6 = (Wha7z6 & X14xx6);
assign Wha7z6 = (!Sqsnv6);
assign Q14xx6 = (Fnsnv6 & Kmsnv6);
assign Kmsnv6 = (E24xx6 & T8tnv6);
assign T8tnv6 = (E6rnv6 & X4snv6);
assign E6rnv6 = (!X477v6);
assign E24xx6 = (Fgzmz6[1] & L24xx6);
assign L24xx6 = (~(S24xx6 & I1c7v6));
assign S24xx6 = (X14xx6 & R0tnv6);
assign C14xx6 = (~(Z24xx6 & G34xx6));
assign G34xx6 = (Fgzmz6[0] ? U34xx6 : N34xx6);
assign U34xx6 = (B44xx6 & I44xx6);
assign I44xx6 = (~(M1tnv6 | X477v6));
assign M1tnv6 = (~(R0tnv6 | I1c7v6));
assign B44xx6 = (P7snv6 & P44xx6);
assign P44xx6 = (Sqsnv6 | Fnsnv6);
assign N34xx6 = (Fnsnv6 & Uia7v6);
assign Uia7v6 = (~(Sqsnv6 & W44xx6));
assign W44xx6 = (~(D54xx6 & Lzb7v6));
assign D54xx6 = (Xw67v6 & R0tnv6);
assign R0tnv6 = (!Z2c7v6);
assign Fnsnv6 = (K54xx6 & P7snv6);
assign P7snv6 = (Jrqnv6 & Ox67v6);
assign Ox67v6 = (~(R54xx6 & Y54xx6));
assign Y54xx6 = (~(F64xx6 & Xw67v6));
assign F64xx6 = (~(Wdtnv6 | O777v6));
assign R54xx6 = (~(Gg77v6 & M64xx6));
assign M64xx6 = (~(T64xx6 & A74xx6));
assign A74xx6 = (~(H74xx6 & O74xx6));
assign O74xx6 = (W577v6 | S677v6);
assign H74xx6 = (~(Pfo7v6 | Kwl8v6));
assign T64xx6 = (~(O777v6 | Xw67v6));
assign K54xx6 = (V74xx6 & C84xx6);
assign C84xx6 = (~(J84xx6 & Q84xx6));
assign Q84xx6 = (~(X84xx6 & Ojymz6[10]));
assign X84xx6 = (S94xx6 ? L94xx6 : E94xx6);
assign L94xx6 = (~(Z94xx6 & Ga4xx6));
assign Z94xx6 = (~(Na4xx6 & Ua4xx6));
assign Ua4xx6 = (!Ojymz6[8]);
assign E94xx6 = (Ojymz6[8] & Bb4xx6);
assign Bb4xx6 = (Ga4xx6 | Na4xx6);
assign Ga4xx6 = (!Ojymz6[9]);
assign J84xx6 = (Ojymz6[8] ? Pb4xx6 : Ib4xx6);
assign Pb4xx6 = (~(S94xx6 & Wb4xx6));
assign Wb4xx6 = (~(Na4xx6 & Dc4xx6));
assign Dc4xx6 = (Ojymz6[10] | Ojymz6[9]);
assign Ib4xx6 = (Kc4xx6 | S94xx6);
assign S94xx6 = (Rc4xx6 & Yc4xx6);
assign Yc4xx6 = (Ojymz6[0] ? Md4xx6 : Fd4xx6);
assign Md4xx6 = (~(Td4xx6 & Ae4xx6));
assign Ae4xx6 = (~(Ojymz6[1] | Ojymz6[3]));
assign Td4xx6 = (Ojymz6[2] & Oasnv6);
assign Fd4xx6 = (~(He4xx6 & Oe4xx6));
assign He4xx6 = (Ojymz6[3] ? Cf4xx6 : Ve4xx6);
assign Cf4xx6 = (Uh77v6 & Jf4xx6);
assign Ve4xx6 = (Ojymz6[2] & Ecsnv6);
assign Rc4xx6 = (Qf4xx6 & Xf4xx6);
assign Xf4xx6 = (~(Tn77v6 & Eg4xx6));
assign Qf4xx6 = (~(Ojymz6[2] & Lg4xx6));
assign Lg4xx6 = (Sg4xx6 | Eg4xx6);
assign Sg4xx6 = (~(Zg4xx6 | Oe4xx6));
assign Oe4xx6 = (!Ojymz6[1]);
assign Zg4xx6 = (Ojymz6[0] ? Iesnv6 : Gh4xx6);
assign Gh4xx6 = (Ojymz6[3] | Pesnv6);
assign Kc4xx6 = (Ojymz6[9] ? Na4xx6 : Ojymz6[10]);
assign Na4xx6 = (Nh4xx6 & Uh4xx6);
assign Uh4xx6 = (Ojymz6[4] ? Ii4xx6 : Bi4xx6);
assign Ii4xx6 = (~(Pi4xx6 & Oasnv6));
assign Oasnv6 = (!Hhsnv6);
assign Hhsnv6 = (B1rnv6 & Lgo7x6);
assign Lgo7x6 = (~(Iwymz6[1] & Zgo7x6));
assign Zgo7x6 = (Zdp7z6[1] ? Wi4xx6 : Sr67z6);
assign B1rnv6 = (!Lfp7z6[1]);
assign Bi4xx6 = (Dj4xx6 & Kj4xx6);
assign Kj4xx6 = (~(Rj4xx6 & Yj4xx6));
assign Yj4xx6 = (~(Ojymz6[5] | Ojymz6[6]));
assign Rj4xx6 = (Uh77v6 & Ojymz6[7]);
assign Dj4xx6 = (~(Pi4xx6 & Ecsnv6));
assign Ecsnv6 = (!Qisnv6);
assign Qisnv6 = (B4o7x6 & Qfo7x6);
assign Qfo7x6 = (~(Iwymz6[0] & Ego7x6));
assign Ego7x6 = (Zdp7z6[0] ? Wi4xx6 : Sr67z6);
assign B4o7x6 = (!Lfp7z6[0]);
assign Pi4xx6 = (Fk4xx6 & Ojymz6[6]);
assign Fk4xx6 = (~(Ojymz6[5] | Ojymz6[7]));
assign Nh4xx6 = (Mk4xx6 & Tk4xx6);
assign Tk4xx6 = (~(Ojymz6[6] & Al4xx6));
assign Al4xx6 = (Hl4xx6 | Ol4xx6);
assign Ol4xx6 = (Vl4xx6 & Ojymz6[5]);
assign Vl4xx6 = (Ojymz6[4] ? Uksnv6 : Cm4xx6);
assign Uksnv6 = (!Iesnv6);
assign Iesnv6 = (U0rnv6 & Bio7x6);
assign Bio7x6 = (~(Iwymz6[3] & Pio7x6));
assign Pio7x6 = (Zdp7z6[3] ? Wi4xx6 : Sr67z6);
assign U0rnv6 = (!Lfp7z6[3]);
assign Cm4xx6 = (~(Pesnv6 | Ojymz6[7]));
assign Pesnv6 = (Aeo7x6 & Gho7x6);
assign Gho7x6 = (~(Iwymz6[2] & Uho7x6));
assign Uho7x6 = (Zdp7z6[2] ? Wi4xx6 : Sr67z6);
assign Wi4xx6 = (!Q087v6);
assign Aeo7x6 = (!Lfp7z6[2]);
assign Mk4xx6 = (~(Tn77v6 & Hl4xx6));
assign V74xx6 = (~(Ok77v6 & Jm4xx6));
assign Jm4xx6 = (~(Qm4xx6 & Tn77v6));
assign Qm4xx6 = (~(Nernv6 | Gernv6));
assign Nernv6 = (~(X5rnv6 | Xu67v6));
assign X5rnv6 = (~(L877v6 & Xm4xx6));
assign X4snv6 = (!Fgzmz6[0]);
assign L5zmz6[7] = (!G3vnv6);
assign G3vnv6 = (Fs3xx6 ? En4xx6 : Ik67z6);
assign En4xx6 = (!Rjzmz6[7]);
assign Hju7v6 = (Xfd7v6 ^ Ln4xx6);
assign Ln4xx6 = (Sn4xx6 & Mz0nz6[4]);
assign Sn4xx6 = (Mz0nz6[3] & Fftnv6);
assign Aju7v6 = (Fftnv6 ? Ux0nz6[0] : E11nz6[0]);
assign Tiu7v6 = (Fftnv6 ? Ux0nz6[1] : E11nz6[1]);
assign Miu7v6 = (Fftnv6 ? Ux0nz6[2] : E11nz6[2]);
assign Fiu7v6 = (!Zn4xx6);
assign Zn4xx6 = (Vicov6 ? No4xx6 : Go4xx6);
assign Go4xx6 = (~(Mz0nz6[3] & Uo4xx6));
assign Yhu7v6 = (!Bp4xx6);
assign Bp4xx6 = (Vicov6 ? Pp4xx6 : Ip4xx6);
assign Ip4xx6 = (Uo4xx6 | Mz0nz6[3]);
assign Uo4xx6 = (!Mz0nz6[4]);
assign Rhu7v6 = (~(Wp4xx6 & Dq4xx6));
assign Dq4xx6 = (~(Uu0nz6[4] & Kq4xx6));
assign Kq4xx6 = (~(Rq4xx6 & Yq4xx6));
assign Yq4xx6 = (!Uu0nz6[3]);
assign Wp4xx6 = (~(Fr4xx6 & Mr4xx6));
assign Mr4xx6 = (~(Tr4xx6 ^ Tvrnv6));
assign Tvrnv6 = (!Zkrnv6);
assign Tr4xx6 = (~(As4xx6 & Hs4xx6));
assign Hs4xx6 = (Imrnv6 | Os4xx6);
assign As4xx6 = (Vs4xx6 | Ct4xx6);
assign Khu7v6 = (Jt4xx6 | Qt4xx6);
assign Qt4xx6 = (Xt4xx6 & Fr4xx6);
assign Xt4xx6 = (Durnv6 ^ Eu4xx6);
assign Jt4xx6 = (Uu0nz6[1] ? Su4xx6 : Lu4xx6);
assign Lu4xx6 = (Zu4xx6 & Gv4xx6);
assign Dhu7v6 = (~(Nv4xx6 & Uv4xx6));
assign Nv4xx6 = (Bw4xx6 & Iw4xx6);
assign Iw4xx6 = (~(Pw4xx6 & Fr4xx6));
assign Pw4xx6 = (Ww4xx6 ^ Dx4xx6);
assign Dx4xx6 = (Eu4xx6 & Durnv6);
assign Bw4xx6 = (~(Uu0nz6[2] & Kx4xx6));
assign Kx4xx6 = (Su4xx6 | Uu0nz6[1]);
assign Su4xx6 = (~(Rx4xx6 & Gv4xx6));
assign Gv4xx6 = (!Uu0nz6[0]);
assign Wgu7v6 = (~(Yx4xx6 & Fy4xx6));
assign Fy4xx6 = (~(My4xx6 & Fr4xx6));
assign My4xx6 = (Ct4xx6 ^ Vs4xx6);
assign Vs4xx6 = (~(Eu4xx6 & Os4xx6));
assign Eu4xx6 = (Errnv6 & A3dov6);
assign A3dov6 = (!Sr5ov6);
assign Ct4xx6 = (~(Imrnv6 ^ Os4xx6));
assign Os4xx6 = (Ww4xx6 & Durnv6);
assign Ww4xx6 = (~(Qqrnv6 ^ Durnv6));
assign Yx4xx6 = (Uu0nz6[3] ? Rq4xx6 : Uv4xx6);
assign Rq4xx6 = (Ty4xx6 & Rx4xx6);
assign Uv4xx6 = (~(Zu4xx6 & Ty4xx6));
assign Ty4xx6 = (~(Az4xx6 | Uu0nz6[0]));
assign Zu4xx6 = (!Hz4xx6);
assign Pgu7v6 = (~(Oz4xx6 & Vz4xx6));
assign Vz4xx6 = (~(C05xx6 & Fr4xx6));
assign C05xx6 = (~(Errnv6 ^ Sr5ov6));
assign Oz4xx6 = (Uu0nz6[0] ? Rx4xx6 : Hz4xx6);
assign Hz4xx6 = (~(J05xx6 & Rx4xx6));
assign Rx4xx6 = (Fr4xx6 | Sr5ov6);
assign Fr4xx6 = (Q05xx6 & X05xx6);
assign X05xx6 = (~(E15xx6 | Kkd7v6));
assign Q05xx6 = (L15xx6 & N6dov6);
assign J05xx6 = (~(L15xx6 & S15xx6));
assign Igu7v6 = (Fftnv6 ? Oha7z6 : T51nz6[0]);
assign Bgu7v6 = (Fftnv6 ? Gha7z6 : T51nz6[1]);
assign Ufu7v6 = (~(Z15xx6 & G25xx6));
assign G25xx6 = (~(T51nz6[2] & Vicov6));
assign Vicov6 = (!Fftnv6);
assign Nfu7v6 = (~(N25xx6 & U25xx6));
assign U25xx6 = (~(B41nz6[1] & B35xx6));
assign Gfu7v6 = (~(I35xx6 & P35xx6));
assign P35xx6 = (~(B41nz6[0] & B35xx6));
assign Zeu7v6 = (D45xx6 ? W35xx6 : Bq0nz6[0]);
assign Seu7v6 = (K45xx6 ? W35xx6 : Lo0nz6[0]);
assign Leu7v6 = (R45xx6 ? W35xx6 : Vm0nz6[0]);
assign W35xx6 = (R21nz6[2] ? F55xx6 : Y45xx6);
assign Eeu7v6 = (D45xx6 ? M55xx6 : Bq0nz6[1]);
assign Xdu7v6 = (K45xx6 ? M55xx6 : Lo0nz6[1]);
assign Qdu7v6 = (R45xx6 ? M55xx6 : Vm0nz6[1]);
assign M55xx6 = (R21nz6[2] ? A65xx6 : T55xx6);
assign Jdu7v6 = (D45xx6 ? H65xx6 : Bq0nz6[2]);
assign Cdu7v6 = (K45xx6 ? H65xx6 : Lo0nz6[2]);
assign Vcu7v6 = (R45xx6 ? H65xx6 : Vm0nz6[2]);
assign H65xx6 = (R21nz6[2] ? V65xx6 : O65xx6);
assign Ocu7v6 = (D45xx6 ? C75xx6 : Bq0nz6[3]);
assign Hcu7v6 = (K45xx6 ? C75xx6 : Lo0nz6[3]);
assign Acu7v6 = (R45xx6 ? C75xx6 : Vm0nz6[3]);
assign C75xx6 = (R21nz6[2] ? Q75xx6 : J75xx6);
assign Tbu7v6 = (D45xx6 ? X75xx6 : Bq0nz6[4]);
assign Mbu7v6 = (K45xx6 ? X75xx6 : Lo0nz6[4]);
assign Fbu7v6 = (R45xx6 ? X75xx6 : Vm0nz6[4]);
assign X75xx6 = (R21nz6[2] ? L85xx6 : E85xx6);
assign Yau7v6 = (D45xx6 ? S85xx6 : Bq0nz6[5]);
assign Rau7v6 = (K45xx6 ? S85xx6 : Lo0nz6[5]);
assign Kau7v6 = (R45xx6 ? S85xx6 : Vm0nz6[5]);
assign S85xx6 = (R21nz6[2] ? G95xx6 : Z85xx6);
assign Dau7v6 = (D45xx6 ? N95xx6 : Bq0nz6[6]);
assign W9u7v6 = (K45xx6 ? N95xx6 : Lo0nz6[6]);
assign P9u7v6 = (R45xx6 ? N95xx6 : Vm0nz6[6]);
assign N95xx6 = (R21nz6[2] ? Ba5xx6 : U95xx6);
assign I9u7v6 = (D45xx6 ? Ia5xx6 : Bq0nz6[7]);
assign D45xx6 = (~(Pa5xx6 | Wa5xx6));
assign Pa5xx6 = (Db5xx6 | Kb5xx6);
assign B9u7v6 = (K45xx6 ? Ia5xx6 : Lo0nz6[7]);
assign K45xx6 = (Rb5xx6 & Wa5xx6);
assign Rb5xx6 = (~(Db5xx6 | Kb5xx6));
assign U8u7v6 = (R45xx6 ? Ia5xx6 : Vm0nz6[7]);
assign R45xx6 = (Yb5xx6 & Db5xx6);
assign Db5xx6 = (Mc5xx6 ? B41nz6[1] : Fc5xx6);
assign Yb5xx6 = (~(Wa5xx6 | Kb5xx6));
assign Kb5xx6 = (Tc5xx6 & Ad5xx6);
assign Ad5xx6 = (~(Mc5xx6 & Hd5xx6));
assign Hd5xx6 = (~(Od5xx6 & Vd5xx6));
assign Vd5xx6 = (~(Oha7z6 & Fftnv6));
assign Tc5xx6 = (~(Ce5xx6 & Je5xx6));
assign Je5xx6 = (~(Qe5xx6 & Xe5xx6));
assign Wa5xx6 = (Mc5xx6 ? B41nz6[0] : Ef5xx6);
assign Mc5xx6 = (~(Lf5xx6 | T51nz6[0]));
assign Ia5xx6 = (R21nz6[2] ? Zf5xx6 : Sf5xx6);
assign N8u7v6 = (Ng5xx6 ? Gg5xx6 : Fl0nz6[0]);
assign G8u7v6 = (Ug5xx6 ? Gg5xx6 : Pj0nz6[0]);
assign Z7u7v6 = (Bh5xx6 ? Gg5xx6 : Zh0nz6[0]);
assign Gg5xx6 = (R21nz6[2] ? Ph5xx6 : Ih5xx6);
assign S7u7v6 = (Ng5xx6 ? Wh5xx6 : Fl0nz6[1]);
assign L7u7v6 = (Ug5xx6 ? Wh5xx6 : Pj0nz6[1]);
assign E7u7v6 = (Bh5xx6 ? Wh5xx6 : Zh0nz6[1]);
assign Wh5xx6 = (R21nz6[2] ? Ki5xx6 : Di5xx6);
assign X6u7v6 = (Ng5xx6 ? Ri5xx6 : Fl0nz6[2]);
assign Q6u7v6 = (Ug5xx6 ? Ri5xx6 : Pj0nz6[2]);
assign J6u7v6 = (Bh5xx6 ? Ri5xx6 : Zh0nz6[2]);
assign Ri5xx6 = (R21nz6[2] ? Fj5xx6 : Yi5xx6);
assign C6u7v6 = (Ng5xx6 ? Mj5xx6 : Fl0nz6[3]);
assign V5u7v6 = (Ug5xx6 ? Mj5xx6 : Pj0nz6[3]);
assign O5u7v6 = (Bh5xx6 ? Mj5xx6 : Zh0nz6[3]);
assign Mj5xx6 = (R21nz6[2] ? Ak5xx6 : Tj5xx6);
assign H5u7v6 = (Ng5xx6 ? Hk5xx6 : Fl0nz6[4]);
assign A5u7v6 = (Ug5xx6 ? Hk5xx6 : Pj0nz6[4]);
assign T4u7v6 = (Bh5xx6 ? Hk5xx6 : Zh0nz6[4]);
assign Hk5xx6 = (R21nz6[2] ? Vk5xx6 : Ok5xx6);
assign M4u7v6 = (Ng5xx6 ? Cl5xx6 : Fl0nz6[5]);
assign F4u7v6 = (Ug5xx6 ? Cl5xx6 : Pj0nz6[5]);
assign Y3u7v6 = (Bh5xx6 ? Cl5xx6 : Zh0nz6[5]);
assign Cl5xx6 = (R21nz6[2] ? Ql5xx6 : Jl5xx6);
assign R3u7v6 = (Ng5xx6 ? Xl5xx6 : Fl0nz6[6]);
assign K3u7v6 = (Ug5xx6 ? Xl5xx6 : Pj0nz6[6]);
assign D3u7v6 = (Bh5xx6 ? Xl5xx6 : Zh0nz6[6]);
assign Xl5xx6 = (R21nz6[2] ? Lm5xx6 : Em5xx6);
assign W2u7v6 = (Ng5xx6 ? Sm5xx6 : Fl0nz6[7]);
assign Ng5xx6 = (Zm5xx6 & Gn5xx6);
assign P2u7v6 = (Ug5xx6 ? Sm5xx6 : Pj0nz6[7]);
assign Ug5xx6 = (Zm5xx6 & Nn5xx6);
assign Zm5xx6 = (Un5xx6 & Bo5xx6);
assign Un5xx6 = (!Io5xx6);
assign I2u7v6 = (Bh5xx6 ? Sm5xx6 : Zh0nz6[7]);
assign Bh5xx6 = (Po5xx6 & Io5xx6);
assign Io5xx6 = (Wo5xx6 ? B41nz6[1] : Fc5xx6);
assign Po5xx6 = (Gn5xx6 & Bo5xx6);
assign Bo5xx6 = (~(Dp5xx6 & Kp5xx6));
assign Kp5xx6 = (B35xx6 | Qe5xx6);
assign Qe5xx6 = (Rp5xx6 & Yp5xx6);
assign Dp5xx6 = (Lf5xx6 | Od5xx6);
assign Od5xx6 = (Fq5xx6 & Mq5xx6);
assign Mq5xx6 = (~(Gha7z6 & Fftnv6));
assign Gn5xx6 = (!Nn5xx6);
assign Nn5xx6 = (Wo5xx6 ? B41nz6[0] : Ef5xx6);
assign Sm5xx6 = (R21nz6[2] ? Ar5xx6 : Tq5xx6);
assign B2u7v6 = (Or5xx6 ? Hr5xx6 : Jg0nz6[0]);
assign U1u7v6 = (Vr5xx6 ? Hr5xx6 : Te0nz6[0]);
assign N1u7v6 = (Cs5xx6 ? Hr5xx6 : Dd0nz6[0]);
assign Hr5xx6 = (R21nz6[2] ? Qs5xx6 : Js5xx6);
assign G1u7v6 = (Or5xx6 ? Xs5xx6 : Jg0nz6[1]);
assign Z0u7v6 = (Vr5xx6 ? Xs5xx6 : Te0nz6[1]);
assign S0u7v6 = (Cs5xx6 ? Xs5xx6 : Dd0nz6[1]);
assign Xs5xx6 = (R21nz6[2] ? Lt5xx6 : Et5xx6);
assign L0u7v6 = (Or5xx6 ? St5xx6 : Jg0nz6[2]);
assign E0u7v6 = (Vr5xx6 ? St5xx6 : Te0nz6[2]);
assign Xzt7v6 = (Cs5xx6 ? St5xx6 : Dd0nz6[2]);
assign St5xx6 = (R21nz6[2] ? Gu5xx6 : Zt5xx6);
assign Qzt7v6 = (Or5xx6 ? Nu5xx6 : Jg0nz6[3]);
assign Jzt7v6 = (Vr5xx6 ? Nu5xx6 : Te0nz6[3]);
assign Czt7v6 = (Cs5xx6 ? Nu5xx6 : Dd0nz6[3]);
assign Nu5xx6 = (R21nz6[2] ? Bv5xx6 : Uu5xx6);
assign Vyt7v6 = (Or5xx6 ? Iv5xx6 : Jg0nz6[4]);
assign Oyt7v6 = (Vr5xx6 ? Iv5xx6 : Te0nz6[4]);
assign Hyt7v6 = (Cs5xx6 ? Iv5xx6 : Dd0nz6[4]);
assign Iv5xx6 = (R21nz6[2] ? Wv5xx6 : Pv5xx6);
assign Ayt7v6 = (Or5xx6 ? Dw5xx6 : Jg0nz6[5]);
assign Txt7v6 = (Vr5xx6 ? Dw5xx6 : Te0nz6[5]);
assign Mxt7v6 = (Cs5xx6 ? Dw5xx6 : Dd0nz6[5]);
assign Dw5xx6 = (R21nz6[2] ? Rw5xx6 : Kw5xx6);
assign Fxt7v6 = (Or5xx6 ? Yw5xx6 : Jg0nz6[6]);
assign Ywt7v6 = (Vr5xx6 ? Yw5xx6 : Te0nz6[6]);
assign Rwt7v6 = (Cs5xx6 ? Yw5xx6 : Dd0nz6[6]);
assign Yw5xx6 = (R21nz6[2] ? Mx5xx6 : Fx5xx6);
assign Kwt7v6 = (Or5xx6 ? Tx5xx6 : Jg0nz6[7]);
assign Or5xx6 = (Ay5xx6 & Hy5xx6);
assign Dwt7v6 = (Vr5xx6 ? Tx5xx6 : Te0nz6[7]);
assign Vr5xx6 = (Ay5xx6 & Oy5xx6);
assign Ay5xx6 = (Vy5xx6 & Cz5xx6);
assign Vy5xx6 = (!Jz5xx6);
assign Wvt7v6 = (Cs5xx6 ? Tx5xx6 : Dd0nz6[7]);
assign Cs5xx6 = (Qz5xx6 & Jz5xx6);
assign Jz5xx6 = (Xz5xx6 ? Fc5xx6 : B41nz6[1]);
assign Qz5xx6 = (Hy5xx6 & Cz5xx6);
assign Cz5xx6 = (~(E06xx6 & L06xx6));
assign E06xx6 = (S06xx6 & Z06xx6);
assign Z06xx6 = (~(G16xx6 & Gha7z6));
assign G16xx6 = (Oha7z6 & N16xx6);
assign N16xx6 = (~(B35xx6 & U16xx6));
assign U16xx6 = (~(Fftnv6 & B26xx6));
assign S06xx6 = (Xz5xx6 | Fq5xx6);
assign Hy5xx6 = (!Oy5xx6);
assign Oy5xx6 = (Xz5xx6 ? Ef5xx6 : B41nz6[0]);
assign Xz5xx6 = (!B26xx6);
assign B26xx6 = (~(I26xx6 & Lf5xx6));
assign Lf5xx6 = (!Wo5xx6);
assign Wo5xx6 = (P26xx6 & W26xx6);
assign I26xx6 = (~(W26xx6 & D36xx6));
assign D36xx6 = (!T51nz6[0]);
assign Tx5xx6 = (R21nz6[2] ? R36xx6 : K36xx6);
assign Pvt7v6 = (F46xx6 ? Y36xx6 : Nb0nz6[0]);
assign Ivt7v6 = (M46xx6 ? Y36xx6 : X90nz6[0]);
assign Bvt7v6 = (T46xx6 ? Y36xx6 : H80nz6[0]);
assign Y36xx6 = (R21nz6[2] ? H56xx6 : A56xx6);
assign Uut7v6 = (F46xx6 ? O56xx6 : Nb0nz6[1]);
assign Nut7v6 = (M46xx6 ? O56xx6 : X90nz6[1]);
assign Gut7v6 = (T46xx6 ? O56xx6 : H80nz6[1]);
assign O56xx6 = (R21nz6[2] ? C66xx6 : V56xx6);
assign Ztt7v6 = (F46xx6 ? J66xx6 : Nb0nz6[2]);
assign Stt7v6 = (M46xx6 ? J66xx6 : X90nz6[2]);
assign Ltt7v6 = (T46xx6 ? J66xx6 : H80nz6[2]);
assign J66xx6 = (R21nz6[2] ? X66xx6 : Q66xx6);
assign Ett7v6 = (F46xx6 ? E76xx6 : Nb0nz6[3]);
assign Xst7v6 = (M46xx6 ? E76xx6 : X90nz6[3]);
assign Qst7v6 = (T46xx6 ? E76xx6 : H80nz6[3]);
assign E76xx6 = (R21nz6[2] ? S76xx6 : L76xx6);
assign Jst7v6 = (F46xx6 ? Z76xx6 : Nb0nz6[4]);
assign Cst7v6 = (M46xx6 ? Z76xx6 : X90nz6[4]);
assign Vrt7v6 = (T46xx6 ? Z76xx6 : H80nz6[4]);
assign Z76xx6 = (R21nz6[2] ? N86xx6 : G86xx6);
assign Ort7v6 = (F46xx6 ? U86xx6 : Nb0nz6[5]);
assign Hrt7v6 = (M46xx6 ? U86xx6 : X90nz6[5]);
assign Art7v6 = (T46xx6 ? U86xx6 : H80nz6[5]);
assign U86xx6 = (R21nz6[2] ? I96xx6 : B96xx6);
assign Tqt7v6 = (F46xx6 ? P96xx6 : Nb0nz6[6]);
assign Mqt7v6 = (M46xx6 ? P96xx6 : X90nz6[6]);
assign Fqt7v6 = (T46xx6 ? P96xx6 : H80nz6[6]);
assign P96xx6 = (R21nz6[2] ? Da6xx6 : W96xx6);
assign Ypt7v6 = (F46xx6 ? Ka6xx6 : Nb0nz6[7]);
assign F46xx6 = (Ra6xx6 & Ya6xx6);
assign Rpt7v6 = (M46xx6 ? Ka6xx6 : X90nz6[7]);
assign M46xx6 = (Ra6xx6 & Fb6xx6);
assign Ra6xx6 = (Mb6xx6 & Tb6xx6);
assign Mb6xx6 = (!Ac6xx6);
assign Kpt7v6 = (T46xx6 ? Ka6xx6 : H80nz6[7]);
assign T46xx6 = (Hc6xx6 & Ac6xx6);
assign Ac6xx6 = (T51nz6[2] ? Fc5xx6 : B41nz6[1]);
assign Hc6xx6 = (Ya6xx6 & Tb6xx6);
assign Tb6xx6 = (~(L06xx6 & Oc6xx6));
assign Oc6xx6 = (Fq5xx6 | T51nz6[2]);
assign Fq5xx6 = (Z15xx6 & B35xx6);
assign Z15xx6 = (!Vc6xx6);
assign L06xx6 = (~(Ce5xx6 & Mho7v6));
assign Ya6xx6 = (!Fb6xx6);
assign Fb6xx6 = (T51nz6[2] ? Ef5xx6 : B41nz6[0]);
assign Ka6xx6 = (R21nz6[2] ? Jd6xx6 : Cd6xx6);
assign Dpt7v6 = (Xd6xx6 ? Qd6xx6 : R60nz6[0]);
assign Wot7v6 = (Ee6xx6 ? Qd6xx6 : B50nz6[0]);
assign Pot7v6 = (Le6xx6 ? Qd6xx6 : L30nz6[0]);
assign Qd6xx6 = (R21nz6[2] ? Y45xx6 : F55xx6);
assign Y45xx6 = (~(Se6xx6 & Ze6xx6));
assign Ze6xx6 = (Gf6xx6 | Nf6xx6);
assign Se6xx6 = (Uf6xx6 & Bg6xx6);
assign Bg6xx6 = (Ig6xx6 | R21nz6[1]);
assign Uf6xx6 = (Pg6xx6 | Wg6xx6);
assign F55xx6 = (~(Dh6xx6 & Kh6xx6));
assign Kh6xx6 = (Rh6xx6 & Yh6xx6);
assign Yh6xx6 = (Pg6xx6 | Fi6xx6);
assign Rh6xx6 = (Gf6xx6 | Mi6xx6);
assign Dh6xx6 = (Ti6xx6 & Aj6xx6);
assign Aj6xx6 = (Hj6xx6 | Oj6xx6);
assign Ti6xx6 = (Vj6xx6 | Ck6xx6);
assign Iot7v6 = (Xd6xx6 ? Jk6xx6 : R60nz6[1]);
assign Bot7v6 = (Ee6xx6 ? Jk6xx6 : B50nz6[1]);
assign Unt7v6 = (Le6xx6 ? Jk6xx6 : L30nz6[1]);
assign Jk6xx6 = (R21nz6[2] ? T55xx6 : A65xx6);
assign T55xx6 = (~(Qk6xx6 & Xk6xx6));
assign Xk6xx6 = (El6xx6 & Ll6xx6);
assign Ll6xx6 = (Sl6xx6 | Vj6xx6);
assign El6xx6 = (Gf6xx6 | Zl6xx6);
assign Qk6xx6 = (Gm6xx6 & Nm6xx6);
assign Nm6xx6 = (Pg6xx6 | Um6xx6);
assign Gm6xx6 = (Hj6xx6 | Bn6xx6);
assign A65xx6 = (~(In6xx6 & Pn6xx6));
assign Pn6xx6 = (Wn6xx6 & Do6xx6);
assign Do6xx6 = (Gf6xx6 | Ko6xx6);
assign Wn6xx6 = (Pg6xx6 | Ro6xx6);
assign In6xx6 = (Yo6xx6 & Fp6xx6);
assign Fp6xx6 = (Hj6xx6 | Mp6xx6);
assign Yo6xx6 = (Vj6xx6 | Tp6xx6);
assign Nnt7v6 = (Xd6xx6 ? Aq6xx6 : R60nz6[2]);
assign Gnt7v6 = (Ee6xx6 ? Aq6xx6 : B50nz6[2]);
assign Zmt7v6 = (Le6xx6 ? Aq6xx6 : L30nz6[2]);
assign Aq6xx6 = (R21nz6[2] ? O65xx6 : V65xx6);
assign O65xx6 = (~(Hq6xx6 & Oq6xx6));
assign Oq6xx6 = (Vq6xx6 & Cr6xx6);
assign Cr6xx6 = (Vj6xx6 | Jr6xx6);
assign Vq6xx6 = (Gf6xx6 | Qr6xx6);
assign Hq6xx6 = (Xr6xx6 & Es6xx6);
assign Es6xx6 = (Pg6xx6 | Ls6xx6);
assign Xr6xx6 = (Hj6xx6 | Ss6xx6);
assign V65xx6 = (~(Zs6xx6 & Gt6xx6));
assign Gt6xx6 = (Nt6xx6 & Ut6xx6);
assign Ut6xx6 = (Gf6xx6 | Bu6xx6);
assign Nt6xx6 = (Pg6xx6 | Iu6xx6);
assign Zs6xx6 = (Pu6xx6 & Wu6xx6);
assign Wu6xx6 = (Hj6xx6 | Dv6xx6);
assign Pu6xx6 = (Vj6xx6 | Kv6xx6);
assign Smt7v6 = (Xd6xx6 ? Rv6xx6 : R60nz6[3]);
assign Lmt7v6 = (Ee6xx6 ? Rv6xx6 : B50nz6[3]);
assign Emt7v6 = (Le6xx6 ? Rv6xx6 : L30nz6[3]);
assign Rv6xx6 = (R21nz6[2] ? J75xx6 : Q75xx6);
assign J75xx6 = (~(Yv6xx6 & Fw6xx6));
assign Fw6xx6 = (Mw6xx6 & Tw6xx6);
assign Tw6xx6 = (Vj6xx6 | Ax6xx6);
assign Mw6xx6 = (Hj6xx6 | Hx6xx6);
assign Yv6xx6 = (Ox6xx6 & Vx6xx6);
assign Vx6xx6 = (Gf6xx6 | Cy6xx6);
assign Ox6xx6 = (Pg6xx6 | Jy6xx6);
assign Q75xx6 = (~(Qy6xx6 & Xy6xx6));
assign Xy6xx6 = (Ez6xx6 & Lz6xx6);
assign Lz6xx6 = (Gf6xx6 | Sz6xx6);
assign Ez6xx6 = (Pg6xx6 | Zz6xx6);
assign Qy6xx6 = (G07xx6 & N07xx6);
assign N07xx6 = (Hj6xx6 | U07xx6);
assign G07xx6 = (Vj6xx6 | B17xx6);
assign Xlt7v6 = (Xd6xx6 ? I17xx6 : R60nz6[4]);
assign Qlt7v6 = (Ee6xx6 ? I17xx6 : B50nz6[4]);
assign Jlt7v6 = (Le6xx6 ? I17xx6 : L30nz6[4]);
assign I17xx6 = (R21nz6[2] ? E85xx6 : L85xx6);
assign E85xx6 = (~(P17xx6 & W17xx6));
assign W17xx6 = (D27xx6 & K27xx6);
assign K27xx6 = (Vj6xx6 | R27xx6);
assign D27xx6 = (Hj6xx6 | Y27xx6);
assign P17xx6 = (F37xx6 & M37xx6);
assign M37xx6 = (Gf6xx6 | T37xx6);
assign F37xx6 = (Pg6xx6 | A47xx6);
assign L85xx6 = (~(H47xx6 & O47xx6));
assign O47xx6 = (V47xx6 & C57xx6);
assign C57xx6 = (Gf6xx6 | J57xx6);
assign V47xx6 = (Pg6xx6 | Q57xx6);
assign H47xx6 = (X57xx6 & E67xx6);
assign E67xx6 = (Hj6xx6 | L67xx6);
assign X57xx6 = (Vj6xx6 | S67xx6);
assign Clt7v6 = (Xd6xx6 ? Z67xx6 : R60nz6[5]);
assign Vkt7v6 = (Ee6xx6 ? Z67xx6 : B50nz6[5]);
assign Okt7v6 = (Le6xx6 ? Z67xx6 : L30nz6[5]);
assign Z67xx6 = (R21nz6[2] ? Z85xx6 : G95xx6);
assign Z85xx6 = (~(G77xx6 & N77xx6));
assign N77xx6 = (U77xx6 & B87xx6);
assign B87xx6 = (Vj6xx6 | I87xx6);
assign U77xx6 = (Hj6xx6 | P87xx6);
assign G77xx6 = (W87xx6 & D97xx6);
assign D97xx6 = (Gf6xx6 | K97xx6);
assign W87xx6 = (Pg6xx6 | R97xx6);
assign G95xx6 = (~(Y97xx6 & Fa7xx6));
assign Fa7xx6 = (Ma7xx6 & Ta7xx6);
assign Ta7xx6 = (Gf6xx6 | Ab7xx6);
assign Ma7xx6 = (Pg6xx6 | Hb7xx6);
assign Y97xx6 = (Ob7xx6 & Vb7xx6);
assign Vb7xx6 = (Hj6xx6 | Cc7xx6);
assign Ob7xx6 = (Vj6xx6 | Jc7xx6);
assign Hkt7v6 = (Xd6xx6 ? Qc7xx6 : R60nz6[6]);
assign Akt7v6 = (Ee6xx6 ? Qc7xx6 : B50nz6[6]);
assign Tjt7v6 = (Le6xx6 ? Qc7xx6 : L30nz6[6]);
assign Qc7xx6 = (R21nz6[2] ? U95xx6 : Ba5xx6);
assign U95xx6 = (~(Xc7xx6 & Ed7xx6));
assign Ed7xx6 = (Ld7xx6 & Sd7xx6);
assign Sd7xx6 = (~(Zd7xx6 & Ge7xx6));
assign Ld7xx6 = (Ne7xx6 | Vj6xx6);
assign Xc7xx6 = (Ue7xx6 & Bf7xx6);
assign Bf7xx6 = (Gf6xx6 | If7xx6);
assign Ue7xx6 = (Pg6xx6 | Pf7xx6);
assign Ba5xx6 = (~(Wf7xx6 & Dg7xx6));
assign Dg7xx6 = (Kg7xx6 & Rg7xx6);
assign Rg7xx6 = (Gf6xx6 | Yg7xx6);
assign Kg7xx6 = (Pg6xx6 | Fh7xx6);
assign Wf7xx6 = (Mh7xx6 & Th7xx6);
assign Th7xx6 = (Hj6xx6 | Ai7xx6);
assign Mh7xx6 = (Vj6xx6 | Hi7xx6);
assign Mjt7v6 = (Xd6xx6 ? Oi7xx6 : R60nz6[7]);
assign Xd6xx6 = (Vi7xx6 & Cj7xx6);
assign Fjt7v6 = (Ee6xx6 ? Oi7xx6 : B50nz6[7]);
assign Ee6xx6 = (Vi7xx6 & Jj7xx6);
assign Vi7xx6 = (Qj7xx6 & Xj7xx6);
assign Qj7xx6 = (!Ek7xx6);
assign Yit7v6 = (Le6xx6 ? Oi7xx6 : L30nz6[7]);
assign Le6xx6 = (Lk7xx6 & Ek7xx6);
assign Ek7xx6 = (Sk7xx6 ? B41nz6[1] : Fc5xx6);
assign Lk7xx6 = (Cj7xx6 & Xj7xx6);
assign Xj7xx6 = (~(Zk7xx6 & Gl7xx6));
assign Gl7xx6 = (~(Sk7xx6 & Ce5xx6));
assign Zk7xx6 = (~(Nl7xx6 & Vc6xx6));
assign Nl7xx6 = (Ul7xx6 & Bm7xx6);
assign Bm7xx6 = (~(Im7xx6 & B35xx6));
assign Ul7xx6 = (~(Rp5xx6 & Xe5xx6));
assign Xe5xx6 = (!Oha7z6);
assign Rp5xx6 = (!Gha7z6);
assign Cj7xx6 = (!Jj7xx6);
assign Jj7xx6 = (Sk7xx6 ? B41nz6[0] : Ef5xx6);
assign Sk7xx6 = (!Im7xx6);
assign Im7xx6 = (~(Pm7xx6 & Wm7xx6));
assign Wm7xx6 = (~(T51nz6[2] & T51nz6[0]));
assign Oi7xx6 = (R21nz6[2] ? Sf5xx6 : Zf5xx6);
assign Sf5xx6 = (~(Dn7xx6 & Kn7xx6));
assign Kn7xx6 = (Pg6xx6 | Rn7xx6);
assign Dn7xx6 = (Yn7xx6 & Fo7xx6);
assign Fo7xx6 = (Mo7xx6 | R21nz6[1]);
assign Yn7xx6 = (Gf6xx6 | To7xx6);
assign Zf5xx6 = (~(Ap7xx6 & Hp7xx6));
assign Hp7xx6 = (Op7xx6 & Vp7xx6);
assign Vp7xx6 = (Gf6xx6 | Cq7xx6);
assign Op7xx6 = (Pg6xx6 | Jq7xx6);
assign Ap7xx6 = (Qq7xx6 & Xq7xx6);
assign Xq7xx6 = (Hj6xx6 | Er7xx6);
assign Qq7xx6 = (Vj6xx6 | Lr7xx6);
assign Rit7v6 = (Zr7xx6 ? Sr7xx6 : V10nz6[0]);
assign Kit7v6 = (Gs7xx6 ? Sr7xx6 : F00nz6[0]);
assign Dit7v6 = (Ns7xx6 ? Sr7xx6 : Pyzmz6[0]);
assign Sr7xx6 = (R21nz6[2] ? Ih5xx6 : Ph5xx6);
assign Ih5xx6 = (~(Us7xx6 & Bt7xx6));
assign Bt7xx6 = (~(Ge7xx6 & It7xx6));
assign Us7xx6 = (Pt7xx6 & Wt7xx6);
assign Wt7xx6 = (Vj6xx6 | Mi6xx6);
assign Pt7xx6 = (Du7xx6 | Ku7xx6);
assign Ph5xx6 = (~(Ru7xx6 & Yu7xx6));
assign Yu7xx6 = (Fv7xx6 & Mv7xx6);
assign Mv7xx6 = (Gf6xx6 | Fi6xx6);
assign Fv7xx6 = (Pg6xx6 | Oj6xx6);
assign Ru7xx6 = (Tv7xx6 & Aw7xx6);
assign Aw7xx6 = (Hj6xx6 | Ck6xx6);
assign Tv7xx6 = (Vj6xx6 | Nf6xx6);
assign Wht7v6 = (Zr7xx6 ? Hw7xx6 : V10nz6[1]);
assign Pht7v6 = (Gs7xx6 ? Hw7xx6 : F00nz6[1]);
assign Iht7v6 = (Ns7xx6 ? Hw7xx6 : Pyzmz6[1]);
assign Hw7xx6 = (R21nz6[2] ? Di5xx6 : Ki5xx6);
assign Di5xx6 = (~(Ow7xx6 & Vw7xx6));
assign Vw7xx6 = (Cx7xx6 & Jx7xx6);
assign Jx7xx6 = (Sl6xx6 | Hj6xx6);
assign Cx7xx6 = (Vj6xx6 | Ko6xx6);
assign Ow7xx6 = (Qx7xx6 & Xx7xx6);
assign Xx7xx6 = (Gf6xx6 | Um6xx6);
assign Qx7xx6 = (Pg6xx6 | Bn6xx6);
assign Ki5xx6 = (~(Ey7xx6 & Ly7xx6));
assign Ly7xx6 = (Sy7xx6 & Zy7xx6);
assign Zy7xx6 = (Gf6xx6 | Ro6xx6);
assign Sy7xx6 = (Pg6xx6 | Mp6xx6);
assign Ey7xx6 = (Gz7xx6 & Nz7xx6);
assign Nz7xx6 = (Vj6xx6 | Zl6xx6);
assign Gz7xx6 = (Hj6xx6 | Tp6xx6);
assign Bht7v6 = (Zr7xx6 ? Uz7xx6 : V10nz6[2]);
assign Ugt7v6 = (Gs7xx6 ? Uz7xx6 : F00nz6[2]);
assign Ngt7v6 = (Ns7xx6 ? Uz7xx6 : Pyzmz6[2]);
assign Uz7xx6 = (R21nz6[2] ? Yi5xx6 : Fj5xx6);
assign Yi5xx6 = (~(B08xx6 & I08xx6));
assign I08xx6 = (P08xx6 & W08xx6);
assign W08xx6 = (Hj6xx6 | Jr6xx6);
assign P08xx6 = (Vj6xx6 | Bu6xx6);
assign B08xx6 = (D18xx6 & K18xx6);
assign K18xx6 = (Gf6xx6 | Ls6xx6);
assign D18xx6 = (Pg6xx6 | Ss6xx6);
assign Fj5xx6 = (~(R18xx6 & Y18xx6));
assign Y18xx6 = (F28xx6 & M28xx6);
assign M28xx6 = (Gf6xx6 | Iu6xx6);
assign F28xx6 = (Pg6xx6 | Dv6xx6);
assign R18xx6 = (T28xx6 & A38xx6);
assign A38xx6 = (Vj6xx6 | Qr6xx6);
assign T28xx6 = (Hj6xx6 | Kv6xx6);
assign Ggt7v6 = (Zr7xx6 ? H38xx6 : V10nz6[3]);
assign Zft7v6 = (Gs7xx6 ? H38xx6 : F00nz6[3]);
assign Sft7v6 = (Ns7xx6 ? H38xx6 : Pyzmz6[3]);
assign H38xx6 = (R21nz6[2] ? Tj5xx6 : Ak5xx6);
assign Tj5xx6 = (~(O38xx6 & V38xx6));
assign V38xx6 = (C48xx6 & J48xx6);
assign J48xx6 = (Hj6xx6 | Ax6xx6);
assign C48xx6 = (Vj6xx6 | Sz6xx6);
assign O38xx6 = (Q48xx6 & X48xx6);
assign X48xx6 = (Pg6xx6 | Hx6xx6);
assign Q48xx6 = (Gf6xx6 | Jy6xx6);
assign Ak5xx6 = (~(E58xx6 & L58xx6));
assign L58xx6 = (S58xx6 & Z58xx6);
assign Z58xx6 = (Gf6xx6 | Zz6xx6);
assign S58xx6 = (Pg6xx6 | U07xx6);
assign E58xx6 = (G68xx6 & N68xx6);
assign N68xx6 = (Vj6xx6 | Cy6xx6);
assign G68xx6 = (Hj6xx6 | B17xx6);
assign Lft7v6 = (Zr7xx6 ? U68xx6 : V10nz6[4]);
assign Eft7v6 = (Gs7xx6 ? U68xx6 : F00nz6[4]);
assign Xet7v6 = (Ns7xx6 ? U68xx6 : Pyzmz6[4]);
assign U68xx6 = (R21nz6[2] ? Ok5xx6 : Vk5xx6);
assign Ok5xx6 = (~(B78xx6 & I78xx6));
assign I78xx6 = (P78xx6 & W78xx6);
assign W78xx6 = (Hj6xx6 | R27xx6);
assign P78xx6 = (Vj6xx6 | J57xx6);
assign B78xx6 = (D88xx6 & K88xx6);
assign K88xx6 = (Pg6xx6 | Y27xx6);
assign D88xx6 = (Gf6xx6 | A47xx6);
assign Vk5xx6 = (~(R88xx6 & Y88xx6));
assign Y88xx6 = (F98xx6 & M98xx6);
assign M98xx6 = (Gf6xx6 | Q57xx6);
assign F98xx6 = (Pg6xx6 | L67xx6);
assign R88xx6 = (T98xx6 & Aa8xx6);
assign Aa8xx6 = (Vj6xx6 | T37xx6);
assign T98xx6 = (Hj6xx6 | S67xx6);
assign Qet7v6 = (Zr7xx6 ? Ha8xx6 : V10nz6[5]);
assign Jet7v6 = (Gs7xx6 ? Ha8xx6 : F00nz6[5]);
assign Cet7v6 = (Ns7xx6 ? Ha8xx6 : Pyzmz6[5]);
assign Ha8xx6 = (R21nz6[2] ? Jl5xx6 : Ql5xx6);
assign Jl5xx6 = (~(Oa8xx6 & Va8xx6));
assign Va8xx6 = (Cb8xx6 & Jb8xx6);
assign Jb8xx6 = (Hj6xx6 | I87xx6);
assign Cb8xx6 = (Vj6xx6 | Ab7xx6);
assign Oa8xx6 = (Qb8xx6 & Xb8xx6);
assign Xb8xx6 = (Pg6xx6 | P87xx6);
assign Qb8xx6 = (Gf6xx6 | R97xx6);
assign Ql5xx6 = (~(Ec8xx6 & Lc8xx6));
assign Lc8xx6 = (Sc8xx6 & Zc8xx6);
assign Zc8xx6 = (Gf6xx6 | Hb7xx6);
assign Sc8xx6 = (Pg6xx6 | Cc7xx6);
assign Ec8xx6 = (Gd8xx6 & Nd8xx6);
assign Nd8xx6 = (Vj6xx6 | K97xx6);
assign Gd8xx6 = (Hj6xx6 | Jc7xx6);
assign Vdt7v6 = (Zr7xx6 ? Ud8xx6 : V10nz6[6]);
assign Odt7v6 = (Gs7xx6 ? Ud8xx6 : F00nz6[6]);
assign Hdt7v6 = (Ns7xx6 ? Ud8xx6 : Pyzmz6[6]);
assign Ud8xx6 = (R21nz6[2] ? Em5xx6 : Lm5xx6);
assign Em5xx6 = (~(Be8xx6 & Ie8xx6));
assign Ie8xx6 = (Pe8xx6 & We8xx6);
assign We8xx6 = (~(Zd7xx6 & Df8xx6));
assign Pe8xx6 = (Ne7xx6 | Hj6xx6);
assign Be8xx6 = (Kf8xx6 & Rf8xx6);
assign Rf8xx6 = (Vj6xx6 | Yg7xx6);
assign Kf8xx6 = (Gf6xx6 | Pf7xx6);
assign Lm5xx6 = (~(Yf8xx6 & Fg8xx6));
assign Fg8xx6 = (Mg8xx6 & Tg8xx6);
assign Tg8xx6 = (Gf6xx6 | Fh7xx6);
assign Mg8xx6 = (Pg6xx6 | Ai7xx6);
assign Yf8xx6 = (Ah8xx6 & Hh8xx6);
assign Hh8xx6 = (Vj6xx6 | If7xx6);
assign Ah8xx6 = (Hj6xx6 | Hi7xx6);
assign Adt7v6 = (Zr7xx6 ? Oh8xx6 : V10nz6[7]);
assign Zr7xx6 = (Vh8xx6 & Ci8xx6);
assign Tct7v6 = (Gs7xx6 ? Oh8xx6 : F00nz6[7]);
assign Gs7xx6 = (Vh8xx6 & Ji8xx6);
assign Vh8xx6 = (Qi8xx6 & Xi8xx6);
assign Qi8xx6 = (!Ej8xx6);
assign Mct7v6 = (Ns7xx6 ? Oh8xx6 : Pyzmz6[7]);
assign Ns7xx6 = (Lj8xx6 & Ej8xx6);
assign Ej8xx6 = (Sj8xx6 ? Fc5xx6 : B41nz6[1]);
assign Lj8xx6 = (Ci8xx6 & Xi8xx6);
assign Xi8xx6 = (~(Zj8xx6 & Gk8xx6));
assign Gk8xx6 = (~(Nk8xx6 & Vc6xx6));
assign Nk8xx6 = (Gha7z6 & Uk8xx6);
assign Uk8xx6 = (~(Sj8xx6 & B35xx6));
assign Zj8xx6 = (~(Ce5xx6 & Pm7xx6));
assign Pm7xx6 = (!Sj8xx6);
assign Ci8xx6 = (!Ji8xx6);
assign Ji8xx6 = (Sj8xx6 ? Ef5xx6 : B41nz6[0]);
assign Oh8xx6 = (R21nz6[2] ? Tq5xx6 : Ar5xx6);
assign Tq5xx6 = (~(Bl8xx6 & Il8xx6));
assign Il8xx6 = (Pl8xx6 & Wl8xx6);
assign Wl8xx6 = (~(Dm8xx6 & Ge7xx6));
assign Pl8xx6 = (Vj6xx6 | Cq7xx6);
assign Bl8xx6 = (Km8xx6 & Rm8xx6);
assign Rm8xx6 = (~(Df8xx6 & Ym8xx6));
assign Km8xx6 = (Gf6xx6 | Rn7xx6);
assign Ar5xx6 = (~(Fn8xx6 & Mn8xx6));
assign Mn8xx6 = (Tn8xx6 & Ao8xx6);
assign Ao8xx6 = (Gf6xx6 | Jq7xx6);
assign Tn8xx6 = (Pg6xx6 | Er7xx6);
assign Fn8xx6 = (Ho8xx6 & Oo8xx6);
assign Oo8xx6 = (Vj6xx6 | To7xx6);
assign Ho8xx6 = (Hj6xx6 | Lr7xx6);
assign Fct7v6 = (Cp8xx6 ? Vo8xx6 : Zwzmz6[0]);
assign Ybt7v6 = (Jp8xx6 ? Vo8xx6 : Jvzmz6[0]);
assign Rbt7v6 = (Qp8xx6 ? Vo8xx6 : Ttzmz6[0]);
assign Vo8xx6 = (R21nz6[2] ? Js5xx6 : Qs5xx6);
assign Js5xx6 = (~(Xp8xx6 & Eq8xx6));
assign Eq8xx6 = (Hj6xx6 | Mi6xx6);
assign Xp8xx6 = (Lq8xx6 & Sq8xx6);
assign Sq8xx6 = (Du7xx6 | Ig6xx6);
assign Ig6xx6 = (R21nz6[0] ? Gr8xx6 : Zq8xx6);
assign Zq8xx6 = (!It7xx6);
assign Lq8xx6 = (Vj6xx6 | Fi6xx6);
assign Qs5xx6 = (~(Nr8xx6 & Ur8xx6));
assign Ur8xx6 = (Bs8xx6 & Is8xx6);
assign Is8xx6 = (Gf6xx6 | Oj6xx6);
assign Bs8xx6 = (Pg6xx6 | Ck6xx6);
assign Nr8xx6 = (Ps8xx6 & Ws8xx6);
assign Ws8xx6 = (Vj6xx6 | Wg6xx6);
assign Ps8xx6 = (Hj6xx6 | Nf6xx6);
assign Kbt7v6 = (Cp8xx6 ? Dt8xx6 : Zwzmz6[1]);
assign Dbt7v6 = (Jp8xx6 ? Dt8xx6 : Jvzmz6[1]);
assign Wat7v6 = (Qp8xx6 ? Dt8xx6 : Ttzmz6[1]);
assign Dt8xx6 = (R21nz6[2] ? Et5xx6 : Lt5xx6);
assign Et5xx6 = (~(Kt8xx6 & Rt8xx6));
assign Rt8xx6 = (Yt8xx6 & Fu8xx6);
assign Fu8xx6 = (Sl6xx6 | Pg6xx6);
assign Yt8xx6 = (Hj6xx6 | Ko6xx6);
assign Kt8xx6 = (Mu8xx6 & Tu8xx6);
assign Tu8xx6 = (Vj6xx6 | Ro6xx6);
assign Mu8xx6 = (Gf6xx6 | Bn6xx6);
assign Lt5xx6 = (~(Av8xx6 & Hv8xx6));
assign Hv8xx6 = (Ov8xx6 & Vv8xx6);
assign Vv8xx6 = (Gf6xx6 | Mp6xx6);
assign Ov8xx6 = (Hj6xx6 | Zl6xx6);
assign Av8xx6 = (Cw8xx6 & Jw8xx6);
assign Jw8xx6 = (Vj6xx6 | Um6xx6);
assign Cw8xx6 = (Pg6xx6 | Tp6xx6);
assign Pat7v6 = (Cp8xx6 ? Qw8xx6 : Zwzmz6[2]);
assign Iat7v6 = (Jp8xx6 ? Qw8xx6 : Jvzmz6[2]);
assign Bat7v6 = (Qp8xx6 ? Qw8xx6 : Ttzmz6[2]);
assign Qw8xx6 = (R21nz6[2] ? Zt5xx6 : Gu5xx6);
assign Zt5xx6 = (~(Xw8xx6 & Ex8xx6));
assign Ex8xx6 = (Lx8xx6 & Sx8xx6);
assign Sx8xx6 = (Pg6xx6 | Jr6xx6);
assign Lx8xx6 = (Hj6xx6 | Bu6xx6);
assign Xw8xx6 = (Zx8xx6 & Gy8xx6);
assign Gy8xx6 = (Vj6xx6 | Iu6xx6);
assign Zx8xx6 = (Gf6xx6 | Ss6xx6);
assign Gu5xx6 = (~(Ny8xx6 & Uy8xx6));
assign Uy8xx6 = (Bz8xx6 & Iz8xx6);
assign Iz8xx6 = (Gf6xx6 | Dv6xx6);
assign Bz8xx6 = (Hj6xx6 | Qr6xx6);
assign Ny8xx6 = (Pz8xx6 & Wz8xx6);
assign Wz8xx6 = (Vj6xx6 | Ls6xx6);
assign Pz8xx6 = (Pg6xx6 | Kv6xx6);
assign U9t7v6 = (Cp8xx6 ? D09xx6 : Zwzmz6[3]);
assign N9t7v6 = (Jp8xx6 ? D09xx6 : Jvzmz6[3]);
assign G9t7v6 = (Qp8xx6 ? D09xx6 : Ttzmz6[3]);
assign D09xx6 = (R21nz6[2] ? Uu5xx6 : Bv5xx6);
assign Uu5xx6 = (~(K09xx6 & R09xx6));
assign R09xx6 = (Y09xx6 & F19xx6);
assign F19xx6 = (Pg6xx6 | Ax6xx6);
assign Y09xx6 = (Hj6xx6 | Sz6xx6);
assign K09xx6 = (M19xx6 & T19xx6);
assign T19xx6 = (Vj6xx6 | Zz6xx6);
assign M19xx6 = (Gf6xx6 | Hx6xx6);
assign Bv5xx6 = (~(A29xx6 & H29xx6));
assign H29xx6 = (O29xx6 & V29xx6);
assign V29xx6 = (Gf6xx6 | U07xx6);
assign O29xx6 = (Hj6xx6 | Cy6xx6);
assign A29xx6 = (C39xx6 & J39xx6);
assign J39xx6 = (Vj6xx6 | Jy6xx6);
assign C39xx6 = (Pg6xx6 | B17xx6);
assign Z8t7v6 = (Cp8xx6 ? Q39xx6 : Zwzmz6[4]);
assign S8t7v6 = (Jp8xx6 ? Q39xx6 : Jvzmz6[4]);
assign L8t7v6 = (Qp8xx6 ? Q39xx6 : Ttzmz6[4]);
assign Q39xx6 = (R21nz6[2] ? Pv5xx6 : Wv5xx6);
assign Pv5xx6 = (~(X39xx6 & E49xx6));
assign E49xx6 = (L49xx6 & S49xx6);
assign S49xx6 = (Pg6xx6 | R27xx6);
assign L49xx6 = (Hj6xx6 | J57xx6);
assign X39xx6 = (Z49xx6 & G59xx6);
assign G59xx6 = (Vj6xx6 | Q57xx6);
assign Z49xx6 = (Gf6xx6 | Y27xx6);
assign Wv5xx6 = (~(N59xx6 & U59xx6));
assign U59xx6 = (B69xx6 & I69xx6);
assign I69xx6 = (Gf6xx6 | L67xx6);
assign B69xx6 = (Hj6xx6 | T37xx6);
assign N59xx6 = (P69xx6 & W69xx6);
assign W69xx6 = (Vj6xx6 | A47xx6);
assign P69xx6 = (Pg6xx6 | S67xx6);
assign E8t7v6 = (Cp8xx6 ? D79xx6 : Zwzmz6[5]);
assign X7t7v6 = (Jp8xx6 ? D79xx6 : Jvzmz6[5]);
assign Q7t7v6 = (Qp8xx6 ? D79xx6 : Ttzmz6[5]);
assign D79xx6 = (R21nz6[2] ? Kw5xx6 : Rw5xx6);
assign Kw5xx6 = (~(K79xx6 & R79xx6));
assign R79xx6 = (Y79xx6 & F89xx6);
assign F89xx6 = (Pg6xx6 | I87xx6);
assign Y79xx6 = (Hj6xx6 | Ab7xx6);
assign K79xx6 = (M89xx6 & T89xx6);
assign T89xx6 = (Vj6xx6 | Hb7xx6);
assign M89xx6 = (Gf6xx6 | P87xx6);
assign Rw5xx6 = (~(A99xx6 & H99xx6));
assign H99xx6 = (O99xx6 & V99xx6);
assign V99xx6 = (Gf6xx6 | Cc7xx6);
assign O99xx6 = (Hj6xx6 | K97xx6);
assign A99xx6 = (Ca9xx6 & Ja9xx6);
assign Ja9xx6 = (Vj6xx6 | R97xx6);
assign Ca9xx6 = (Pg6xx6 | Jc7xx6);
assign J7t7v6 = (Cp8xx6 ? Qa9xx6 : Zwzmz6[6]);
assign C7t7v6 = (Jp8xx6 ? Qa9xx6 : Jvzmz6[6]);
assign V6t7v6 = (Qp8xx6 ? Qa9xx6 : Ttzmz6[6]);
assign Qa9xx6 = (R21nz6[2] ? Fx5xx6 : Mx5xx6);
assign Fx5xx6 = (~(Xa9xx6 & Eb9xx6));
assign Eb9xx6 = (Lb9xx6 & Sb9xx6);
assign Sb9xx6 = (~(Zd7xx6 & Zb9xx6));
assign Lb9xx6 = (Ne7xx6 | Pg6xx6);
assign Xa9xx6 = (Gc9xx6 & Nc9xx6);
assign Nc9xx6 = (Hj6xx6 | Yg7xx6);
assign Gc9xx6 = (Vj6xx6 | Fh7xx6);
assign Mx5xx6 = (~(Uc9xx6 & Bd9xx6));
assign Bd9xx6 = (Id9xx6 & Pd9xx6);
assign Pd9xx6 = (Gf6xx6 | Ai7xx6);
assign Id9xx6 = (Hj6xx6 | If7xx6);
assign Uc9xx6 = (Wd9xx6 & De9xx6);
assign De9xx6 = (Vj6xx6 | Pf7xx6);
assign Wd9xx6 = (Pg6xx6 | Hi7xx6);
assign O6t7v6 = (Cp8xx6 ? Ke9xx6 : Zwzmz6[7]);
assign Cp8xx6 = (Re9xx6 & Ye9xx6);
assign H6t7v6 = (Jp8xx6 ? Ke9xx6 : Jvzmz6[7]);
assign Jp8xx6 = (Re9xx6 & Ff9xx6);
assign Re9xx6 = (Mf9xx6 & Tf9xx6);
assign Mf9xx6 = (!Ag9xx6);
assign A6t7v6 = (Qp8xx6 ? Ke9xx6 : Ttzmz6[7]);
assign Qp8xx6 = (Hg9xx6 & Ag9xx6);
assign Ag9xx6 = (Og9xx6 ? Fc5xx6 : B41nz6[1]);
assign Hg9xx6 = (Ye9xx6 & Tf9xx6);
assign Tf9xx6 = (~(Vg9xx6 & Ch9xx6));
assign Ch9xx6 = (~(Jh9xx6 & Qh9xx6));
assign Qh9xx6 = (Oha7z6 & Xh9xx6);
assign Xh9xx6 = (~(Og9xx6 & B35xx6));
assign Oha7z6 = (~(Ei9xx6 | Li9xx6));
assign Li9xx6 = (~(Wsc7v6 | T51nz6[0]));
assign Jh9xx6 = (Gha7z6 & Vc6xx6);
assign Vc6xx6 = (Mho7v6 & Fftnv6);
assign Gha7z6 = (Si9xx6 ^ Ei9xx6);
assign Si9xx6 = (Zi9xx6 ^ P26xx6);
assign Vg9xx6 = (~(Ce5xx6 & Gj9xx6));
assign Gj9xx6 = (!Og9xx6);
assign Ye9xx6 = (!Ff9xx6);
assign Ff9xx6 = (Og9xx6 ? Ef5xx6 : B41nz6[0]);
assign Og9xx6 = (Sj8xx6 & T51nz6[0]);
assign Sj8xx6 = (T51nz6[2] & T51nz6[1]);
assign Ke9xx6 = (R21nz6[2] ? K36xx6 : R36xx6);
assign K36xx6 = (~(Nj9xx6 & Uj9xx6));
assign Uj9xx6 = (Vj6xx6 | Jq7xx6);
assign Nj9xx6 = (Bk9xx6 & Ik9xx6);
assign Ik9xx6 = (Du7xx6 | Mo7xx6);
assign Mo7xx6 = (Pk9xx6 & Wk9xx6);
assign Wk9xx6 = (~(Dl9xx6 & Kl9xx6));
assign Pk9xx6 = (~(R21nz6[0] & Ym8xx6));
assign Bk9xx6 = (Hj6xx6 | Cq7xx6);
assign R36xx6 = (~(Rl9xx6 & Yl9xx6));
assign Yl9xx6 = (Fm9xx6 & Mm9xx6);
assign Mm9xx6 = (Gf6xx6 | Er7xx6);
assign Fm9xx6 = (Hj6xx6 | To7xx6);
assign Rl9xx6 = (Tm9xx6 & An9xx6);
assign An9xx6 = (Pg6xx6 | Lr7xx6);
assign Tm9xx6 = (Vj6xx6 | Rn7xx6);
assign T5t7v6 = (I35xx6 ? Dszmz6[0] : Hn9xx6);
assign M5t7v6 = (N25xx6 ? Nqzmz6[0] : Hn9xx6);
assign F5t7v6 = (On9xx6 ? Hn9xx6 : Xozmz6[0]);
assign Hn9xx6 = (R21nz6[2] ? A56xx6 : H56xx6);
assign A56xx6 = (~(Vn9xx6 & Co9xx6));
assign Co9xx6 = (Jo9xx6 & Qo9xx6);
assign Qo9xx6 = (Hj6xx6 | Fi6xx6);
assign Fi6xx6 = (Xo9xx6 & Ep9xx6);
assign Ep9xx6 = (~(Gnzmz6[8] & Lp9xx6));
assign Xo9xx6 = (Sp9xx6 & Zp9xx6);
assign Sp9xx6 = (~(Gq9xx6 & Jezmz6[16]));
assign Gq9xx6 = (Dl9xx6 & Nq9xx6);
assign Jo9xx6 = (Pg6xx6 | Mi6xx6);
assign Mi6xx6 = (Uq9xx6 & Br9xx6);
assign Br9xx6 = (~(Gnzmz6[0] & Lp9xx6));
assign Uq9xx6 = (Ir9xx6 & Zp9xx6);
assign Ir9xx6 = (~(Jezmz6[8] & Pr9xx6));
assign Vn9xx6 = (Wr9xx6 & Ds9xx6);
assign Ds9xx6 = (Vj6xx6 | Oj6xx6);
assign Oj6xx6 = (Ks9xx6 & Rs9xx6);
assign Rs9xx6 = (Ys9xx6 & Ft9xx6);
assign Ft9xx6 = (~(Jezmz6[8] & Mt9xx6));
assign Ys9xx6 = (~(Tt9xx6 & Jezmz6[24]));
assign Tt9xx6 = (Dl9xx6 & Au9xx6);
assign Ks9xx6 = (Hu9xx6 & Ou9xx6);
assign Ou9xx6 = (~(Vu9xx6 & Cv9xx6));
assign Hu9xx6 = (~(Gnzmz6[16] & Lp9xx6));
assign Wr9xx6 = (~(Zb9xx6 & It7xx6));
assign H56xx6 = (~(Jv9xx6 & Qv9xx6));
assign Qv9xx6 = (Pg6xx6 | Nf6xx6);
assign Nf6xx6 = (Xv9xx6 & Ew9xx6);
assign Ew9xx6 = (~(Jezmz6[24] & Mt9xx6));
assign Xv9xx6 = (Lw9xx6 & Sw9xx6);
assign Sw9xx6 = (~(Zw9xx6 & Cv9xx6));
assign Lw9xx6 = (~(Gnzmz6[32] & Lp9xx6));
assign Jv9xx6 = (Gx9xx6 & Nx9xx6);
assign Nx9xx6 = (Gf6xx6 | Ck6xx6);
assign Ck6xx6 = (Ux9xx6 & By9xx6);
assign By9xx6 = (Iy9xx6 & Py9xx6);
assign Py9xx6 = (~(Jezmz6[16] & Mt9xx6));
assign Iy9xx6 = (~(Wy9xx6 & Jezmz6[32]));
assign Wy9xx6 = (Dl9xx6 & Dz9xx6);
assign Ux9xx6 = (Kz9xx6 & Rz9xx6);
assign Rz9xx6 = (~(Yz9xx6 & Cv9xx6));
assign Kz9xx6 = (~(Gnzmz6[24] & Lp9xx6));
assign Gx9xx6 = (Ku7xx6 | R21nz6[1]);
assign Ku7xx6 = (R21nz6[0] ? Wg6xx6 : Gr8xx6);
assign Wg6xx6 = (F0axx6 & M0axx6);
assign M0axx6 = (~(T0axx6 & Cv9xx6));
assign Cv9xx6 = (Pazmz6[4] & Dl9xx6);
assign F0axx6 = (~(Gnzmz6[40] & Lp9xx6));
assign Gr8xx6 = (~(Cfc7v6 & Lp9xx6));
assign Y4t7v6 = (I35xx6 ? Dszmz6[1] : A1axx6);
assign R4t7v6 = (N25xx6 ? Nqzmz6[1] : A1axx6);
assign K4t7v6 = (On9xx6 ? A1axx6 : Xozmz6[1]);
assign A1axx6 = (R21nz6[2] ? V56xx6 : C66xx6);
assign V56xx6 = (~(H1axx6 & O1axx6));
assign O1axx6 = (V1axx6 & C2axx6);
assign C2axx6 = (Sl6xx6 | Gf6xx6);
assign Sl6xx6 = (~(J2axx6 & Q2axx6));
assign Q2axx6 = (~(X2axx6 & E3axx6));
assign E3axx6 = (~(Dl9xx6 & L3axx6));
assign L3axx6 = (S3axx6 | Jezmz6[1]);
assign S3axx6 = (~(Ro87v6 | Z3axx6));
assign J2axx6 = (G4axx6 | N4axx6);
assign V1axx6 = (Pg6xx6 | Ko6xx6);
assign Ko6xx6 = (U4axx6 & B5axx6);
assign B5axx6 = (~(Gnzmz6[1] & Lp9xx6));
assign U4axx6 = (~(I5axx6 | P5axx6));
assign I5axx6 = (W5axx6 & Dl9xx6);
assign W5axx6 = (D6axx6 & K6axx6);
assign K6axx6 = (R6axx6 | Jezmz6[9]);
assign R6axx6 = (~(Y6axx6 | Z3axx6));
assign D6axx6 = (~(Z3axx6 & F7axx6));
assign H1axx6 = (M7axx6 & T7axx6);
assign T7axx6 = (Hj6xx6 | Ro6xx6);
assign Ro6xx6 = (A8axx6 & H8axx6);
assign H8axx6 = (~(Dl9xx6 & O8axx6));
assign O8axx6 = (~(V8axx6 & C9axx6));
assign C9axx6 = (~(Pazmz6[0] & J9axx6));
assign V8axx6 = (Q9axx6 & X9axx6);
assign X9axx6 = (Z3axx6 | Eaaxx6);
assign Q9axx6 = (~(Jezmz6[17] & Nq9xx6));
assign A8axx6 = (Laaxx6 & Saaxx6);
assign Saaxx6 = (~(Zaaxx6 & Gbaxx6));
assign Gbaxx6 = (P5axx6 | Gnzmz6[9]);
assign Laaxx6 = (~(Jezmz6[1] & Mt9xx6));
assign M7axx6 = (Vj6xx6 | Mp6xx6);
assign Mp6xx6 = (Nbaxx6 & Ubaxx6);
assign Ubaxx6 = (~(Dl9xx6 & Bcaxx6));
assign Bcaxx6 = (~(Icaxx6 & Pcaxx6));
assign Pcaxx6 = (Wcaxx6 & Ddaxx6);
assign Ddaxx6 = (Kdaxx6 | Z3axx6);
assign Wcaxx6 = (~(Jezmz6[25] & Au9xx6));
assign Icaxx6 = (Rdaxx6 & Ydaxx6);
assign Ydaxx6 = (~(Pazmz6[0] & Feaxx6));
assign Rdaxx6 = (~(Pazmz6[5] & Vu9xx6));
assign Nbaxx6 = (Meaxx6 & Teaxx6);
assign Teaxx6 = (~(Zaaxx6 & Afaxx6));
assign Afaxx6 = (P5axx6 | Gnzmz6[17]);
assign Meaxx6 = (~(Jezmz6[9] & Mt9xx6));
assign C66xx6 = (~(Hfaxx6 & Ofaxx6));
assign Ofaxx6 = (Vfaxx6 & Cgaxx6);
assign Cgaxx6 = (Pg6xx6 | Zl6xx6);
assign Zl6xx6 = (Jgaxx6 & Qgaxx6);
assign Qgaxx6 = (~(Dl9xx6 & Xgaxx6));
assign Xgaxx6 = (~(Ehaxx6 & Lhaxx6));
assign Lhaxx6 = (~(Pazmz6[5] & Zw9xx6));
assign Ehaxx6 = (Shaxx6 & Zhaxx6);
assign Zhaxx6 = (Z3axx6 | Giaxx6);
assign Shaxx6 = (~(Pazmz6[0] & Niaxx6));
assign Jgaxx6 = (Uiaxx6 & Bjaxx6);
assign Bjaxx6 = (~(Zaaxx6 & Ijaxx6));
assign Ijaxx6 = (P5axx6 | Gnzmz6[33]);
assign Uiaxx6 = (~(Jezmz6[25] & Mt9xx6));
assign Vfaxx6 = (Hj6xx6 | Um6xx6);
assign Um6xx6 = (Pjaxx6 & Wjaxx6);
assign Wjaxx6 = (Dkaxx6 & Kkaxx6);
assign Dkaxx6 = (~(Gnzmz6[41] & Lp9xx6));
assign Pjaxx6 = (Rkaxx6 & Ykaxx6);
assign Ykaxx6 = (Flaxx6 | Z3axx6);
assign Rkaxx6 = (~(Mlaxx6 & Dl9xx6));
assign Mlaxx6 = (Tlaxx6 & Amaxx6);
assign Amaxx6 = (~(Hmaxx6 & Omaxx6));
assign Omaxx6 = (!Pazmz6[5]);
assign Hmaxx6 = (Vmaxx6 | Z3axx6);
assign Tlaxx6 = (~(Z3axx6 & Cnaxx6));
assign Hfaxx6 = (Jnaxx6 & Qnaxx6);
assign Qnaxx6 = (Vj6xx6 | Bn6xx6);
assign Bn6xx6 = (Xnaxx6 & Eoaxx6);
assign Eoaxx6 = (~(Ym8xx6 & G4axx6));
assign Xnaxx6 = (~(Wgc7v6 & Lp9xx6));
assign Jnaxx6 = (Gf6xx6 | Tp6xx6);
assign Tp6xx6 = (Loaxx6 & Soaxx6);
assign Soaxx6 = (~(Dl9xx6 & Zoaxx6));
assign Zoaxx6 = (~(Gpaxx6 & Npaxx6));
assign Npaxx6 = (Upaxx6 & Bqaxx6);
assign Bqaxx6 = (~(G4axx6 & Iqaxx6));
assign Upaxx6 = (~(Pazmz6[5] & Yz9xx6));
assign Gpaxx6 = (Pqaxx6 & Wqaxx6);
assign Wqaxx6 = (~(Pazmz6[0] & Draxx6));
assign Pqaxx6 = (~(Jezmz6[33] & Dz9xx6));
assign Loaxx6 = (Kraxx6 & Rraxx6);
assign Rraxx6 = (~(Zaaxx6 & Yraxx6));
assign Yraxx6 = (P5axx6 | Gnzmz6[25]);
assign Zaaxx6 = (P5axx6 | Lp9xx6);
assign P5axx6 = (Fsaxx6 & G4axx6);
assign G4axx6 = (!Z3axx6);
assign Kraxx6 = (~(Jezmz6[17] & Mt9xx6));
assign D4t7v6 = (I35xx6 ? Dszmz6[2] : Msaxx6);
assign W3t7v6 = (N25xx6 ? Nqzmz6[2] : Msaxx6);
assign P3t7v6 = (On9xx6 ? Msaxx6 : Xozmz6[2]);
assign Msaxx6 = (R21nz6[2] ? Q66xx6 : X66xx6);
assign Q66xx6 = (~(Tsaxx6 & Ataxx6));
assign Ataxx6 = (Htaxx6 & Otaxx6);
assign Otaxx6 = (Gf6xx6 | Jr6xx6);
assign Jr6xx6 = (Vtaxx6 & Cuaxx6);
assign Vtaxx6 = (~(Juaxx6 & Dl9xx6));
assign Juaxx6 = (Quaxx6 & Xuaxx6);
assign Xuaxx6 = (~(Evaxx6 & Lvaxx6));
assign Lvaxx6 = (~(Jezmz6[2] & Svaxx6));
assign Svaxx6 = (~(F7axx6 & Zvaxx6));
assign Quaxx6 = (Zvaxx6 | Jezmz6[2]);
assign Htaxx6 = (Pg6xx6 | Bu6xx6);
assign Bu6xx6 = (Gwaxx6 & Nwaxx6);
assign Nwaxx6 = (~(Gnzmz6[2] & Lp9xx6));
assign Gwaxx6 = (~(Uwaxx6 | Bxaxx6));
assign Uwaxx6 = (Ixaxx6 & Dl9xx6);
assign Ixaxx6 = (Pxaxx6 & Wxaxx6);
assign Wxaxx6 = (Dyaxx6 | Jezmz6[10]);
assign Dyaxx6 = (~(Y6axx6 | Evaxx6));
assign Pxaxx6 = (~(Evaxx6 & F7axx6));
assign Tsaxx6 = (Kyaxx6 & Ryaxx6);
assign Ryaxx6 = (Hj6xx6 | Iu6xx6);
assign Iu6xx6 = (Yyaxx6 & Fzaxx6);
assign Fzaxx6 = (~(Dl9xx6 & Mzaxx6));
assign Mzaxx6 = (~(Tzaxx6 & A0bxx6));
assign A0bxx6 = (~(Pazmz6[1] & J9axx6));
assign Tzaxx6 = (H0bxx6 & O0bxx6);
assign O0bxx6 = (Evaxx6 | Eaaxx6);
assign H0bxx6 = (~(Jezmz6[18] & Nq9xx6));
assign Yyaxx6 = (V0bxx6 & C1bxx6);
assign C1bxx6 = (~(J1bxx6 & Q1bxx6));
assign Q1bxx6 = (Bxaxx6 | Gnzmz6[10]);
assign V0bxx6 = (~(Jezmz6[2] & Mt9xx6));
assign Kyaxx6 = (Vj6xx6 | Dv6xx6);
assign Dv6xx6 = (X1bxx6 & E2bxx6);
assign E2bxx6 = (~(Dl9xx6 & L2bxx6));
assign L2bxx6 = (~(S2bxx6 & Z2bxx6));
assign Z2bxx6 = (G3bxx6 & N3bxx6);
assign N3bxx6 = (Kdaxx6 | Evaxx6);
assign G3bxx6 = (~(Jezmz6[26] & Au9xx6));
assign S2bxx6 = (U3bxx6 & B4bxx6);
assign B4bxx6 = (~(Pazmz6[1] & Feaxx6));
assign U3bxx6 = (~(Pazmz6[6] & Vu9xx6));
assign X1bxx6 = (I4bxx6 & P4bxx6);
assign P4bxx6 = (~(J1bxx6 & W4bxx6));
assign W4bxx6 = (Bxaxx6 | Gnzmz6[18]);
assign I4bxx6 = (~(Jezmz6[10] & Mt9xx6));
assign X66xx6 = (~(D5bxx6 & K5bxx6));
assign K5bxx6 = (R5bxx6 & Y5bxx6);
assign Y5bxx6 = (Pg6xx6 | Qr6xx6);
assign Qr6xx6 = (F6bxx6 & M6bxx6);
assign M6bxx6 = (~(Dl9xx6 & T6bxx6));
assign T6bxx6 = (~(A7bxx6 & H7bxx6));
assign H7bxx6 = (~(Pazmz6[6] & Zw9xx6));
assign A7bxx6 = (O7bxx6 & V7bxx6);
assign V7bxx6 = (Evaxx6 | Giaxx6);
assign O7bxx6 = (~(Pazmz6[1] & Niaxx6));
assign F6bxx6 = (C8bxx6 & J8bxx6);
assign J8bxx6 = (~(J1bxx6 & Q8bxx6));
assign Q8bxx6 = (Bxaxx6 | Gnzmz6[34]);
assign C8bxx6 = (~(Jezmz6[26] & Mt9xx6));
assign R5bxx6 = (Hj6xx6 | Ls6xx6);
assign Ls6xx6 = (X8bxx6 & E9bxx6);
assign E9bxx6 = (L9bxx6 & Kkaxx6);
assign L9bxx6 = (~(Gnzmz6[42] & Lp9xx6));
assign X8bxx6 = (S9bxx6 & Z9bxx6);
assign Z9bxx6 = (Flaxx6 | Evaxx6);
assign S9bxx6 = (~(Gabxx6 & Dl9xx6));
assign Gabxx6 = (Nabxx6 & Uabxx6);
assign Uabxx6 = (~(Bbbxx6 & Ibbxx6));
assign Bbbxx6 = (Vmaxx6 | Evaxx6);
assign Nabxx6 = (~(Evaxx6 & Cnaxx6));
assign Evaxx6 = (!Pbbxx6);
assign D5bxx6 = (Wbbxx6 & Dcbxx6);
assign Dcbxx6 = (Vj6xx6 | Ss6xx6);
assign Ss6xx6 = (Kcbxx6 & Rcbxx6);
assign Rcbxx6 = (~(Ym8xx6 & Pbbxx6));
assign Kcbxx6 = (~(Qic7v6 & Lp9xx6));
assign Wbbxx6 = (Gf6xx6 | Kv6xx6);
assign Kv6xx6 = (Ycbxx6 & Fdbxx6);
assign Fdbxx6 = (~(Dl9xx6 & Mdbxx6));
assign Mdbxx6 = (~(Tdbxx6 & Aebxx6));
assign Aebxx6 = (Hebxx6 & Oebxx6);
assign Oebxx6 = (~(Pbbxx6 & Iqaxx6));
assign Hebxx6 = (~(Pazmz6[6] & Yz9xx6));
assign Tdbxx6 = (Vebxx6 & Cfbxx6);
assign Cfbxx6 = (~(Pazmz6[1] & Draxx6));
assign Vebxx6 = (~(Jezmz6[34] & Dz9xx6));
assign Ycbxx6 = (Jfbxx6 & Qfbxx6);
assign Qfbxx6 = (~(J1bxx6 & Xfbxx6));
assign Xfbxx6 = (Bxaxx6 | Gnzmz6[26]);
assign J1bxx6 = (Bxaxx6 | Lp9xx6);
assign Bxaxx6 = (Fsaxx6 & Pbbxx6);
assign Pbbxx6 = (~(Egbxx6 & Lgbxx6));
assign Egbxx6 = (~(Lczmz6[0] & Sgbxx6));
assign Jfbxx6 = (~(Jezmz6[18] & Mt9xx6));
assign I3t7v6 = (I35xx6 ? Dszmz6[3] : Zgbxx6);
assign B3t7v6 = (N25xx6 ? Nqzmz6[3] : Zgbxx6);
assign U2t7v6 = (On9xx6 ? Zgbxx6 : Xozmz6[3]);
assign Zgbxx6 = (R21nz6[2] ? L76xx6 : S76xx6);
assign L76xx6 = (~(Ghbxx6 & Nhbxx6));
assign Nhbxx6 = (Uhbxx6 & Bibxx6);
assign Bibxx6 = (Gf6xx6 | Ax6xx6);
assign Ax6xx6 = (Iibxx6 & Pibxx6);
assign Pibxx6 = (~(Wibxx6 & Djbxx6));
assign Iibxx6 = (Kjbxx6 & Zp9xx6);
assign Kjbxx6 = (~(Jezmz6[3] & It7xx6));
assign Uhbxx6 = (Pg6xx6 | Sz6xx6);
assign Sz6xx6 = (Rjbxx6 & Yjbxx6);
assign Yjbxx6 = (~(Fkbxx6 | Mkbxx6));
assign Fkbxx6 = (Jezmz6[11] & Pr9xx6);
assign Rjbxx6 = (Tkbxx6 & Albxx6);
assign Albxx6 = (~(Gnzmz6[3] & Lp9xx6));
assign Tkbxx6 = (~(Hlbxx6 & Djbxx6));
assign Ghbxx6 = (Olbxx6 & Vlbxx6);
assign Vlbxx6 = (Hj6xx6 | Zz6xx6);
assign Zz6xx6 = (Cmbxx6 & Jmbxx6);
assign Jmbxx6 = (~(Dl9xx6 & Qmbxx6));
assign Qmbxx6 = (~(Xmbxx6 & Enbxx6));
assign Enbxx6 = (~(Pazmz6[2] & J9axx6));
assign Xmbxx6 = (Lnbxx6 & Snbxx6);
assign Snbxx6 = (Znbxx6 | Eaaxx6);
assign Lnbxx6 = (~(Jezmz6[19] & Nq9xx6));
assign Cmbxx6 = (Gobxx6 & Nobxx6);
assign Nobxx6 = (~(Uobxx6 & Bpbxx6));
assign Bpbxx6 = (Mkbxx6 | Gnzmz6[11]);
assign Gobxx6 = (~(Jezmz6[3] & Mt9xx6));
assign Olbxx6 = (Vj6xx6 | U07xx6);
assign U07xx6 = (Ipbxx6 & Ppbxx6);
assign Ppbxx6 = (~(Dl9xx6 & Wpbxx6));
assign Wpbxx6 = (~(Dqbxx6 & Kqbxx6));
assign Kqbxx6 = (Rqbxx6 & Yqbxx6);
assign Yqbxx6 = (Kdaxx6 | Znbxx6);
assign Rqbxx6 = (~(Jezmz6[27] & Au9xx6));
assign Dqbxx6 = (Frbxx6 & Mrbxx6);
assign Mrbxx6 = (~(Pazmz6[2] & Feaxx6));
assign Frbxx6 = (~(Pazmz6[7] & Vu9xx6));
assign Ipbxx6 = (Trbxx6 & Asbxx6);
assign Asbxx6 = (~(Uobxx6 & Hsbxx6));
assign Hsbxx6 = (Mkbxx6 | Gnzmz6[19]);
assign Trbxx6 = (~(Jezmz6[11] & Mt9xx6));
assign S76xx6 = (~(Osbxx6 & Vsbxx6));
assign Vsbxx6 = (Ctbxx6 & Jtbxx6);
assign Jtbxx6 = (Vj6xx6 | Hx6xx6);
assign Hx6xx6 = (Qtbxx6 & Xtbxx6);
assign Xtbxx6 = (~(Ym8xx6 & Djbxx6));
assign Qtbxx6 = (~(Kkc7v6 & Lp9xx6));
assign Ctbxx6 = (Pg6xx6 | Cy6xx6);
assign Cy6xx6 = (Eubxx6 & Lubxx6);
assign Lubxx6 = (~(Dl9xx6 & Subxx6));
assign Subxx6 = (~(Zubxx6 & Gvbxx6));
assign Gvbxx6 = (~(Pazmz6[7] & Zw9xx6));
assign Zubxx6 = (Nvbxx6 & Uvbxx6);
assign Uvbxx6 = (Znbxx6 | Giaxx6);
assign Nvbxx6 = (~(Pazmz6[2] & Niaxx6));
assign Eubxx6 = (Bwbxx6 & Iwbxx6);
assign Iwbxx6 = (~(Uobxx6 & Pwbxx6));
assign Pwbxx6 = (Mkbxx6 | Gnzmz6[35]);
assign Bwbxx6 = (~(Jezmz6[27] & Mt9xx6));
assign Osbxx6 = (Wwbxx6 & Dxbxx6);
assign Dxbxx6 = (Hj6xx6 | Jy6xx6);
assign Jy6xx6 = (Kxbxx6 & Rxbxx6);
assign Rxbxx6 = (~(Gnzmz6[43] & Lp9xx6));
assign Kxbxx6 = (Yxbxx6 & Fybxx6);
assign Fybxx6 = (~(Mybxx6 & Dl9xx6));
assign Mybxx6 = (Tybxx6 & Azbxx6);
assign Azbxx6 = (~(Hzbxx6 & Ozbxx6));
assign Ozbxx6 = (!Pazmz6[7]);
assign Hzbxx6 = (Vmaxx6 | Znbxx6);
assign Tybxx6 = (~(Znbxx6 & Cnaxx6));
assign Yxbxx6 = (~(Vzbxx6 & Djbxx6));
assign Wwbxx6 = (Gf6xx6 | B17xx6);
assign B17xx6 = (C0cxx6 & J0cxx6);
assign J0cxx6 = (~(Dl9xx6 & Q0cxx6));
assign Q0cxx6 = (~(X0cxx6 & E1cxx6));
assign E1cxx6 = (L1cxx6 & S1cxx6);
assign S1cxx6 = (~(Djbxx6 & Iqaxx6));
assign L1cxx6 = (~(Pazmz6[7] & Yz9xx6));
assign X0cxx6 = (Z1cxx6 & G2cxx6);
assign G2cxx6 = (~(Pazmz6[2] & Draxx6));
assign Z1cxx6 = (~(Jezmz6[35] & Dz9xx6));
assign C0cxx6 = (N2cxx6 & U2cxx6);
assign U2cxx6 = (~(Uobxx6 & B3cxx6));
assign B3cxx6 = (Mkbxx6 | Gnzmz6[27]);
assign Uobxx6 = (Mkbxx6 | Lp9xx6);
assign Mkbxx6 = (Fsaxx6 & Djbxx6);
assign Djbxx6 = (!Znbxx6);
assign Znbxx6 = (Z3axx6 & Tusnv6);
assign Z3axx6 = (Lgbxx6 & Sgbxx6);
assign Lgbxx6 = (~(Ifb7v6 & Fgzmz6[0]));
assign N2cxx6 = (~(Jezmz6[19] & Mt9xx6));
assign N2t7v6 = (I35xx6 ? Dszmz6[4] : I3cxx6);
assign G2t7v6 = (N25xx6 ? Nqzmz6[4] : I3cxx6);
assign Z1t7v6 = (On9xx6 ? I3cxx6 : Xozmz6[4]);
assign I3cxx6 = (R21nz6[2] ? G86xx6 : N86xx6);
assign G86xx6 = (~(P3cxx6 & W3cxx6));
assign W3cxx6 = (D4cxx6 & K4cxx6);
assign K4cxx6 = (Gf6xx6 | R27xx6);
assign R27xx6 = (R4cxx6 & Y4cxx6);
assign Y4cxx6 = (~(Wibxx6 & Lczmz6[2]));
assign R4cxx6 = (F5cxx6 & Cuaxx6);
assign F5cxx6 = (~(Jezmz6[4] & It7xx6));
assign D4cxx6 = (Pg6xx6 | J57xx6);
assign J57xx6 = (M5cxx6 & T5cxx6);
assign T5cxx6 = (~(A6cxx6 | H6cxx6));
assign A6cxx6 = (Jezmz6[12] & Pr9xx6);
assign M5cxx6 = (O6cxx6 & V6cxx6);
assign V6cxx6 = (~(Gnzmz6[4] & Lp9xx6));
assign O6cxx6 = (~(Hlbxx6 & Lczmz6[2]));
assign P3cxx6 = (C7cxx6 & J7cxx6);
assign J7cxx6 = (Hj6xx6 | Q57xx6);
assign Q57xx6 = (Q7cxx6 & X7cxx6);
assign X7cxx6 = (~(Dl9xx6 & E8cxx6));
assign E8cxx6 = (~(L8cxx6 & S8cxx6));
assign S8cxx6 = (Z8cxx6 | Eaaxx6);
assign L8cxx6 = (G9cxx6 & N9cxx6);
assign N9cxx6 = (~(Jezmz6[20] & Nq9xx6));
assign G9cxx6 = (~(Pazmz6[3] & J9axx6));
assign Q7cxx6 = (U9cxx6 & Bacxx6);
assign Bacxx6 = (~(Iacxx6 & Pacxx6));
assign Pacxx6 = (H6cxx6 | Gnzmz6[12]);
assign U9cxx6 = (~(Jezmz6[4] & Mt9xx6));
assign C7cxx6 = (Vj6xx6 | L67xx6);
assign L67xx6 = (Wacxx6 & Dbcxx6);
assign Dbcxx6 = (~(Dl9xx6 & Kbcxx6));
assign Kbcxx6 = (~(Rbcxx6 & Ybcxx6));
assign Ybcxx6 = (Fccxx6 & Mccxx6);
assign Mccxx6 = (~(Jezmz6[28] & Au9xx6));
assign Fccxx6 = (~(Pazmz6[3] & Feaxx6));
assign Rbcxx6 = (Tccxx6 & Adcxx6);
assign Adcxx6 = (~(Pazmz6[8] & Vu9xx6));
assign Tccxx6 = (Z8cxx6 | Kdaxx6);
assign Wacxx6 = (Hdcxx6 & Odcxx6);
assign Odcxx6 = (~(Iacxx6 & Vdcxx6));
assign Vdcxx6 = (H6cxx6 | Gnzmz6[20]);
assign Hdcxx6 = (~(Jezmz6[12] & Mt9xx6));
assign N86xx6 = (~(Cecxx6 & Jecxx6));
assign Jecxx6 = (Qecxx6 & Xecxx6);
assign Xecxx6 = (Vj6xx6 | Y27xx6);
assign Y27xx6 = (Efcxx6 & Z8cxx6);
assign Efcxx6 = (~(Emc7v6 & Lp9xx6));
assign Qecxx6 = (Pg6xx6 | T37xx6);
assign T37xx6 = (Lfcxx6 & Sfcxx6);
assign Sfcxx6 = (~(Dl9xx6 & Zfcxx6));
assign Zfcxx6 = (~(Ggcxx6 & Ngcxx6));
assign Ngcxx6 = (~(Pazmz6[8] & Zw9xx6));
assign Zw9xx6 = (!Ugcxx6);
assign Ggcxx6 = (Bhcxx6 & Ihcxx6);
assign Ihcxx6 = (~(Pazmz6[3] & Niaxx6));
assign Bhcxx6 = (Z8cxx6 | Giaxx6);
assign Lfcxx6 = (Phcxx6 & Whcxx6);
assign Whcxx6 = (~(Iacxx6 & Dicxx6));
assign Dicxx6 = (H6cxx6 | Gnzmz6[36]);
assign Phcxx6 = (~(Jezmz6[28] & Mt9xx6));
assign Cecxx6 = (Kicxx6 & Ricxx6);
assign Ricxx6 = (Hj6xx6 | A47xx6);
assign A47xx6 = (Yicxx6 & Fjcxx6);
assign Fjcxx6 = (Mjcxx6 & Kkaxx6);
assign Mjcxx6 = (~(Gnzmz6[44] & Lp9xx6));
assign Yicxx6 = (Tjcxx6 & Akcxx6);
assign Akcxx6 = (~(Lczmz6[2] & Hkcxx6));
assign Tjcxx6 = (~(Okcxx6 & Pazmz6[8]));
assign Okcxx6 = (T0axx6 & Dl9xx6);
assign Kicxx6 = (Gf6xx6 | S67xx6);
assign S67xx6 = (Vkcxx6 & Clcxx6);
assign Clcxx6 = (~(Dl9xx6 & Jlcxx6));
assign Jlcxx6 = (~(Qlcxx6 & Xlcxx6));
assign Xlcxx6 = (Emcxx6 & Lmcxx6);
assign Emcxx6 = (~(Pazmz6[8] & Yz9xx6));
assign Qlcxx6 = (Smcxx6 & Zmcxx6);
assign Zmcxx6 = (~(Pazmz6[3] & Draxx6));
assign Smcxx6 = (~(Lczmz6[2] & Iqaxx6));
assign Vkcxx6 = (Gncxx6 & Nncxx6);
assign Nncxx6 = (~(Iacxx6 & Uncxx6));
assign Uncxx6 = (H6cxx6 | Gnzmz6[28]);
assign Iacxx6 = (H6cxx6 | Lp9xx6);
assign H6cxx6 = (Fsaxx6 & Lczmz6[2]);
assign Gncxx6 = (~(Jezmz6[20] & Mt9xx6));
assign S1t7v6 = (I35xx6 ? Dszmz6[5] : Bocxx6);
assign L1t7v6 = (N25xx6 ? Nqzmz6[5] : Bocxx6);
assign E1t7v6 = (On9xx6 ? Bocxx6 : Xozmz6[5]);
assign Bocxx6 = (R21nz6[2] ? B96xx6 : I96xx6);
assign B96xx6 = (~(Iocxx6 & Pocxx6));
assign Pocxx6 = (Wocxx6 & Dpcxx6);
assign Dpcxx6 = (Gf6xx6 | I87xx6);
assign I87xx6 = (Kpcxx6 & Rpcxx6);
assign Rpcxx6 = (~(Wibxx6 & Lczmz6[3]));
assign Wibxx6 = (~(Ypcxx6 | Ro87v6));
assign Kpcxx6 = (Fqcxx6 & Cuaxx6);
assign Fqcxx6 = (~(Jezmz6[5] & It7xx6));
assign It7xx6 = (Pr9xx6 | Mqcxx6);
assign Mqcxx6 = (Dl9xx6 & Ro87v6);
assign Wocxx6 = (Pg6xx6 | Ab7xx6);
assign Ab7xx6 = (Tqcxx6 & Arcxx6);
assign Arcxx6 = (Hrcxx6 & Orcxx6);
assign Orcxx6 = (~(Gnzmz6[5] & Lp9xx6));
assign Hrcxx6 = (Vrcxx6 & Cscxx6);
assign Vrcxx6 = (~(Jezmz6[13] & Pr9xx6));
assign Pr9xx6 = (Dl9xx6 & Jscxx6);
assign Jscxx6 = (!F7axx6);
assign Tqcxx6 = (Qscxx6 & Xscxx6);
assign Xscxx6 = (~(Jezmz6[32] & Mt9xx6));
assign Qscxx6 = (~(Hlbxx6 & Lczmz6[3]));
assign Iocxx6 = (Etcxx6 & Ltcxx6);
assign Ltcxx6 = (Hj6xx6 | Hb7xx6);
assign Hb7xx6 = (Stcxx6 & Ztcxx6);
assign Ztcxx6 = (Gucxx6 & Cscxx6);
assign Gucxx6 = (~(Jezmz6[5] & Mt9xx6));
assign Stcxx6 = (Nucxx6 & Uucxx6);
assign Uucxx6 = (~(Dl9xx6 & Bvcxx6));
assign Bvcxx6 = (~(Ivcxx6 & Pvcxx6));
assign Pvcxx6 = (Wvcxx6 | Eaaxx6);
assign Ivcxx6 = (Dwcxx6 & Kwcxx6);
assign Kwcxx6 = (~(Jezmz6[21] & Nq9xx6));
assign Dwcxx6 = (~(W1a7v6 & J9axx6));
assign Nucxx6 = (~(Gnzmz6[13] & Lp9xx6));
assign Etcxx6 = (Vj6xx6 | Cc7xx6);
assign Cc7xx6 = (Rwcxx6 & Ywcxx6);
assign Ywcxx6 = (Fxcxx6 & Cscxx6);
assign Cscxx6 = (~(Fsaxx6 & Lczmz6[3]));
assign Fxcxx6 = (~(Jezmz6[13] & Mt9xx6));
assign Rwcxx6 = (Mxcxx6 & Txcxx6);
assign Txcxx6 = (~(Dl9xx6 & Aycxx6));
assign Aycxx6 = (~(Hycxx6 & Oycxx6));
assign Oycxx6 = (Wvcxx6 | Kdaxx6);
assign Hycxx6 = (Vycxx6 & Czcxx6);
assign Czcxx6 = (~(Jezmz6[29] & Au9xx6));
assign Vycxx6 = (~(W1a7v6 & Feaxx6));
assign Mxcxx6 = (~(Gnzmz6[21] & Lp9xx6));
assign I96xx6 = (~(Jzcxx6 & Qzcxx6));
assign Qzcxx6 = (Xzcxx6 & E0dxx6);
assign E0dxx6 = (Vj6xx6 | P87xx6);
assign P87xx6 = (L0dxx6 & Wvcxx6);
assign L0dxx6 = (~(Ync7v6 & Lp9xx6));
assign Xzcxx6 = (Pg6xx6 | K97xx6);
assign K97xx6 = (S0dxx6 & Z0dxx6);
assign Z0dxx6 = (G1dxx6 & N1dxx6);
assign N1dxx6 = (~(Jezmz6[29] & Mt9xx6));
assign G1dxx6 = (~(U1dxx6 & W1a7v6));
assign U1dxx6 = (Dl9xx6 & Niaxx6);
assign S0dxx6 = (B2dxx6 & I2dxx6);
assign I2dxx6 = (~(Lczmz6[3] & P2dxx6));
assign B2dxx6 = (~(Gnzmz6[37] & Lp9xx6));
assign Jzcxx6 = (W2dxx6 & D3dxx6);
assign D3dxx6 = (Hj6xx6 | R97xx6);
assign R97xx6 = (K3dxx6 & R3dxx6);
assign R3dxx6 = (~(Gnzmz6[45] & Lp9xx6));
assign K3dxx6 = (Y3dxx6 & Kkaxx6);
assign Y3dxx6 = (~(Lczmz6[3] & Hkcxx6));
assign W2dxx6 = (Gf6xx6 | Jc7xx6);
assign Jc7xx6 = (F4dxx6 & M4dxx6);
assign M4dxx6 = (T4dxx6 & A5dxx6);
assign A5dxx6 = (~(Jezmz6[21] & Mt9xx6));
assign T4dxx6 = (~(H5dxx6 & W1a7v6));
assign H5dxx6 = (Dl9xx6 & Draxx6);
assign F4dxx6 = (O5dxx6 & V5dxx6);
assign V5dxx6 = (~(Lczmz6[3] & C6dxx6));
assign C6dxx6 = (~(J6dxx6 & Cuaxx6));
assign J6dxx6 = (~(Dl9xx6 & Iqaxx6));
assign O5dxx6 = (~(Gnzmz6[29] & Lp9xx6));
assign X0t7v6 = (I35xx6 ? Dszmz6[6] : Q6dxx6);
assign Q0t7v6 = (N25xx6 ? Nqzmz6[6] : Q6dxx6);
assign J0t7v6 = (On9xx6 ? Q6dxx6 : Xozmz6[6]);
assign Q6dxx6 = (R21nz6[2] ? W96xx6 : Da6xx6);
assign W96xx6 = (~(X6dxx6 & E7dxx6));
assign E7dxx6 = (L7dxx6 & S7dxx6);
assign S7dxx6 = (Ne7xx6 | Gf6xx6);
assign Ne7xx6 = (~(Z7dxx6 & G8dxx6));
assign G8dxx6 = (~(X2axx6 & N8dxx6));
assign N8dxx6 = (~(Dl9xx6 & U8dxx6));
assign U8dxx6 = (B9dxx6 | Jezmz6[6]);
assign B9dxx6 = (~(I9dxx6 | Ro87v6));
assign Z7dxx6 = (P9dxx6 | N4axx6);
assign N4axx6 = (~(W9dxx6 & F7axx6));
assign W9dxx6 = (X2axx6 & Zvaxx6);
assign L7dxx6 = (Pg6xx6 | Yg7xx6);
assign Yg7xx6 = (Dadxx6 & Kadxx6);
assign Kadxx6 = (~(Radxx6 & Dl9xx6));
assign Radxx6 = (Yadxx6 & Fbdxx6);
assign Fbdxx6 = (Mbdxx6 | Jezmz6[14]);
assign Mbdxx6 = (~(I9dxx6 | Y6axx6));
assign Yadxx6 = (~(I9dxx6 & F7axx6));
assign F7axx6 = (~(Tbdxx6 | J9axx6));
assign Tbdxx6 = (Nq9xx6 | Y6axx6);
assign Dadxx6 = (Acdxx6 & Hcdxx6);
assign Hcdxx6 = (~(Jezmz6[33] & Mt9xx6));
assign Acdxx6 = (~(Ocdxx6 & Vcdxx6));
assign Vcdxx6 = (Cddxx6 | Gnzmz6[6]);
assign X6dxx6 = (Jddxx6 & Qddxx6);
assign Qddxx6 = (Hj6xx6 | Fh7xx6);
assign Fh7xx6 = (Xddxx6 & Eedxx6);
assign Eedxx6 = (~(Dl9xx6 & Ledxx6));
assign Ledxx6 = (~(Sedxx6 & Zedxx6));
assign Zedxx6 = (I9dxx6 | Eaaxx6);
assign Sedxx6 = (~(Jezmz6[22] & Nq9xx6));
assign Nq9xx6 = (Gfdxx6 | Au9xx6);
assign Gfdxx6 = (Feaxx6 | Nfdxx6);
assign Xddxx6 = (Ufdxx6 & Bgdxx6);
assign Bgdxx6 = (~(Jezmz6[6] & Mt9xx6));
assign Ufdxx6 = (~(Ocdxx6 & Igdxx6));
assign Igdxx6 = (Cddxx6 | Gnzmz6[14]);
assign Jddxx6 = (Vj6xx6 | Ai7xx6);
assign Ai7xx6 = (Pgdxx6 & Wgdxx6);
assign Wgdxx6 = (~(Dl9xx6 & Dhdxx6));
assign Dhdxx6 = (~(Khdxx6 & Rhdxx6));
assign Rhdxx6 = (I9dxx6 | Kdaxx6);
assign Khdxx6 = (~(Jezmz6[30] & Au9xx6));
assign Au9xx6 = (Yhdxx6 | Draxx6);
assign Yhdxx6 = (~(Fidxx6 & Lmcxx6));
assign Pgdxx6 = (Midxx6 & Tidxx6);
assign Tidxx6 = (~(Jezmz6[14] & Mt9xx6));
assign Midxx6 = (~(Ocdxx6 & Ajdxx6));
assign Ajdxx6 = (Cddxx6 | Gnzmz6[22]);
assign Da6xx6 = (~(Hjdxx6 & Ojdxx6));
assign Ojdxx6 = (Vjdxx6 & Ckdxx6);
assign Ckdxx6 = (~(Zd7xx6 & Jkdxx6));
assign Zd7xx6 = (P9dxx6 & Ym8xx6);
assign Vjdxx6 = (Pg6xx6 | If7xx6);
assign If7xx6 = (Qkdxx6 & Xkdxx6);
assign Xkdxx6 = (~(Jezmz6[30] & Mt9xx6));
assign Qkdxx6 = (Eldxx6 & Lldxx6);
assign Lldxx6 = (~(P9dxx6 & P2dxx6));
assign P2dxx6 = (~(Sldxx6 & Cuaxx6));
assign Sldxx6 = (Ypcxx6 | Giaxx6);
assign Eldxx6 = (~(Gnzmz6[38] & Lp9xx6));
assign Hjdxx6 = (Zldxx6 & Gmdxx6);
assign Gmdxx6 = (Hj6xx6 | Pf7xx6);
assign Pf7xx6 = (Nmdxx6 & Umdxx6);
assign Umdxx6 = (~(Gnzmz6[46] & Lp9xx6));
assign Nmdxx6 = (Bndxx6 & Kkaxx6);
assign Bndxx6 = (~(Indxx6 & P9dxx6));
assign Indxx6 = (Hkcxx6 & Ym8xx6);
assign Hkcxx6 = (~(Vmaxx6 & Flaxx6));
assign Zldxx6 = (Gf6xx6 | Hi7xx6);
assign Hi7xx6 = (Pndxx6 & Wndxx6);
assign Wndxx6 = (~(Dl9xx6 & Dodxx6));
assign Dodxx6 = (~(Kodxx6 & Rodxx6));
assign Rodxx6 = (~(P9dxx6 & Iqaxx6));
assign P9dxx6 = (!I9dxx6);
assign Kodxx6 = (~(Dz9xx6 & Yodxx6));
assign Pndxx6 = (Fpdxx6 & Mpdxx6);
assign Mpdxx6 = (~(Jezmz6[22] & Mt9xx6));
assign Fpdxx6 = (~(Ocdxx6 & Tpdxx6));
assign Tpdxx6 = (Cddxx6 | Gnzmz6[30]);
assign Ocdxx6 = (Cddxx6 | Lp9xx6);
assign Cddxx6 = (~(Cuaxx6 | I9dxx6));
assign I9dxx6 = (Ifb7v6 ? Fgzmz6[0] : Aqdxx6);
assign Aqdxx6 = (~(Pdtnv6 & Sgbxx6));
assign C0t7v6 = (I35xx6 ? Dszmz6[7] : Hqdxx6);
assign I35xx6 = (~(Ef5xx6 & Ce5xx6));
assign Ef5xx6 = (Oqdxx6 & Vqdxx6);
assign Oqdxx6 = (!B41nz6[1]);
assign Vzs7v6 = (N25xx6 ? Nqzmz6[7] : Hqdxx6);
assign N25xx6 = (~(Ce5xx6 & Fc5xx6));
assign Fc5xx6 = (~(Vqdxx6 | B41nz6[1]));
assign Ozs7v6 = (On9xx6 ? Hqdxx6 : Xozmz6[7]);
assign On9xx6 = (Crdxx6 & Ce5xx6);
assign Ce5xx6 = (!B35xx6);
assign B35xx6 = (~(Jrdxx6 & Fftnv6));
assign Fftnv6 = (~(Qrdxx6 & Zkrnv6));
assign Zkrnv6 = (Xrdxx6 ? K6d7v6 : Cuc7v6);
assign Qrdxx6 = (Esdxx6 & Lsdxx6);
assign Lsdxx6 = (~(Ssdxx6 & Zsdxx6));
assign Zsdxx6 = (Bgt8v6 ? Ntdxx6 : Gtdxx6);
assign Ntdxx6 = (Qqrnv6 | Skcov6);
assign Qqrnv6 = (!Zrrnv6);
assign Gtdxx6 = (~(Skcov6 & Utdxx6));
assign Utdxx6 = (Budxx6 | Zrrnv6);
assign Ssdxx6 = (Iudxx6 & Pudxx6);
assign Pudxx6 = (~(Wudxx6 & Budxx6));
assign Budxx6 = (~(Durnv6 & Dvdxx6));
assign Dvdxx6 = (~(Skcov6 & Errnv6));
assign Durnv6 = (!Kvdxx6);
assign Kvdxx6 = (Xrdxx6 ? Cad7v6 : Uxc7v6);
assign Wudxx6 = (~(Rvdxx6 & Yvdxx6));
assign Yvdxx6 = (~(Fwdxx6 & Mwdxx6));
assign Mwdxx6 = (~(Gsrnv6 & Twdxx6));
assign Gsrnv6 = (!Errnv6);
assign Errnv6 = (Xrdxx6 ? Ibd7v6 : Azc7v6);
assign Fwdxx6 = (Axdxx6 & Let8v6);
assign Axdxx6 = (Zrrnv6 | Bgt8v6);
assign Rvdxx6 = (~(Skcov6 & Zrrnv6));
assign Zrrnv6 = (Xrdxx6 ? W8d7v6 : Owc7v6);
assign Iudxx6 = (~(Fvrnv6 & Hxdxx6));
assign Esdxx6 = (~(Oxdxx6 & Imrnv6));
assign Imrnv6 = (!Fvrnv6);
assign Fvrnv6 = (Xrdxx6 ? Q7d7v6 : Ivc7v6);
assign Xrdxx6 = (~(Vxdxx6 & Cydxx6));
assign Cydxx6 = (~(E11nz6[4] & Owrnv6));
assign Vxdxx6 = (Jydxx6 & Nlcov6);
assign Jydxx6 = (~(Qydxx6 & Xydxx6));
assign Xydxx6 = (~(Rr0nz6[1] & Pp4xx6));
assign Pp4xx6 = (!E11nz6[4]);
assign Qydxx6 = (Ezdxx6 & Lzdxx6);
assign Lzdxx6 = (~(Szdxx6 & Zzdxx6));
assign Zzdxx6 = (~(E11nz6[3] & Cxrnv6));
assign Szdxx6 = (G0exx6 & N0exx6);
assign N0exx6 = (~(U0exx6 & B1exx6));
assign B1exx6 = (E11nz6[1] | I1exx6);
assign I1exx6 = (P1exx6 & E11nz6[0]);
assign P1exx6 = (Lyrnv6 & Qqcov6);
assign U0exx6 = (~(W1exx6 & D2exx6));
assign D2exx6 = (~(E11nz6[2] & Qqcov6));
assign W1exx6 = (K2exx6 & Jxrnv6);
assign K2exx6 = (~(R2exx6 & E11nz6[0]));
assign R2exx6 = (Y2exx6 & Lyrnv6);
assign Y2exx6 = (~(Hw0nz6[2] & Mocov6));
assign Mocov6 = (!E11nz6[2]);
assign G0exx6 = (~(E11nz6[2] & Ercov6));
assign Ezdxx6 = (~(Rr0nz6[0] & No4xx6));
assign No4xx6 = (!E11nz6[3]);
assign Oxdxx6 = (!Hxdxx6);
assign Hxdxx6 = (~(Qjcov6 & Skcov6));
assign Skcov6 = (Twdxx6 & Zi9xx6);
assign Twdxx6 = (!Wsc7v6);
assign Qjcov6 = (~(Bgt8v6 | Rht8v6));
assign Jrdxx6 = (~(F3exx6 & M3exx6));
assign M3exx6 = (~(T51nz6[2] & T3exx6));
assign F3exx6 = (~(A4exx6 | Rht8v6));
assign Rht8v6 = (H4exx6 | O4exx6);
assign H4exx6 = (V4exx6 & C5exx6);
assign A4exx6 = (~(J5exx6 | Q5exx6));
assign Q5exx6 = (!Bgt8v6);
assign Crdxx6 = (B41nz6[1] & Vqdxx6);
assign Vqdxx6 = (!B41nz6[0]);
assign Hqdxx6 = (R21nz6[2] ? Cd6xx6 : Jd6xx6);
assign Cd6xx6 = (~(X5exx6 & E6exx6));
assign E6exx6 = (L6exx6 & S6exx6);
assign S6exx6 = (~(Dm8xx6 & Zb9xx6));
assign Dm8xx6 = (Dl9xx6 & Kl9xx6);
assign Kl9xx6 = (Zvaxx6 | Jezmz6[7]);
assign L6exx6 = (Pg6xx6 | Cq7xx6);
assign Cq7xx6 = (Z6exx6 & G7exx6);
assign G7exx6 = (~(Hlbxx6 | Fsaxx6));
assign Hlbxx6 = (~(Ypcxx6 | Y6axx6));
assign Z6exx6 = (N7exx6 & U7exx6);
assign U7exx6 = (~(Dl9xx6 & Jezmz6[15]));
assign N7exx6 = (~(B987v6 & Lp9xx6));
assign X5exx6 = (B8exx6 & I8exx6);
assign I8exx6 = (Hj6xx6 | Jq7xx6);
assign Jq7xx6 = (P8exx6 & W8exx6);
assign W8exx6 = (~(Dl9xx6 & D9exx6));
assign D9exx6 = (~(K9exx6 & Eaaxx6));
assign K9exx6 = (~(R9exx6 | Jezmz6[23]));
assign R9exx6 = (Y9exx6 & J9axx6);
assign J9axx6 = (Vu9xx6 | Faexx6);
assign Faexx6 = (Maexx6 & Taexx6);
assign P8exx6 = (Abexx6 & Hbexx6);
assign Hbexx6 = (~(Mt9xx6 & Jezmz6[7]));
assign Abexx6 = (~(Obexx6 & Vbexx6));
assign Vbexx6 = (Fsaxx6 | Gnzmz6[15]);
assign B8exx6 = (Vj6xx6 | Er7xx6);
assign Er7xx6 = (Ccexx6 & Jcexx6);
assign Jcexx6 = (~(Dl9xx6 & Qcexx6));
assign Qcexx6 = (~(Xcexx6 & Kdaxx6));
assign Xcexx6 = (Edexx6 & Ldexx6);
assign Ldexx6 = (!Jezmz6[31]);
assign Edexx6 = (~(Y9exx6 & Feaxx6));
assign Feaxx6 = (Yz9xx6 | Sdexx6);
assign Ccexx6 = (Zdexx6 & Geexx6);
assign Geexx6 = (~(Mt9xx6 & Jezmz6[15]));
assign Zdexx6 = (~(Obexx6 & Neexx6));
assign Neexx6 = (~(Cuaxx6 & Ueexx6));
assign Vj6xx6 = (!Jkdxx6);
assign Jd6xx6 = (~(Bfexx6 & Ifexx6));
assign Ifexx6 = (Pfexx6 & Wfexx6);
assign Wfexx6 = (Pg6xx6 | To7xx6);
assign To7xx6 = (Dgexx6 & Kgexx6);
assign Kgexx6 = (~(Dl9xx6 & Rgexx6));
assign Rgexx6 = (~(Giaxx6 & Ygexx6));
assign Ygexx6 = (~(Y9exx6 & Niaxx6));
assign Niaxx6 = (~(Cnaxx6 & Fhexx6));
assign Fhexx6 = (~(Maexx6 & Dz9xx6));
assign Cnaxx6 = (!T0axx6);
assign T0axx6 = (Mhexx6 & Dz9xx6);
assign Dgexx6 = (Thexx6 & Aiexx6);
assign Aiexx6 = (~(Mt9xx6 & Jezmz6[31]));
assign Thexx6 = (~(Obexx6 & Hiexx6));
assign Hiexx6 = (~(Cuaxx6 & Oiexx6));
assign Pg6xx6 = (!Df8xx6);
assign Df8xx6 = (~(Du7xx6 | R21nz6[0]));
assign Pfexx6 = (Hj6xx6 | Rn7xx6);
assign Rn7xx6 = (Viexx6 & Cjexx6);
assign Cjexx6 = (Ypcxx6 | Vmaxx6);
assign Vmaxx6 = (Jjexx6 & Giaxx6);
assign Giaxx6 = (Qjexx6 & Xjexx6);
assign Xjexx6 = (Ekexx6 & Lkexx6);
assign Lkexx6 = (!Yz9xx6);
assign Yz9xx6 = (Mhexx6 & Skexx6);
assign Qjexx6 = (Zkexx6 & Yodxx6);
assign Jjexx6 = (Ugcxx6 & Glexx6);
assign Viexx6 = (~(Vzbxx6 | O4exx6));
assign O4exx6 = (Ka87v6 & Lp9xx6);
assign Vzbxx6 = (~(Flaxx6 | Nlexx6));
assign Nlexx6 = (Ztb7v6 & Cuaxx6);
assign Hj6xx6 = (!Ge7xx6);
assign Ge7xx6 = (~(Ulexx6 | R21nz6[1]));
assign Bfexx6 = (Bmexx6 & Imexx6);
assign Imexx6 = (Gf6xx6 | Lr7xx6);
assign Lr7xx6 = (Pmexx6 & Wmexx6);
assign Wmexx6 = (~(Dl9xx6 & Dnexx6));
assign Dnexx6 = (~(Zkexx6 & Knexx6));
assign Knexx6 = (~(Y9exx6 & Draxx6));
assign Draxx6 = (~(Ugcxx6 & Ekexx6));
assign Ekexx6 = (~(Rnexx6 & Maexx6));
assign Ugcxx6 = (~(Rnexx6 & Mhexx6));
assign Rnexx6 = (Ynexx6 & Lmcxx6);
assign Zkexx6 = (!Iqaxx6);
assign Iqaxx6 = (~(Foexx6 & Moexx6));
assign Moexx6 = (~(Sdexx6 | Vu9xx6));
assign Vu9xx6 = (Mhexx6 & Taexx6);
assign Sdexx6 = (~(Glexx6 | Toexx6));
assign Foexx6 = (Kdaxx6 & Apexx6);
assign Apexx6 = (Fidxx6 | Dz9xx6);
assign Fidxx6 = (~(Ynexx6 & Hpexx6));
assign Kdaxx6 = (Opexx6 & Eaaxx6);
assign Eaaxx6 = (Y6axx6 & Vpexx6);
assign Vpexx6 = (~(Hpexx6 & Taexx6));
assign Opexx6 = (Cqexx6 & Jqexx6);
assign Cqexx6 = (~(Maexx6 & Taexx6));
assign Pmexx6 = (Qqexx6 & Xqexx6);
assign Xqexx6 = (~(Mt9xx6 & Jezmz6[23]));
assign Qqexx6 = (~(Obexx6 & Erexx6));
assign Erexx6 = (~(Cuaxx6 & Lrexx6));
assign Obexx6 = (!X2axx6);
assign X2axx6 = (Cuaxx6 & I0snv6);
assign Gf6xx6 = (!Zb9xx6);
assign Zb9xx6 = (~(Du7xx6 | Ulexx6));
assign Ulexx6 = (!R21nz6[0]);
assign Du7xx6 = (!R21nz6[1]);
assign Bmexx6 = (~(Jkdxx6 & Ym8xx6));
assign Ym8xx6 = (~(Flaxx6 & Ypcxx6));
assign Ypcxx6 = (!Dl9xx6);
assign Flaxx6 = (Zp9xx6 & Cuaxx6);
assign Jkdxx6 = (~(R21nz6[0] | R21nz6[1]));
assign Hzs7v6 = (~(Srexx6 & Zrexx6));
assign Zrexx6 = (~(Gsexx6 & Nsexx6));
assign Nsexx6 = (~(Usexx6 & Btexx6));
assign Btexx6 = (Itexx6 & Ptexx6);
assign Ptexx6 = (Wtexx6 & Duexx6);
assign Duexx6 = (Kuexx6 & Ruexx6);
assign Ruexx6 = (~(Yuexx6 & Bq0nz6[0]));
assign Kuexx6 = (Fvexx6 & Mvexx6);
assign Mvexx6 = (~(Tvexx6 & Fl0nz6[0]));
assign Fvexx6 = (~(Awexx6 & Jg0nz6[0]));
assign Wtexx6 = (Hwexx6 & Owexx6);
assign Owexx6 = (~(Vwexx6 & Nb0nz6[0]));
assign Hwexx6 = (Cxexx6 & Jxexx6);
assign Jxexx6 = (~(Qxexx6 & R60nz6[0]));
assign Cxexx6 = (~(Xxexx6 & V10nz6[0]));
assign Itexx6 = (Eyexx6 & Lyexx6);
assign Lyexx6 = (Syexx6 & Zyexx6);
assign Zyexx6 = (~(Gzexx6 & Zwzmz6[0]));
assign Syexx6 = (Nzexx6 & Uzexx6);
assign Uzexx6 = (~(B0fxx6 & Dszmz6[0]));
assign Nzexx6 = (~(I0fxx6 & Lo0nz6[0]));
assign Eyexx6 = (P0fxx6 & W0fxx6);
assign W0fxx6 = (~(D1fxx6 & Pj0nz6[0]));
assign P0fxx6 = (K1fxx6 & R1fxx6);
assign R1fxx6 = (~(Y1fxx6 & Te0nz6[0]));
assign K1fxx6 = (~(F2fxx6 & X90nz6[0]));
assign Usexx6 = (M2fxx6 & T2fxx6);
assign T2fxx6 = (A3fxx6 & H3fxx6);
assign H3fxx6 = (O3fxx6 & V3fxx6);
assign V3fxx6 = (~(C4fxx6 & B50nz6[0]));
assign O3fxx6 = (J4fxx6 & Q4fxx6);
assign Q4fxx6 = (~(X4fxx6 & F00nz6[0]));
assign J4fxx6 = (~(E5fxx6 & Jvzmz6[0]));
assign A3fxx6 = (L5fxx6 & S5fxx6);
assign S5fxx6 = (~(Z5fxx6 & Nqzmz6[0]));
assign L5fxx6 = (G6fxx6 & N6fxx6);
assign N6fxx6 = (~(U6fxx6 & Vm0nz6[0]));
assign G6fxx6 = (~(B7fxx6 & Zh0nz6[0]));
assign M2fxx6 = (I7fxx6 & P7fxx6);
assign P7fxx6 = (W7fxx6 & D8fxx6);
assign D8fxx6 = (~(K8fxx6 & Dd0nz6[0]));
assign W7fxx6 = (R8fxx6 & Y8fxx6);
assign Y8fxx6 = (~(F9fxx6 & H80nz6[0]));
assign R8fxx6 = (~(M9fxx6 & L30nz6[0]));
assign I7fxx6 = (T9fxx6 & Aafxx6);
assign Aafxx6 = (~(Xozmz6[0] & Hafxx6));
assign T9fxx6 = (Oafxx6 & Vafxx6);
assign Vafxx6 = (~(Cbfxx6 & Ttzmz6[0]));
assign Oafxx6 = (~(Jbfxx6 & Pyzmz6[0]));
assign Srexx6 = (~(Ak67z6 & Lr5ov6));
assign Azs7v6 = (Cmtiw6 ? D7hdt6 : L0g7z6[32]);
assign Tys7v6 = (~(Qbfxx6 & Xbfxx6));
assign Xbfxx6 = (~(Yj2ov6 & Yxf7z6[0]));
assign Qbfxx6 = (Ecfxx6 & Lcfxx6);
assign Lcfxx6 = (Scfxx6 | Wi2ov6);
assign Scfxx6 = (T1lhw6 ? Ubpdt6 : Epmdt6);
assign T1lhw6 = (Pcg7z6[31] ^ Elgdt6);
assign Pcg7z6[31] = (Qamnv6 ? Wiudt6 : Ixrdt6);
assign Qamnv6 = (~(D4wnv6 ^ Zfg7z6[32]));
assign D4wnv6 = (!Elgdt6);
assign Ecfxx6 = (~(Bnmdt6 & Rj2ov6));
assign Mys7v6 = (~(Zcfxx6 & Gdfxx6));
assign Gdfxx6 = (~(Y3bov6 & Yxf7z6[0]));
assign Zcfxx6 = (Ndfxx6 & Udfxx6);
assign Udfxx6 = (~(Rj2ov6 & Pemdt6));
assign Ndfxx6 = (~(Yj2ov6 & Yxf7z6[4]));
assign Fys7v6 = (~(Befxx6 & Iefxx6));
assign Iefxx6 = (~(Y3bov6 & Yxf7z6[4]));
assign Befxx6 = (Pefxx6 & Wefxx6);
assign Wefxx6 = (~(Rj2ov6 & D6mdt6));
assign Pefxx6 = (~(Yj2ov6 & Yxf7z6[8]));
assign Yxs7v6 = (~(Dffxx6 & Kffxx6));
assign Kffxx6 = (~(Y3bov6 & Yxf7z6[8]));
assign Dffxx6 = (Rffxx6 & Yffxx6);
assign Yffxx6 = (~(Rj2ov6 & Rxldt6));
assign Rffxx6 = (~(Yj2ov6 & Yxf7z6[12]));
assign Rxs7v6 = (~(Fgfxx6 & Mgfxx6));
assign Mgfxx6 = (~(Y3bov6 & Yxf7z6[12]));
assign Fgfxx6 = (Tgfxx6 & Ahfxx6);
assign Ahfxx6 = (~(Rj2ov6 & Fpldt6));
assign Tgfxx6 = (~(Yj2ov6 & Yxf7z6[16]));
assign Kxs7v6 = (~(Hhfxx6 & Ohfxx6));
assign Ohfxx6 = (~(Y3bov6 & Yxf7z6[16]));
assign Hhfxx6 = (Vhfxx6 & Cifxx6);
assign Cifxx6 = (~(Rj2ov6 & Tgldt6));
assign Vhfxx6 = (~(Yj2ov6 & Yxf7z6[20]));
assign Dxs7v6 = (~(Jifxx6 & Qifxx6));
assign Qifxx6 = (~(Y3bov6 & Yxf7z6[20]));
assign Jifxx6 = (Xifxx6 & Ejfxx6);
assign Ejfxx6 = (~(Rj2ov6 & H8ldt6));
assign Xifxx6 = (~(Yj2ov6 & Yxf7z6[24]));
assign Wws7v6 = (~(Ljfxx6 & Sjfxx6));
assign Sjfxx6 = (~(Y3bov6 & Yxf7z6[24]));
assign Ljfxx6 = (Zjfxx6 & Gkfxx6);
assign Gkfxx6 = (~(Rj2ov6 & Vzkdt6));
assign Rj2ov6 = (Nkfxx6 & Ukfxx6);
assign Ukfxx6 = (~(Blfxx6 | Yj2ov6));
assign Blfxx6 = (Ijnnv6 | Rabov6);
assign Ijnnv6 = (!Kxtiw6);
assign Nkfxx6 = (Dfkov6 & Ilfxx6);
assign Zjfxx6 = (~(Yj2ov6 & Yxf7z6[28]));
assign Pws7v6 = (~(Plfxx6 & Wlfxx6));
assign Wlfxx6 = (~(Yj2ov6 & Yxf7z6[32]));
assign Yj2ov6 = (Yzm7x6 & Dmfxx6);
assign Dmfxx6 = (Kmfxx6 & Yqtiw6);
assign Yqtiw6 = (~(Rabov6 & Rmfxx6));
assign Rmfxx6 = (~(Ymfxx6 & Fnfxx6));
assign Ymfxx6 = (~(Go37x6 & Mnfxx6));
assign Rabov6 = (!Z6jhw6);
assign Kmfxx6 = (Wi2ov6 & Kxtiw6);
assign Yzm7x6 = (~(L7bov6 | E7bov6));
assign E7bov6 = (~(Tnfxx6 & Ts27x6));
assign Tnfxx6 = (Aofxx6 & Qariw6);
assign Qariw6 = (~(Dqtiw6 & Ehgdt6));
assign L7bov6 = (~(Ilfxx6 & A127x6));
assign Plfxx6 = (~(Y3bov6 & Yxf7z6[28]));
assign Iws7v6 = (Diaov6 ? Hofxx6 : Pmc7z6[2]);
assign Diaov6 = (!Riaov6);
assign Riaov6 = (Oofxx6 & Phaov6);
assign Phaov6 = (Pooov6 & Vofxx6);
assign Vofxx6 = (Cpfxx6 & Jpfxx6);
assign Jpfxx6 = (D61ov6 | Qpfxx6);
assign Qpfxx6 = (Xpfxx6 & Eqfxx6);
assign Xpfxx6 = (Hkoov6 & Lqfxx6);
assign D61ov6 = (Sqfxx6 & Qv0ov6);
assign Sqfxx6 = (!G8xnv6);
assign G8xnv6 = (~(Zqfxx6 & Grfxx6));
assign Zqfxx6 = (~(Jamnv6 & A9mnv6));
assign Cpfxx6 = (Jsoov6 & Pj1ov6);
assign Pooov6 = (Q0wnv6 & O4piw6);
assign Oofxx6 = (Femhw6 & Ij1ov6);
assign Ij1ov6 = (!Cg1ov6);
assign Femhw6 = (~(Nrfxx6 & N3onv6));
assign Nrfxx6 = (Urfxx6 & Fetov6);
assign Urfxx6 = (~(Bsfxx6 & Isfxx6));
assign Bsfxx6 = (Tao7v6 & J9tov6);
assign Bws7v6 = (~(Psfxx6 & Wsfxx6));
assign Wsfxx6 = (~(Dtfxx6 & Ktfxx6));
assign Dtfxx6 = (Osd7z6[2] & Vs9ov6);
assign Psfxx6 = (~(Rtfxx6 & Rem7x6));
assign Rtfxx6 = (Zec7z6[11] & Fetov6);
assign Uvs7v6 = (~(Ytfxx6 & Fufxx6));
assign Fufxx6 = (~(Mufxx6 & Ktfxx6));
assign Mufxx6 = (Osd7z6[1] & Vs9ov6);
assign Ytfxx6 = (~(Tufxx6 & Rem7x6));
assign Rem7x6 = (~(Bsrov6 | Jbd8x6));
assign Bsrov6 = (!Yxd7z6[0]);
assign Yxd7z6[0] = (Btpiw6 & N3onv6);
assign Tufxx6 = (Gginv6 & Fetov6);
assign Nvs7v6 = (Pkkiw6 ? N6znv6 : Avfxx6);
assign Avfxx6 = (!W977z6);
assign Gvs7v6 = (!Hvfxx6);
assign Hvfxx6 = (Tqoov6 ? Gt67z6 : Ovfxx6);
assign Zus7v6 = (!Vvfxx6);
assign Vvfxx6 = (As9ov6 ? Wt67z6 : Ovfxx6);
assign Ovfxx6 = (!Y1znv6);
assign Sus7v6 = (Tqoov6 ? Cwfxx6 : Jxynv6);
assign Cwfxx6 = (!Mu67z6);
assign Lus7v6 = (As9ov6 ? Jwfxx6 : Jxynv6);
assign Jwfxx6 = (!Cv67z6);
assign Eus7v6 = (Pkkiw6 ? Usynv6 : Qwfxx6);
assign Qwfxx6 = (!Sv67z6);
assign Xts7v6 = (Klkiw6 ? Usynv6 : Xwfxx6);
assign Xwfxx6 = (!Iw67z6);
assign Qts7v6 = (Pkkiw6 ? Foynv6 : Exfxx6);
assign Exfxx6 = (!Yw67z6);
assign Jts7v6 = (Klkiw6 ? Foynv6 : Lxfxx6);
assign Lxfxx6 = (!Ox67z6);
assign Cts7v6 = (Pkkiw6 ? Qjynv6 : Sxfxx6);
assign Sxfxx6 = (!Ey67z6);
assign Vss7v6 = (Klkiw6 ? Qjynv6 : Zxfxx6);
assign Zxfxx6 = (!Uy67z6);
assign Oss7v6 = (Pkkiw6 ? Bfynv6 : Gyfxx6);
assign Gyfxx6 = (!Kz67z6);
assign Hss7v6 = (Klkiw6 ? Bfynv6 : Nyfxx6);
assign Nyfxx6 = (!A077z6);
assign Ass7v6 = (Pkkiw6 ? Maynv6 : Uyfxx6);
assign Uyfxx6 = (!Q077z6);
assign Trs7v6 = (Klkiw6 ? Maynv6 : Bzfxx6);
assign Bzfxx6 = (!G177z6);
assign Mrs7v6 = (Pkkiw6 ? P9xnv6 : Izfxx6);
assign Izfxx6 = (!W177z6);
assign Frs7v6 = (Klkiw6 ? P9xnv6 : Pzfxx6);
assign Pzfxx6 = (!M277z6);
assign Yqs7v6 = (!Wzfxx6);
assign Wzfxx6 = (Pkkiw6 ? D0gxx6 : C377z6);
assign Rqs7v6 = (!K0gxx6);
assign K0gxx6 = (Klkiw6 ? D0gxx6 : S377z6);
assign D0gxx6 = (!W1ynv6);
assign Kqs7v6 = (!R0gxx6);
assign R0gxx6 = (Pkkiw6 ? Y0gxx6 : I477z6);
assign Dqs7v6 = (!F1gxx6);
assign F1gxx6 = (Klkiw6 ? Y0gxx6 : Y477z6);
assign Y0gxx6 = (!Hxxnv6);
assign Wps7v6 = (Pkkiw6 ? Ssxnv6 : M1gxx6);
assign M1gxx6 = (!O577z6);
assign Pps7v6 = (Klkiw6 ? Ssxnv6 : T1gxx6);
assign T1gxx6 = (!E677z6);
assign Ips7v6 = (Pkkiw6 ? Doxnv6 : A2gxx6);
assign A2gxx6 = (!U677z6);
assign Bps7v6 = (Klkiw6 ? Doxnv6 : H2gxx6);
assign H2gxx6 = (!K777z6);
assign Uos7v6 = (Pkkiw6 ? Ojxnv6 : O2gxx6);
assign O2gxx6 = (!A877z6);
assign Nos7v6 = (Klkiw6 ? Ojxnv6 : V2gxx6);
assign V2gxx6 = (!Q877z6);
assign Gos7v6 = (Pkkiw6 ? Zexnv6 : C3gxx6);
assign C3gxx6 = (!G977z6);
assign Zns7v6 = (Mr9ov6 ? Bvtet6 : J3gxx6);
assign J3gxx6 = (Q3gxx6 | Rekiw6);
assign Rekiw6 = (X3gxx6 & Nh1ft6);
assign X3gxx6 = (Rr1ft6 & E4gxx6);
assign Q3gxx6 = (Pdkiw6 | Ogkiw6);
assign Sns7v6 = (Mr9ov6 ? Attet6 : L4gxx6);
assign L4gxx6 = (Pdkiw6 | Kekiw6);
assign Kekiw6 = (S4gxx6 & Z4gxx6);
assign Pdkiw6 = (G5gxx6 & N5gxx6);
assign N5gxx6 = (Xo1ft6 & U5gxx6);
assign G5gxx6 = (Z4gxx6 & Rf1ft6);
assign Lns7v6 = (Mr9ov6 ? Zqtet6 : B6gxx6);
assign B6gxx6 = (Ogkiw6 | Hgkiw6);
assign Hgkiw6 = (I6gxx6 & P6gxx6);
assign P6gxx6 = (W6gxx6 & U5gxx6);
assign I6gxx6 = (D7gxx6 & Z4gxx6);
assign Ens7v6 = (S3eiw6 ? T52iw6 : K6uet6);
assign S3eiw6 = (K7gxx6 & R7gxx6);
assign R7gxx6 = (~(Y7gxx6 & F8gxx6));
assign F8gxx6 = (Pp9ov6 & Wp9ov6);
assign Pp9ov6 = (~(Hryet6 | Woyet6));
assign Y7gxx6 = (M8gxx6 & T8gxx6);
assign M8gxx6 = (A9gxx6 & Qakiw6);
assign K7gxx6 = (Yjonv6 & O1eiw6);
assign Xms7v6 = (~(H9gxx6 & O9gxx6));
assign O9gxx6 = (~(Wzxet6 & B32iw6));
assign Qms7v6 = (V9gxx6 | Cagxx6);
assign Cagxx6 = (Jagxx6 & Qagxx6);
assign Qagxx6 = (Xagxx6 | Wlvet6);
assign Xagxx6 = (~(Cfxet6 | Ebgxx6));
assign Ebgxx6 = (!Yca7z6);
assign V9gxx6 = (Sbgxx6 ? Tim7z6[7] : Lbgxx6);
assign Lbgxx6 = (~(Zbgxx6 & Gcgxx6));
assign Gcgxx6 = (~(Fs1ov6 & Itb7z6[7]));
assign Zbgxx6 = (Ncgxx6 & Ucgxx6);
assign Ucgxx6 = (~(At1ov6 & Yca7z6));
assign Ncgxx6 = (~(Kwp7x6 & Ot1ov6));
assign Jms7v6 = (Bdgxx6 | Idgxx6);
assign Idgxx6 = (Jagxx6 & Pdgxx6);
assign Pdgxx6 = (Wdgxx6 | Xnvet6);
assign Wdgxx6 = (~(Dhxet6 | Degxx6));
assign Degxx6 = (!Gda7z6);
assign Bdgxx6 = (Sbgxx6 ? Tim7z6[6] : Kegxx6);
assign Kegxx6 = (~(Regxx6 & Yegxx6));
assign Yegxx6 = (~(Fs1ov6 & Itb7z6[6]));
assign Regxx6 = (Ffgxx6 & Mfgxx6);
assign Mfgxx6 = (~(At1ov6 & Gda7z6));
assign Ffgxx6 = (~(Lzq7x6 & Ot1ov6));
assign Cms7v6 = (Tfgxx6 | Aggxx6);
assign Aggxx6 = (Jagxx6 & Hggxx6);
assign Hggxx6 = (Oggxx6 | Ypvet6);
assign Oggxx6 = (~(Ejxet6 | Vggxx6));
assign Vggxx6 = (!Oda7z6);
assign Tfgxx6 = (Sbgxx6 ? Tim7z6[5] : Chgxx6);
assign Chgxx6 = (~(Jhgxx6 & Qhgxx6));
assign Qhgxx6 = (~(Fs1ov6 & Itb7z6[5]));
assign Jhgxx6 = (Xhgxx6 & Eigxx6);
assign Eigxx6 = (~(At1ov6 & Oda7z6));
assign Xhgxx6 = (~(Zsq7x6 & Ot1ov6));
assign Vls7v6 = (Ligxx6 | Sigxx6);
assign Sigxx6 = (Jagxx6 & Zigxx6);
assign Zigxx6 = (Gjgxx6 | Zrvet6);
assign Gjgxx6 = (~(Flxet6 | Njgxx6));
assign Njgxx6 = (!Qco7v6);
assign Ligxx6 = (Sbgxx6 ? Tim7z6[4] : Ujgxx6);
assign Ujgxx6 = (~(Bkgxx6 & Ikgxx6));
assign Ikgxx6 = (~(Fs1ov6 & Itb7z6[4]));
assign Bkgxx6 = (Pkgxx6 & Wkgxx6);
assign Wkgxx6 = (~(At1ov6 & Qco7v6));
assign Pkgxx6 = (~(Pnq7x6 & Ot1ov6));
assign Ols7v6 = (Dlgxx6 | Klgxx6);
assign Klgxx6 = (Jagxx6 & Rlgxx6);
assign Rlgxx6 = (Ylgxx6 | Auvet6);
assign Ylgxx6 = (Fmgxx6 & Wda7z6);
assign Fmgxx6 = (!Gnxet6);
assign Dlgxx6 = (Sbgxx6 ? Tim7z6[3] : Mmgxx6);
assign Mmgxx6 = (~(Tmgxx6 & Angxx6));
assign Angxx6 = (~(Fs1ov6 & Itb7z6[3]));
assign Tmgxx6 = (Hngxx6 & Ongxx6);
assign Ongxx6 = (~(At1ov6 & Wda7z6));
assign Hngxx6 = (~(Fiq7x6 & Ot1ov6));
assign Hls7v6 = (~(Vngxx6 & Cogxx6));
assign Cogxx6 = (~(Jagxx6 & Jogxx6));
assign Jogxx6 = (Qogxx6 | Bwvet6);
assign Qogxx6 = (Xogxx6 & Eea7z6);
assign Xogxx6 = (!Hpxet6);
assign Vngxx6 = (Sbgxx6 ? Lpgxx6 : Epgxx6);
assign Lpgxx6 = (!Tim7z6[2]);
assign Epgxx6 = (Spgxx6 & Zpgxx6);
assign Zpgxx6 = (~(Fs1ov6 & Itb7z6[2]));
assign Spgxx6 = (Gqgxx6 & Nqgxx6);
assign Nqgxx6 = (~(At1ov6 & Eea7z6));
assign Gqgxx6 = (~(Vcq7x6 & Ot1ov6));
assign Als7v6 = (Uqgxx6 | Brgxx6);
assign Brgxx6 = (Jagxx6 & Irgxx6);
assign Irgxx6 = (Prgxx6 | Cyvet6);
assign Prgxx6 = (~(Irxet6 | Wrgxx6));
assign Wrgxx6 = (!Mea7z6);
assign Uqgxx6 = (Sbgxx6 ? Tim7z6[1] : Dsgxx6);
assign Dsgxx6 = (~(Ksgxx6 & Rsgxx6));
assign Rsgxx6 = (~(Fs1ov6 & Itb7z6[1]));
assign Ksgxx6 = (Ysgxx6 & Ftgxx6);
assign Ftgxx6 = (~(At1ov6 & Mea7z6));
assign Ysgxx6 = (~(L7q7x6 & Ot1ov6));
assign Tks7v6 = (Mtgxx6 | Ttgxx6);
assign Ttgxx6 = (Jagxx6 & Augxx6);
assign Augxx6 = (Hugxx6 | D0wet6);
assign Hugxx6 = (~(Jtxet6 | Ougxx6));
assign Ougxx6 = (!Uea7z6);
assign Jagxx6 = (~(Vugxx6 | Sbgxx6));
assign Mtgxx6 = (Sbgxx6 ? Tim7z6[0] : Cvgxx6);
assign Cvgxx6 = (~(Jvgxx6 & Qvgxx6));
assign Qvgxx6 = (~(I8r7x6 & Xvgxx6));
assign Jvgxx6 = (Ewgxx6 & Lwgxx6);
assign Lwgxx6 = (~(Znn7z6[1] & Asonv6));
assign Asonv6 = (~(Swgxx6 & Zwgxx6));
assign Zwgxx6 = (~(Styet6 & I8r7x6));
assign Swgxx6 = (~(Ewyet6 & Itb7z6[0]));
assign Ewgxx6 = (~(At1ov6 & Uea7z6));
assign Mks7v6 = (Gxgxx6 | Nxgxx6);
assign Nxgxx6 = (Uxgxx6 & Bygxx6);
assign Bygxx6 = (Iygxx6 | O5vet6);
assign Iygxx6 = (~(Uywet6 | Pygxx6));
assign Pygxx6 = (!Uaa7z6);
assign Gxgxx6 = (Dzgxx6 ? Wygxx6 : Tim7z6[15]);
assign Wygxx6 = (~(Kzgxx6 & Rzgxx6));
assign Rzgxx6 = (~(Fs1ov6 & Itb7z6[15]));
assign Kzgxx6 = (Yzgxx6 & F0hxx6);
assign F0hxx6 = (~(At1ov6 & Uaa7z6));
assign Yzgxx6 = (~(Oyp7x6 & Ot1ov6));
assign Fks7v6 = (M0hxx6 | T0hxx6);
assign T0hxx6 = (Uxgxx6 & A1hxx6);
assign A1hxx6 = (H1hxx6 | P7vet6);
assign H1hxx6 = (~(V0xet6 | O1hxx6));
assign O1hxx6 = (!Cba7z6);
assign M0hxx6 = (Dzgxx6 ? V1hxx6 : Tim7z6[14]);
assign V1hxx6 = (~(C2hxx6 & J2hxx6));
assign J2hxx6 = (~(Fs1ov6 & Itb7z6[14]));
assign C2hxx6 = (Q2hxx6 & X2hxx6);
assign X2hxx6 = (~(At1ov6 & Cba7z6));
assign Q2hxx6 = (~(Twq7x6 & Ot1ov6));
assign Yjs7v6 = (E3hxx6 | L3hxx6);
assign L3hxx6 = (Uxgxx6 & S3hxx6);
assign S3hxx6 = (Z3hxx6 | Q9vet6);
assign Z3hxx6 = (~(W2xet6 | G4hxx6));
assign G4hxx6 = (!Kba7z6);
assign E3hxx6 = (Dzgxx6 ? N4hxx6 : Tim7z6[13]);
assign N4hxx6 = (~(U4hxx6 & B5hxx6));
assign B5hxx6 = (~(Fs1ov6 & Itb7z6[13]));
assign U4hxx6 = (I5hxx6 & P5hxx6);
assign P5hxx6 = (~(At1ov6 & Kba7z6));
assign I5hxx6 = (~(Vqq7x6 & Ot1ov6));
assign Rjs7v6 = (W5hxx6 | D6hxx6);
assign D6hxx6 = (Uxgxx6 & K6hxx6);
assign K6hxx6 = (R6hxx6 | Rbvet6);
assign R6hxx6 = (~(X4xet6 | Y6hxx6));
assign Y6hxx6 = (!Jco7v6);
assign W5hxx6 = (Dzgxx6 ? F7hxx6 : Tim7z6[12]);
assign F7hxx6 = (~(M7hxx6 & T7hxx6));
assign T7hxx6 = (~(Fs1ov6 & Itb7z6[12]));
assign M7hxx6 = (A8hxx6 & H8hxx6);
assign H8hxx6 = (~(At1ov6 & Jco7v6));
assign A8hxx6 = (~(Llq7x6 & Ot1ov6));
assign Kjs7v6 = (O8hxx6 | V8hxx6);
assign V8hxx6 = (Uxgxx6 & C9hxx6);
assign C9hxx6 = (J9hxx6 | Sdvet6);
assign J9hxx6 = (Q9hxx6 & Sba7z6);
assign Q9hxx6 = (!Y6xet6);
assign O8hxx6 = (Dzgxx6 ? X9hxx6 : Tim7z6[11]);
assign X9hxx6 = (~(Eahxx6 & Lahxx6));
assign Lahxx6 = (~(Fs1ov6 & Itb7z6[11]));
assign Eahxx6 = (Sahxx6 & Zahxx6);
assign Zahxx6 = (~(At1ov6 & Sba7z6));
assign Sahxx6 = (~(Bgq7x6 & Ot1ov6));
assign Djs7v6 = (~(Gbhxx6 & Nbhxx6));
assign Nbhxx6 = (~(Uxgxx6 & Ubhxx6));
assign Ubhxx6 = (Bchxx6 | Tfvet6);
assign Bchxx6 = (Ichxx6 & Aca7z6);
assign Ichxx6 = (!Z8xet6);
assign Gbhxx6 = (Dzgxx6 ? Wchxx6 : Pchxx6);
assign Wchxx6 = (Ddhxx6 & Kdhxx6);
assign Kdhxx6 = (~(Fs1ov6 & Itb7z6[10]));
assign Ddhxx6 = (Rdhxx6 & Ydhxx6);
assign Ydhxx6 = (~(At1ov6 & Aca7z6));
assign Rdhxx6 = (~(Raq7x6 & Ot1ov6));
assign Pchxx6 = (!Tim7z6[10]);
assign Wis7v6 = (Fehxx6 | Mehxx6);
assign Mehxx6 = (Uxgxx6 & Tehxx6);
assign Tehxx6 = (Afhxx6 | Uhvet6);
assign Afhxx6 = (~(Abxet6 | Hfhxx6));
assign Hfhxx6 = (!Ica7z6);
assign Fehxx6 = (Dzgxx6 ? Ofhxx6 : Tim7z6[9]);
assign Ofhxx6 = (~(Vfhxx6 & Cghxx6));
assign Cghxx6 = (~(Fs1ov6 & Itb7z6[9]));
assign Vfhxx6 = (Jghxx6 & Qghxx6);
assign Qghxx6 = (~(At1ov6 & Ica7z6));
assign Jghxx6 = (~(H5q7x6 & Ot1ov6));
assign Pis7v6 = (Xghxx6 | Ehhxx6);
assign Ehhxx6 = (Uxgxx6 & Lhhxx6);
assign Lhhxx6 = (Shhxx6 | Vjvet6);
assign Shhxx6 = (~(Bdxet6 | Zhhxx6));
assign Zhhxx6 = (!Qca7z6);
assign Uxgxx6 = (Znn7z6[2] & Dzgxx6);
assign Xghxx6 = (Dzgxx6 ? Gihxx6 : Tim7z6[8]);
assign Dzgxx6 = (~(Sbgxx6 & Nihxx6));
assign Nihxx6 = (~(Uihxx6 & Eia7z6));
assign Uihxx6 = (Bjhxx6 & Ijhxx6);
assign Sbgxx6 = (Pjhxx6 & Wjhxx6);
assign Pjhxx6 = (Dkhxx6 & Kkhxx6);
assign Dkhxx6 = (~(Rkhxx6 & Ykhxx6));
assign Rkhxx6 = (Djonv6 & Mia7z6);
assign Gihxx6 = (~(Flhxx6 & Mlhxx6));
assign Mlhxx6 = (~(Fs1ov6 & Itb7z6[8]));
assign Flhxx6 = (Tlhxx6 & Amhxx6);
assign Amhxx6 = (~(At1ov6 & Qca7z6));
assign Tlhxx6 = (~(Kqonv6 & Ot1ov6));
assign Iis7v6 = (Hmhxx6 | Omhxx6);
assign Omhxx6 = (Vmhxx6 & Cnhxx6);
assign Cnhxx6 = (Jnhxx6 | Gpuet6);
assign Jnhxx6 = (~(Miwet6 | Qnhxx6));
assign Qnhxx6 = (!Q8a7z6);
assign Hmhxx6 = (Eohxx6 ? Xnhxx6 : Tim7z6[23]);
assign Xnhxx6 = (~(Lohxx6 & Sohxx6));
assign Sohxx6 = (~(Fs1ov6 & Itb7z6[23]));
assign Lohxx6 = (Zohxx6 & Gphxx6);
assign Gphxx6 = (~(At1ov6 & Q8a7z6));
assign Zohxx6 = (~(Xzp7x6 & Ot1ov6));
assign Bis7v6 = (Nphxx6 | Uphxx6);
assign Uphxx6 = (Vmhxx6 & Bqhxx6);
assign Bqhxx6 = (Iqhxx6 | Hruet6);
assign Iqhxx6 = (~(Nkwet6 | Pqhxx6));
assign Pqhxx6 = (!Y8a7z6);
assign Nphxx6 = (Eohxx6 ? Wqhxx6 : Tim7z6[22]);
assign Wqhxx6 = (~(Drhxx6 & Krhxx6));
assign Krhxx6 = (~(Fs1ov6 & Itb7z6[22]));
assign Drhxx6 = (Rrhxx6 & Yrhxx6);
assign Yrhxx6 = (~(At1ov6 & Y8a7z6));
assign Rrhxx6 = (~(Wuq7x6 & Ot1ov6));
assign Uhs7v6 = (Fshxx6 | Mshxx6);
assign Mshxx6 = (Vmhxx6 & Tshxx6);
assign Tshxx6 = (Athxx6 | Ituet6);
assign Athxx6 = (~(Omwet6 | Hthxx6));
assign Hthxx6 = (!G9a7z6);
assign Fshxx6 = (Eohxx6 ? Othxx6 : Tim7z6[21]);
assign Othxx6 = (~(Vthxx6 & Cuhxx6));
assign Cuhxx6 = (~(Fs1ov6 & Itb7z6[21]));
assign Vthxx6 = (Juhxx6 & Quhxx6);
assign Quhxx6 = (~(At1ov6 & G9a7z6));
assign Juhxx6 = (~(Mpq7x6 & Ot1ov6));
assign Nhs7v6 = (Xuhxx6 | Evhxx6);
assign Evhxx6 = (Vmhxx6 & Lvhxx6);
assign Lvhxx6 = (Svhxx6 | Jvuet6);
assign Svhxx6 = (~(Powet6 | Zvhxx6));
assign Zvhxx6 = (!Cco7v6);
assign Xuhxx6 = (Eohxx6 ? Gwhxx6 : Tim7z6[20]);
assign Gwhxx6 = (~(Nwhxx6 & Uwhxx6));
assign Uwhxx6 = (~(Fs1ov6 & Itb7z6[20]));
assign Nwhxx6 = (Bxhxx6 & Ixhxx6);
assign Ixhxx6 = (~(At1ov6 & Cco7v6));
assign Bxhxx6 = (~(Ckq7x6 & Ot1ov6));
assign Ghs7v6 = (Pxhxx6 | Wxhxx6);
assign Wxhxx6 = (Vmhxx6 & Dyhxx6);
assign Dyhxx6 = (Kyhxx6 | Kxuet6);
assign Kyhxx6 = (Ryhxx6 & O9a7z6);
assign Ryhxx6 = (!Qqwet6);
assign Pxhxx6 = (Eohxx6 ? Yyhxx6 : Tim7z6[19]);
assign Yyhxx6 = (~(Fzhxx6 & Mzhxx6));
assign Mzhxx6 = (~(Fs1ov6 & Itb7z6[19]));
assign Fzhxx6 = (Tzhxx6 & A0ixx6);
assign A0ixx6 = (~(At1ov6 & O9a7z6));
assign Tzhxx6 = (~(Seq7x6 & Ot1ov6));
assign Zgs7v6 = (~(H0ixx6 & O0ixx6));
assign O0ixx6 = (~(Vmhxx6 & V0ixx6));
assign V0ixx6 = (C1ixx6 | Lzuet6);
assign C1ixx6 = (J1ixx6 & W9a7z6);
assign J1ixx6 = (!Rswet6);
assign H0ixx6 = (Eohxx6 ? X1ixx6 : Q1ixx6);
assign X1ixx6 = (E2ixx6 & L2ixx6);
assign L2ixx6 = (~(Fs1ov6 & Itb7z6[18]));
assign E2ixx6 = (S2ixx6 & Z2ixx6);
assign Z2ixx6 = (~(At1ov6 & W9a7z6));
assign S2ixx6 = (~(I9q7x6 & Ot1ov6));
assign Q1ixx6 = (!Tim7z6[18]);
assign Sgs7v6 = (G3ixx6 | N3ixx6);
assign N3ixx6 = (Vmhxx6 & U3ixx6);
assign U3ixx6 = (B4ixx6 | M1vet6);
assign B4ixx6 = (~(Suwet6 | I4ixx6));
assign I4ixx6 = (!Eaa7z6);
assign G3ixx6 = (Eohxx6 ? P4ixx6 : Tim7z6[17]);
assign P4ixx6 = (~(W4ixx6 & D5ixx6));
assign D5ixx6 = (~(Fs1ov6 & Itb7z6[17]));
assign W4ixx6 = (K5ixx6 & R5ixx6);
assign R5ixx6 = (~(At1ov6 & Eaa7z6));
assign K5ixx6 = (~(Y3q7x6 & Ot1ov6));
assign Lgs7v6 = (Y5ixx6 | F6ixx6);
assign F6ixx6 = (Vmhxx6 & M6ixx6);
assign M6ixx6 = (T6ixx6 | N3vet6);
assign T6ixx6 = (~(Twwet6 | A7ixx6));
assign A7ixx6 = (!Maa7z6);
assign Vmhxx6 = (Znn7z6[2] & Eohxx6);
assign Y5ixx6 = (Eohxx6 ? H7ixx6 : Tim7z6[16]);
assign Eohxx6 = (~(O7ixx6 & V7ixx6));
assign V7ixx6 = (~(C8ixx6 & J8ixx6));
assign J8ixx6 = (Q8ixx6 & Ijhxx6);
assign C8ixx6 = (Bjhxx6 & Ven7z6[0]);
assign H7ixx6 = (~(X8ixx6 & E9ixx6));
assign E9ixx6 = (~(Fs1ov6 & Itb7z6[16]));
assign X8ixx6 = (L9ixx6 & S9ixx6);
assign S9ixx6 = (~(At1ov6 & Maa7z6));
assign L9ixx6 = (~(V4r7x6 & Ot1ov6));
assign Egs7v6 = (Z9ixx6 | Gaixx6);
assign Gaixx6 = (Bq1ov6 & Naixx6);
assign Naixx6 = (Uaixx6 | Zauet6);
assign Uaixx6 = (~(F4wet6 | Bbixx6));
assign Bbixx6 = (!M6a7z6);
assign Z9ixx6 = (Kr1ov6 ? Ibixx6 : Tim7z6[30]);
assign Ibixx6 = (~(Pbixx6 & Wbixx6));
assign Wbixx6 = (~(Fs1ov6 & Itb7z6[30]));
assign Pbixx6 = (Dcixx6 & Kcixx6);
assign Kcixx6 = (~(At1ov6 & M6a7z6));
assign Dcixx6 = (~(Vxq7x6 & Ot1ov6));
assign Xfs7v6 = (Rcixx6 | Ycixx6);
assign Ycixx6 = (Bq1ov6 & Fdixx6);
assign Fdixx6 = (Mdixx6 | Aduet6);
assign Mdixx6 = (~(G6wet6 | Tdixx6));
assign Tdixx6 = (!U6a7z6);
assign Rcixx6 = (Kr1ov6 ? Aeixx6 : Tim7z6[29]);
assign Aeixx6 = (~(Heixx6 & Oeixx6));
assign Oeixx6 = (~(Fs1ov6 & Itb7z6[29]));
assign Heixx6 = (Veixx6 & Cfixx6);
assign Cfixx6 = (~(At1ov6 & U6a7z6));
assign Veixx6 = (~(Qrq7x6 & Ot1ov6));
assign Qfs7v6 = (Jfixx6 | Qfixx6);
assign Qfixx6 = (Bq1ov6 & Xfixx6);
assign Xfixx6 = (Egixx6 | Bfuet6);
assign Egixx6 = (~(H8wet6 | Lgixx6));
assign Lgixx6 = (!C7a7z6);
assign Jfixx6 = (Kr1ov6 ? Sgixx6 : Tim7z6[28]);
assign Sgixx6 = (~(Zgixx6 & Ghixx6));
assign Ghixx6 = (~(Fs1ov6 & Itb7z6[28]));
assign Zgixx6 = (Nhixx6 & Uhixx6);
assign Uhixx6 = (~(At1ov6 & C7a7z6));
assign Nhixx6 = (~(Gmq7x6 & Ot1ov6));
assign Jfs7v6 = (Biixx6 | Iiixx6);
assign Iiixx6 = (Bq1ov6 & Piixx6);
assign Piixx6 = (Wiixx6 | Chuet6);
assign Wiixx6 = (~(Iawet6 | Djixx6));
assign Djixx6 = (!K7a7z6);
assign Biixx6 = (Kr1ov6 ? Kjixx6 : Tim7z6[27]);
assign Kjixx6 = (~(Rjixx6 & Yjixx6));
assign Yjixx6 = (~(Fs1ov6 & Itb7z6[27]));
assign Rjixx6 = (Fkixx6 & Mkixx6);
assign Mkixx6 = (~(At1ov6 & K7a7z6));
assign Fkixx6 = (~(Wgq7x6 & Ot1ov6));
assign Cfs7v6 = (~(Tkixx6 & Alixx6));
assign Alixx6 = (~(Bq1ov6 & Hlixx6));
assign Hlixx6 = (Olixx6 | Djuet6);
assign Olixx6 = (Vlixx6 & S7a7z6);
assign Vlixx6 = (!Jcwet6);
assign Tkixx6 = (Kr1ov6 ? Jmixx6 : Cmixx6);
assign Jmixx6 = (Qmixx6 & Xmixx6);
assign Xmixx6 = (~(Fs1ov6 & Itb7z6[26]));
assign Qmixx6 = (Enixx6 & Lnixx6);
assign Lnixx6 = (~(At1ov6 & S7a7z6));
assign Enixx6 = (~(Mbq7x6 & Ot1ov6));
assign Cmixx6 = (!Tim7z6[26]);
assign Ves7v6 = (Snixx6 | Znixx6);
assign Znixx6 = (Bq1ov6 & Goixx6);
assign Goixx6 = (Noixx6 | Eluet6);
assign Noixx6 = (~(Kewet6 | Uoixx6));
assign Uoixx6 = (!A8a7z6);
assign Snixx6 = (Kr1ov6 ? Bpixx6 : Tim7z6[25]);
assign Bpixx6 = (~(Ipixx6 & Ppixx6));
assign Ppixx6 = (~(Fs1ov6 & Itb7z6[25]));
assign Ipixx6 = (Wpixx6 & Dqixx6);
assign Dqixx6 = (~(At1ov6 & A8a7z6));
assign Wpixx6 = (~(C6q7x6 & Ot1ov6));
assign Oes7v6 = (Kqixx6 | Rqixx6);
assign Rqixx6 = (Bq1ov6 & Yqixx6);
assign Yqixx6 = (Frixx6 | Fnuet6);
assign Frixx6 = (~(Lgwet6 | Mrixx6));
assign Mrixx6 = (!I8a7z6);
assign Bq1ov6 = (Znn7z6[2] & Kr1ov6);
assign Kqixx6 = (Kr1ov6 ? Trixx6 : Tim7z6[24]);
assign Kr1ov6 = (~(O7ixx6 & Asixx6));
assign Asixx6 = (~(Hsixx6 & Bjhxx6));
assign Hsixx6 = (~(Eia7z6 | Wzxet6));
assign Eia7z6 = (Osixx6 & Vsixx6);
assign Vsixx6 = (~(Ven7z6[2] & Ven7z6[1]));
assign O7ixx6 = (Ctixx6 & Wjhxx6);
assign Wjhxx6 = (Jtixx6 & H9gxx6);
assign H9gxx6 = (~(B32iw6 & Qtixx6));
assign B32iw6 = (!O1eiw6);
assign Jtixx6 = (~(Ijhxx6 & Xtixx6));
assign Xtixx6 = (~(Euixx6 & Luixx6));
assign Euixx6 = (~(Suixx6 & Cmonv6));
assign Cmonv6 = (Bp9ov6 ? Zuixx6 : Goonv6);
assign Bp9ov6 = (!L3eiw6);
assign L3eiw6 = (~(Gvixx6 & Nvixx6));
assign Gvixx6 = (Uvixx6 & Bwixx6);
assign Ctixx6 = (Iwixx6 & Kkhxx6);
assign Kkhxx6 = (~(Pwixx6 & Bjhxx6));
assign Pwixx6 = (I2yet6 & Ijhxx6);
assign Iwixx6 = (~(Wwixx6 & Ykhxx6));
assign Ykhxx6 = (Dxixx6 & Kxixx6);
assign Dxixx6 = (Rxixx6 & Ijhxx6);
assign Ijhxx6 = (!Wzxet6);
assign Wwixx6 = (Djonv6 & Kjonv6);
assign Kjonv6 = (!Mia7z6);
assign Mia7z6 = (Yxixx6 | Ven7z6[0]);
assign Trixx6 = (~(Fyixx6 & Myixx6));
assign Myixx6 = (~(Fs1ov6 & Itb7z6[24]));
assign Fs1ov6 = (Tyixx6 & I2yet6);
assign Tyixx6 = (Ewyet6 & Znn7z6[1]);
assign Fyixx6 = (Azixx6 & Hzixx6);
assign Hzixx6 = (~(At1ov6 & I8a7z6));
assign At1ov6 = (Rxixx6 ? Ozixx6 : Kxixx6);
assign Azixx6 = (~(Yqonv6 & Ot1ov6));
assign Ot1ov6 = (~(Znn7z6[3] & Vzixx6));
assign Vzixx6 = (~(C0jxx6 & I2yet6));
assign C0jxx6 = (Styet6 & Znn7z6[1]);
assign Hes7v6 = (Mk9ov6 ? Kyn7z6[2] : J0jxx6);
assign Mk9ov6 = (~(H6l8v6 | Gazet6));
assign H6l8v6 = (HTRANSS[1] & Zuixx6);
assign Aes7v6 = (~(Q0jxx6 & X0jxx6));
assign X0jxx6 = (~(E1jxx6 & L1jxx6));
assign E1jxx6 = (~(Cfonv6 | S1jxx6));
assign Q0jxx6 = (~(Z1jxx6 & Svn7z6[0]));
assign Tds7v6 = (~(G2jxx6 & N2jxx6));
assign N2jxx6 = (~(U2jxx6 & L1jxx6));
assign U2jxx6 = (~(Zn9ov6 | S1jxx6));
assign G2jxx6 = (~(Svn7z6[1] & Z1jxx6));
assign Mds7v6 = (~(B3jxx6 & I3jxx6));
assign I3jxx6 = (P3jxx6 | W3jxx6);
assign B3jxx6 = (D4jxx6 & K4jxx6);
assign K4jxx6 = (~(L1jxx6 & J0jxx6));
assign L1jxx6 = (HWRITES & W3jxx6);
assign W3jxx6 = (!Z1jxx6);
assign Z1jxx6 = (~(R4jxx6 | HREADYS));
assign R4jxx6 = (!Y4jxx6);
assign D4jxx6 = (~(S1jxx6 & HWRITES));
assign S1jxx6 = (~(Y4jxx6 | HREADYS));
assign Y4jxx6 = (~(Svn7z6[0] & Qtixx6));
assign Fds7v6 = (U0jhw6 ? R3h7z6[1] : F5jxx6);
assign U0jhw6 = (G0jhw6 & M5jxx6);
assign M5jxx6 = (~(T5jxx6 & R3h7z6[0]));
assign T5jxx6 = (~(Ypinv6 | Bqmov6));
assign Bqmov6 = (A6jxx6 & K2d7x6);
assign A6jxx6 = (I3wnv6 & U3a7x6);
assign G0jhw6 = (~(H6jxx6 & Zpdiw6));
assign Zpdiw6 = (Ii9ov6 & Fsmov6);
assign Fsmov6 = (~(O6jxx6 & V6jxx6));
assign V6jxx6 = (~(Sv97x6 & C7jxx6));
assign O6jxx6 = (Iqmov6 & U3a7x6);
assign H6jxx6 = (Msmov6 & Bi9ov6);
assign Ycs7v6 = (~(J7jxx6 & Q7jxx6));
assign Q7jxx6 = (Hbpiw6 | X7jxx6);
assign X7jxx6 = (E8jxx6 & L8jxx6);
assign L8jxx6 = (~(S8jxx6 & Cmm7z6[0]));
assign E8jxx6 = (Z8jxx6 & G9jxx6);
assign G9jxx6 = (~(N9jxx6 & U9jxx6));
assign N9jxx6 = (~(Bajxx6 | R3ihw6));
assign R3ihw6 = (Iajxx6 & Pajxx6);
assign Pajxx6 = (Wajxx6 & Dbjxx6);
assign Dbjxx6 = (~(Kbjxx6 & Td9ov6));
assign Wajxx6 = (~(Rbjxx6 & Jf9ov6));
assign Iajxx6 = (Ybjxx6 & Fcjxx6);
assign Fcjxx6 = (~(Mcjxx6 & Ve9ov6));
assign Ybjxx6 = (~(Tcjxx6 & Fd9ov6));
assign Z8jxx6 = (Adjxx6 | I2bov6);
assign I2bov6 = (Hdjxx6 & Odjxx6);
assign Odjxx6 = (Vdjxx6 & Cejxx6);
assign Cejxx6 = (Jejxx6 & Qejxx6);
assign Qejxx6 = (Xejxx6 & Efjxx6);
assign Efjxx6 = (~(Lfjxx6 & Pic7z6[0]));
assign Xejxx6 = (~(Sfjxx6 & vis_r12_o[0]));
assign Jejxx6 = (Zfjxx6 & Ggjxx6);
assign Ggjxx6 = (~(Ngjxx6 & vis_r11_o[0]));
assign Zfjxx6 = (~(Ugjxx6 & vis_r10_o[0]));
assign Vdjxx6 = (Bhjxx6 & Ihjxx6);
assign Ihjxx6 = (~(Phjxx6 & vis_r8_o[0]));
assign Bhjxx6 = (Whjxx6 & Dijxx6);
assign Dijxx6 = (~(Kijxx6 & vis_r7_o[0]));
assign Whjxx6 = (~(Rijxx6 & vis_r9_o[0]));
assign Hdjxx6 = (Yijxx6 & Fjjxx6);
assign Fjjxx6 = (Mjjxx6 & Tjjxx6);
assign Tjjxx6 = (Akjxx6 & Hkjxx6);
assign Hkjxx6 = (~(Okjxx6 & vis_r6_o[0]));
assign Akjxx6 = (~(Vkjxx6 & vis_r5_o[0]));
assign Mjjxx6 = (Cljxx6 & Jljxx6);
assign Jljxx6 = (~(Qljxx6 & vis_r4_o[0]));
assign Cljxx6 = (~(Xljxx6 & vis_r3_o[0]));
assign Yijxx6 = (Emjxx6 & Lmjxx6);
assign Lmjxx6 = (~(Smjxx6 & vis_r1_o[0]));
assign Emjxx6 = (Zmjxx6 & Gnjxx6);
assign Gnjxx6 = (~(Nnjxx6 & vis_r0_o[0]));
assign Zmjxx6 = (~(Unjxx6 & vis_r2_o[0]));
assign J7jxx6 = (~(K1i7z6[0] & Zs4ov6));
assign Rcs7v6 = (~(Bojxx6 & Iojxx6));
assign Iojxx6 = (Hbpiw6 | Pojxx6);
assign Pojxx6 = (Wojxx6 & Dpjxx6);
assign Dpjxx6 = (Kpjxx6 & Rpjxx6);
assign Rpjxx6 = (~(Ypjxx6 & U9jxx6));
assign Ypjxx6 = (~(Bajxx6 | J5knv6));
assign J5knv6 = (Fqjxx6 & Mqjxx6);
assign Mqjxx6 = (Tqjxx6 & Arjxx6);
assign Arjxx6 = (~(Ex77x6 & Kbjxx6));
assign Tqjxx6 = (~(Ab67x6 & Rbjxx6));
assign Fqjxx6 = (Hrjxx6 & Orjxx6);
assign Orjxx6 = (~(Ob67x6 & Mcjxx6));
assign Hrjxx6 = (~(Vv77x6 & Tcjxx6));
assign Bajxx6 = (Vrjxx6 & Csjxx6);
assign Kpjxx6 = (Adjxx6 | Lu9ov6);
assign Lu9ov6 = (Jsjxx6 & Qsjxx6);
assign Qsjxx6 = (Xsjxx6 & Etjxx6);
assign Etjxx6 = (Ltjxx6 & Stjxx6);
assign Stjxx6 = (Ztjxx6 & Gujxx6);
assign Gujxx6 = (~(Lfjxx6 & Pic7z6[1]));
assign Ztjxx6 = (~(Sfjxx6 & vis_r12_o[1]));
assign Ltjxx6 = (Nujxx6 & Uujxx6);
assign Uujxx6 = (~(Ngjxx6 & vis_r11_o[1]));
assign Nujxx6 = (~(Ugjxx6 & vis_r10_o[1]));
assign Xsjxx6 = (Bvjxx6 & Ivjxx6);
assign Ivjxx6 = (~(Phjxx6 & vis_r8_o[1]));
assign Bvjxx6 = (Pvjxx6 & Wvjxx6);
assign Wvjxx6 = (~(Kijxx6 & vis_r7_o[1]));
assign Pvjxx6 = (~(Rijxx6 & vis_r9_o[1]));
assign Jsjxx6 = (Dwjxx6 & Kwjxx6);
assign Kwjxx6 = (Rwjxx6 & Ywjxx6);
assign Ywjxx6 = (Fxjxx6 & Mxjxx6);
assign Mxjxx6 = (~(Okjxx6 & vis_r6_o[1]));
assign Fxjxx6 = (~(Vkjxx6 & vis_r5_o[1]));
assign Rwjxx6 = (Txjxx6 & Ayjxx6);
assign Ayjxx6 = (~(Qljxx6 & vis_r4_o[1]));
assign Txjxx6 = (~(Xljxx6 & vis_r3_o[1]));
assign Dwjxx6 = (Hyjxx6 & Oyjxx6);
assign Oyjxx6 = (~(Smjxx6 & vis_r1_o[1]));
assign Hyjxx6 = (Vyjxx6 & Czjxx6);
assign Czjxx6 = (~(Nnjxx6 & vis_r0_o[1]));
assign Vyjxx6 = (~(Unjxx6 & vis_r2_o[1]));
assign Wojxx6 = (Jzjxx6 & Qzjxx6);
assign Qzjxx6 = (~(Xzjxx6 & vis_pc_o[1]));
assign Jzjxx6 = (~(S8jxx6 & Cmm7z6[1]));
assign Hbpiw6 = (~(E0kxx6 & L0kxx6));
assign L0kxx6 = (~(K0riw6 & S0kxx6));
assign S0kxx6 = (~(Prsov6 & T1riw6));
assign E0kxx6 = (Z0kxx6 & G1kxx6);
assign Bojxx6 = (~(K1i7z6[1] & Zs4ov6));
assign Kcs7v6 = (~(N1kxx6 & U1kxx6));
assign U1kxx6 = (B2kxx6 & I2kxx6);
assign I2kxx6 = (~(Xzjxx6 & vis_pc_o[2]));
assign B2kxx6 = (P2kxx6 & W2kxx6);
assign W2kxx6 = (~(U9jxx6 & Nmjnv6));
assign Nmjnv6 = (~(D3kxx6 & K3kxx6));
assign K3kxx6 = (R3kxx6 & Y3kxx6);
assign Y3kxx6 = (~(Kbjxx6 & Icfov6));
assign R3kxx6 = (~(Kdfov6 & Rbjxx6));
assign D3kxx6 = (F4kxx6 & M4kxx6);
assign M4kxx6 = (~(Ddfov6 & Mcjxx6));
assign F4kxx6 = (~(Tcjxx6 & Bcfov6));
assign P2kxx6 = (Adjxx6 | N5yiw6);
assign N5yiw6 = (T4kxx6 & A5kxx6);
assign A5kxx6 = (H5kxx6 & O5kxx6);
assign O5kxx6 = (V5kxx6 & C6kxx6);
assign C6kxx6 = (J6kxx6 & Q6kxx6);
assign Q6kxx6 = (~(X6kxx6 & vis_psp_o[2]));
assign J6kxx6 = (~(E7kxx6 & vis_msp_o[2]));
assign V5kxx6 = (L7kxx6 & S7kxx6);
assign S7kxx6 = (~(Lfjxx6 & Pic7z6[2]));
assign L7kxx6 = (~(Sfjxx6 & vis_r12_o[2]));
assign H5kxx6 = (Z7kxx6 & G8kxx6);
assign G8kxx6 = (N8kxx6 & U8kxx6);
assign U8kxx6 = (~(Ngjxx6 & vis_r11_o[2]));
assign N8kxx6 = (~(Ugjxx6 & vis_r10_o[2]));
assign Z7kxx6 = (B9kxx6 & I9kxx6);
assign I9kxx6 = (~(Kijxx6 & vis_r7_o[2]));
assign B9kxx6 = (~(Rijxx6 & vis_r9_o[2]));
assign T4kxx6 = (P9kxx6 & W9kxx6);
assign W9kxx6 = (Dakxx6 & Kakxx6);
assign Kakxx6 = (Rakxx6 & Yakxx6);
assign Yakxx6 = (~(Phjxx6 & vis_r8_o[2]));
assign Rakxx6 = (~(Okjxx6 & vis_r6_o[2]));
assign Dakxx6 = (Fbkxx6 & Mbkxx6);
assign Mbkxx6 = (~(Vkjxx6 & vis_r5_o[2]));
assign Fbkxx6 = (~(Qljxx6 & vis_r4_o[2]));
assign P9kxx6 = (Tbkxx6 & Ackxx6);
assign Ackxx6 = (Hckxx6 & Ockxx6);
assign Ockxx6 = (~(Xljxx6 & vis_r3_o[2]));
assign Hckxx6 = (~(Nnjxx6 & vis_r0_o[2]));
assign Tbkxx6 = (Vckxx6 & Cdkxx6);
assign Cdkxx6 = (~(Unjxx6 & vis_r2_o[2]));
assign Vckxx6 = (~(Smjxx6 & vis_r1_o[2]));
assign N1kxx6 = (Jdkxx6 & Qdkxx6);
assign Qdkxx6 = (~(S8jxx6 & Yefnv6));
assign Jdkxx6 = (~(K1i7z6[2] & Zs4ov6));
assign Dcs7v6 = (~(Xdkxx6 & Eekxx6));
assign Eekxx6 = (Lekxx6 & Sekxx6);
assign Sekxx6 = (~(U9jxx6 & Rhjnv6));
assign Rhjnv6 = (~(Zekxx6 & Gfkxx6));
assign Gfkxx6 = (Nfkxx6 & Ufkxx6);
assign Ufkxx6 = (~(Mmlov6 & Kbjxx6));
assign Nfkxx6 = (~(Onlov6 & Rbjxx6));
assign Zekxx6 = (Bgkxx6 & Igkxx6);
assign Igkxx6 = (~(Hnlov6 & Mcjxx6));
assign Bgkxx6 = (~(Fmlov6 & Tcjxx6));
assign Lekxx6 = (Pgkxx6 & Wgkxx6);
assign Pgkxx6 = (Adjxx6 | Zhh6x6);
assign Zhh6x6 = (Dhkxx6 & Khkxx6);
assign Khkxx6 = (Rhkxx6 & Yhkxx6);
assign Yhkxx6 = (Fikxx6 & Mikxx6);
assign Mikxx6 = (Tikxx6 & Ajkxx6);
assign Ajkxx6 = (~(X6kxx6 & vis_psp_o[3]));
assign Tikxx6 = (~(E7kxx6 & vis_msp_o[3]));
assign Fikxx6 = (Hjkxx6 & Ojkxx6);
assign Ojkxx6 = (~(Lfjxx6 & Pic7z6[3]));
assign Hjkxx6 = (~(Sfjxx6 & vis_r12_o[3]));
assign Rhkxx6 = (Vjkxx6 & Ckkxx6);
assign Ckkxx6 = (Jkkxx6 & Qkkxx6);
assign Qkkxx6 = (~(Ngjxx6 & vis_r11_o[3]));
assign Jkkxx6 = (~(Ugjxx6 & vis_r10_o[3]));
assign Vjkxx6 = (Xkkxx6 & Elkxx6);
assign Elkxx6 = (~(Kijxx6 & vis_r7_o[3]));
assign Xkkxx6 = (~(Rijxx6 & vis_r9_o[3]));
assign Dhkxx6 = (Llkxx6 & Slkxx6);
assign Slkxx6 = (Zlkxx6 & Gmkxx6);
assign Gmkxx6 = (Nmkxx6 & Umkxx6);
assign Umkxx6 = (~(Phjxx6 & vis_r8_o[3]));
assign Nmkxx6 = (~(Okjxx6 & vis_r6_o[3]));
assign Zlkxx6 = (Bnkxx6 & Inkxx6);
assign Inkxx6 = (~(Vkjxx6 & vis_r5_o[3]));
assign Bnkxx6 = (~(Qljxx6 & vis_r4_o[3]));
assign Llkxx6 = (Pnkxx6 & Wnkxx6);
assign Wnkxx6 = (Dokxx6 & Kokxx6);
assign Kokxx6 = (~(Xljxx6 & vis_r3_o[3]));
assign Dokxx6 = (~(Nnjxx6 & vis_r0_o[3]));
assign Pnkxx6 = (Rokxx6 & Yokxx6);
assign Yokxx6 = (~(Unjxx6 & vis_r2_o[3]));
assign Rokxx6 = (~(Smjxx6 & vis_r1_o[3]));
assign Xdkxx6 = (Fpkxx6 & Mpkxx6);
assign Mpkxx6 = (~(K1i7z6[3] & Zs4ov6));
assign Fpkxx6 = (Tpkxx6 & Aqkxx6);
assign Aqkxx6 = (~(Xzjxx6 & vis_pc_o[3]));
assign Tpkxx6 = (~(S8jxx6 & Cmm7z6[3]));
assign Wbs7v6 = (~(Hqkxx6 & Oqkxx6));
assign Oqkxx6 = (Vqkxx6 & Crkxx6);
assign Crkxx6 = (~(U9jxx6 & Bgjnv6));
assign Bgjnv6 = (~(Jrkxx6 & Qrkxx6));
assign Qrkxx6 = (Xrkxx6 & Eskxx6);
assign Eskxx6 = (~(Cb77x6 & Kbjxx6));
assign Xrkxx6 = (~(Tw57x6 & Rbjxx6));
assign Jrkxx6 = (Lskxx6 & Sskxx6);
assign Sskxx6 = (~(Ax57x6 & Mcjxx6));
assign Lskxx6 = (~(T977x6 & Tcjxx6));
assign Vqkxx6 = (Zskxx6 & Wgkxx6);
assign Zskxx6 = (Adjxx6 | Jy2jw6);
assign Jy2jw6 = (Gtkxx6 & Ntkxx6);
assign Ntkxx6 = (Utkxx6 & Bukxx6);
assign Bukxx6 = (Iukxx6 & Pukxx6);
assign Pukxx6 = (Wukxx6 & Dvkxx6);
assign Dvkxx6 = (~(X6kxx6 & vis_psp_o[4]));
assign Wukxx6 = (~(E7kxx6 & vis_msp_o[4]));
assign Iukxx6 = (Kvkxx6 & Rvkxx6);
assign Rvkxx6 = (~(Lfjxx6 & Pic7z6[4]));
assign Kvkxx6 = (~(Sfjxx6 & vis_r12_o[4]));
assign Utkxx6 = (Yvkxx6 & Fwkxx6);
assign Fwkxx6 = (Mwkxx6 & Twkxx6);
assign Twkxx6 = (~(Ngjxx6 & vis_r11_o[4]));
assign Mwkxx6 = (~(Ugjxx6 & vis_r10_o[4]));
assign Yvkxx6 = (Axkxx6 & Hxkxx6);
assign Hxkxx6 = (~(Kijxx6 & vis_r7_o[4]));
assign Axkxx6 = (~(Rijxx6 & vis_r9_o[4]));
assign Gtkxx6 = (Oxkxx6 & Vxkxx6);
assign Vxkxx6 = (Cykxx6 & Jykxx6);
assign Jykxx6 = (Qykxx6 & Xykxx6);
assign Xykxx6 = (~(Phjxx6 & vis_r8_o[4]));
assign Qykxx6 = (~(Okjxx6 & vis_r6_o[4]));
assign Cykxx6 = (Ezkxx6 & Lzkxx6);
assign Lzkxx6 = (~(Vkjxx6 & vis_r5_o[4]));
assign Ezkxx6 = (~(Qljxx6 & vis_r4_o[4]));
assign Oxkxx6 = (Szkxx6 & Zzkxx6);
assign Zzkxx6 = (G0lxx6 & N0lxx6);
assign N0lxx6 = (~(Xljxx6 & vis_r3_o[4]));
assign G0lxx6 = (~(Nnjxx6 & vis_r0_o[4]));
assign Szkxx6 = (U0lxx6 & B1lxx6);
assign B1lxx6 = (~(Unjxx6 & vis_r2_o[4]));
assign U0lxx6 = (~(Smjxx6 & vis_r1_o[4]));
assign Hqkxx6 = (I1lxx6 & P1lxx6);
assign P1lxx6 = (~(K1i7z6[4] & Zs4ov6));
assign I1lxx6 = (W1lxx6 & D2lxx6);
assign D2lxx6 = (~(Xzjxx6 & vis_pc_o[4]));
assign W1lxx6 = (~(S8jxx6 & Cmm7z6[4]));
assign Pbs7v6 = (~(K2lxx6 & R2lxx6));
assign R2lxx6 = (Y2lxx6 & F3lxx6);
assign F3lxx6 = (~(U9jxx6 & Lejnv6));
assign Lejnv6 = (~(M3lxx6 & T3lxx6));
assign T3lxx6 = (A4lxx6 & H4lxx6);
assign H4lxx6 = (~(C477x6 & Kbjxx6));
assign A4lxx6 = (~(Qr57x6 & Rbjxx6));
assign M3lxx6 = (O4lxx6 & V4lxx6);
assign V4lxx6 = (~(Xr57x6 & Mcjxx6));
assign O4lxx6 = (~(T277x6 & Tcjxx6));
assign Y2lxx6 = (C5lxx6 & Wgkxx6);
assign C5lxx6 = (Adjxx6 | Hei6x6);
assign Hei6x6 = (J5lxx6 & Q5lxx6);
assign Q5lxx6 = (X5lxx6 & E6lxx6);
assign E6lxx6 = (L6lxx6 & S6lxx6);
assign S6lxx6 = (Z6lxx6 & G7lxx6);
assign G7lxx6 = (~(X6kxx6 & vis_psp_o[5]));
assign Z6lxx6 = (~(E7kxx6 & vis_msp_o[5]));
assign L6lxx6 = (N7lxx6 & U7lxx6);
assign U7lxx6 = (~(Lfjxx6 & Pic7z6[5]));
assign N7lxx6 = (~(Sfjxx6 & vis_r12_o[5]));
assign X5lxx6 = (B8lxx6 & I8lxx6);
assign I8lxx6 = (P8lxx6 & W8lxx6);
assign W8lxx6 = (~(Ngjxx6 & vis_r11_o[5]));
assign P8lxx6 = (~(Ugjxx6 & vis_r10_o[5]));
assign B8lxx6 = (D9lxx6 & K9lxx6);
assign K9lxx6 = (~(Kijxx6 & vis_r7_o[5]));
assign D9lxx6 = (~(Rijxx6 & vis_r9_o[5]));
assign J5lxx6 = (R9lxx6 & Y9lxx6);
assign Y9lxx6 = (Falxx6 & Malxx6);
assign Malxx6 = (Talxx6 & Ablxx6);
assign Ablxx6 = (~(Phjxx6 & vis_r8_o[5]));
assign Talxx6 = (~(Okjxx6 & vis_r6_o[5]));
assign Falxx6 = (Hblxx6 & Oblxx6);
assign Oblxx6 = (~(Vkjxx6 & vis_r5_o[5]));
assign Hblxx6 = (~(Qljxx6 & vis_r4_o[5]));
assign R9lxx6 = (Vblxx6 & Cclxx6);
assign Cclxx6 = (Jclxx6 & Qclxx6);
assign Qclxx6 = (~(Xljxx6 & vis_r3_o[5]));
assign Jclxx6 = (~(Nnjxx6 & vis_r0_o[5]));
assign Vblxx6 = (Xclxx6 & Edlxx6);
assign Edlxx6 = (~(Unjxx6 & vis_r2_o[5]));
assign Xclxx6 = (~(Smjxx6 & vis_r1_o[5]));
assign K2lxx6 = (Ldlxx6 & Sdlxx6);
assign Sdlxx6 = (~(K1i7z6[5] & Zs4ov6));
assign Ldlxx6 = (Zdlxx6 & Gelxx6);
assign Gelxx6 = (~(Xzjxx6 & vis_pc_o[5]));
assign Zdlxx6 = (~(S8jxx6 & Cmm7z6[5]));
assign Ibs7v6 = (~(Nelxx6 & Uelxx6));
assign Uelxx6 = (Bflxx6 & Iflxx6);
assign Iflxx6 = (~(U9jxx6 & Vcjnv6));
assign Vcjnv6 = (~(Pflxx6 & Wflxx6));
assign Wflxx6 = (Dglxx6 & Kglxx6);
assign Kglxx6 = (~(Cx67x6 & Kbjxx6));
assign Dglxx6 = (~(Nm57x6 & Rbjxx6));
assign Pflxx6 = (Rglxx6 & Yglxx6);
assign Yglxx6 = (~(Um57x6 & Mcjxx6));
assign Rglxx6 = (~(Tv67x6 & Tcjxx6));
assign Bflxx6 = (Fhlxx6 & Wgkxx6);
assign Fhlxx6 = (Adjxx6 | F3l6x6);
assign F3l6x6 = (Mhlxx6 & Thlxx6);
assign Thlxx6 = (Ailxx6 & Hilxx6);
assign Hilxx6 = (Oilxx6 & Vilxx6);
assign Vilxx6 = (Cjlxx6 & Jjlxx6);
assign Jjlxx6 = (~(X6kxx6 & vis_psp_o[6]));
assign Cjlxx6 = (~(E7kxx6 & vis_msp_o[6]));
assign Oilxx6 = (Qjlxx6 & Xjlxx6);
assign Xjlxx6 = (~(Lfjxx6 & Pic7z6[6]));
assign Qjlxx6 = (~(Sfjxx6 & vis_r12_o[6]));
assign Ailxx6 = (Eklxx6 & Lklxx6);
assign Lklxx6 = (Sklxx6 & Zklxx6);
assign Zklxx6 = (~(Ngjxx6 & vis_r11_o[6]));
assign Sklxx6 = (~(Ugjxx6 & vis_r10_o[6]));
assign Eklxx6 = (Gllxx6 & Nllxx6);
assign Nllxx6 = (~(Kijxx6 & vis_r7_o[6]));
assign Gllxx6 = (~(Rijxx6 & vis_r9_o[6]));
assign Mhlxx6 = (Ullxx6 & Bmlxx6);
assign Bmlxx6 = (Imlxx6 & Pmlxx6);
assign Pmlxx6 = (Wmlxx6 & Dnlxx6);
assign Dnlxx6 = (~(Phjxx6 & vis_r8_o[6]));
assign Wmlxx6 = (~(Okjxx6 & vis_r6_o[6]));
assign Imlxx6 = (Knlxx6 & Rnlxx6);
assign Rnlxx6 = (~(Vkjxx6 & vis_r5_o[6]));
assign Knlxx6 = (~(Qljxx6 & vis_r4_o[6]));
assign Ullxx6 = (Ynlxx6 & Folxx6);
assign Folxx6 = (Molxx6 & Tolxx6);
assign Tolxx6 = (~(Xljxx6 & vis_r3_o[6]));
assign Molxx6 = (~(Nnjxx6 & vis_r0_o[6]));
assign Ynlxx6 = (Aplxx6 & Hplxx6);
assign Hplxx6 = (~(Unjxx6 & vis_r2_o[6]));
assign Aplxx6 = (~(Smjxx6 & vis_r1_o[6]));
assign Nelxx6 = (Oplxx6 & Vplxx6);
assign Vplxx6 = (~(K1i7z6[6] & Zs4ov6));
assign Oplxx6 = (Cqlxx6 & Jqlxx6);
assign Jqlxx6 = (~(Xzjxx6 & vis_pc_o[6]));
assign Cqlxx6 = (~(S8jxx6 & Cmm7z6[6]));
assign Bbs7v6 = (~(Qqlxx6 & Xqlxx6));
assign Xqlxx6 = (Erlxx6 & Lrlxx6);
assign Lrlxx6 = (~(U9jxx6 & Fbjnv6));
assign Fbjnv6 = (~(Srlxx6 & Zrlxx6));
assign Zrlxx6 = (Gslxx6 & Nslxx6);
assign Nslxx6 = (~(Hp67x6 & Kbjxx6));
assign Kbjxx6 = (~(Uslxx6 & Btlxx6));
assign Btlxx6 = (~(Itlxx6 & Gaa7x6));
assign Uslxx6 = (Ptlxx6 & Wtlxx6);
assign Ptlxx6 = (~(Av77x6 & Dulxx6));
assign Gslxx6 = (~(Dh57x6 & Rbjxx6));
assign Rbjxx6 = (~(Kulxx6 & Rulxx6));
assign Rulxx6 = (~(Itlxx6 & Av77x6));
assign Kulxx6 = (Yulxx6 & Fvlxx6);
assign Yulxx6 = (~(Dca7x6 & Dulxx6));
assign Srlxx6 = (Mvlxx6 & Tvlxx6);
assign Tvlxx6 = (~(Mcjxx6 & Rh57x6));
assign Mcjxx6 = (~(Awlxx6 & Hwlxx6));
assign Hwlxx6 = (~(Itlxx6 & Dca7x6));
assign Awlxx6 = (Owlxx6 & Vwlxx6);
assign Owlxx6 = (~(H287x6 & Dulxx6));
assign Mvlxx6 = (~(Kn67x6 & Tcjxx6));
assign Tcjxx6 = (~(Cxlxx6 & Jxlxx6));
assign Jxlxx6 = (~(Itlxx6 & H287x6));
assign Cxlxx6 = (Qxlxx6 & Xxlxx6);
assign Qxlxx6 = (~(Gaa7x6 & Dulxx6));
assign Dulxx6 = (Xgmov6 | Eylxx6);
assign Erlxx6 = (Lylxx6 & Wgkxx6);
assign Lylxx6 = (Adjxx6 | Brn6x6);
assign Brn6x6 = (Sylxx6 & Zylxx6);
assign Zylxx6 = (Gzlxx6 & Nzlxx6);
assign Nzlxx6 = (Uzlxx6 & B0mxx6);
assign B0mxx6 = (I0mxx6 & P0mxx6);
assign P0mxx6 = (~(X6kxx6 & vis_psp_o[7]));
assign I0mxx6 = (~(E7kxx6 & vis_msp_o[7]));
assign Uzlxx6 = (W0mxx6 & D1mxx6);
assign D1mxx6 = (~(Lfjxx6 & Pic7z6[7]));
assign W0mxx6 = (~(Sfjxx6 & vis_r12_o[7]));
assign Gzlxx6 = (K1mxx6 & R1mxx6);
assign R1mxx6 = (Y1mxx6 & F2mxx6);
assign F2mxx6 = (~(Ngjxx6 & vis_r11_o[7]));
assign Y1mxx6 = (~(Ugjxx6 & vis_r10_o[7]));
assign K1mxx6 = (M2mxx6 & T2mxx6);
assign T2mxx6 = (~(Kijxx6 & vis_r7_o[7]));
assign M2mxx6 = (~(Rijxx6 & vis_r9_o[7]));
assign Sylxx6 = (A3mxx6 & H3mxx6);
assign H3mxx6 = (O3mxx6 & V3mxx6);
assign V3mxx6 = (C4mxx6 & J4mxx6);
assign J4mxx6 = (~(Phjxx6 & vis_r8_o[7]));
assign C4mxx6 = (~(Okjxx6 & vis_r6_o[7]));
assign O3mxx6 = (Q4mxx6 & X4mxx6);
assign X4mxx6 = (~(Vkjxx6 & vis_r5_o[7]));
assign Q4mxx6 = (~(Qljxx6 & vis_r4_o[7]));
assign A3mxx6 = (E5mxx6 & L5mxx6);
assign L5mxx6 = (S5mxx6 & Z5mxx6);
assign Z5mxx6 = (~(Xljxx6 & vis_r3_o[7]));
assign S5mxx6 = (~(Nnjxx6 & vis_r0_o[7]));
assign E5mxx6 = (G6mxx6 & N6mxx6);
assign N6mxx6 = (~(Unjxx6 & vis_r2_o[7]));
assign G6mxx6 = (~(Smjxx6 & vis_r1_o[7]));
assign Qqlxx6 = (U6mxx6 & B7mxx6);
assign B7mxx6 = (~(K1i7z6[7] & Zs4ov6));
assign U6mxx6 = (I7mxx6 & P7mxx6);
assign P7mxx6 = (~(Xzjxx6 & vis_pc_o[7]));
assign I7mxx6 = (~(S8jxx6 & Cmm7z6[7]));
assign Uas7v6 = (~(W7mxx6 & D8mxx6));
assign D8mxx6 = (K8mxx6 & R8mxx6);
assign R8mxx6 = (~(U9jxx6 & P9jnv6));
assign P9jnv6 = (~(Y8mxx6 & F9mxx6));
assign F9mxx6 = (M9mxx6 & T9mxx6);
assign T9mxx6 = (~(Aamxx6 & Td9ov6));
assign M9mxx6 = (Hamxx6 & Oamxx6);
assign Oamxx6 = (~(Vamxx6 & Jf9ov6));
assign Hamxx6 = (~(Cbmxx6 & Ve9ov6));
assign Y8mxx6 = (Jbmxx6 & Qbmxx6);
assign Qbmxx6 = (~(Xbmxx6 & Fd9ov6));
assign K8mxx6 = (Ecmxx6 & Wgkxx6);
assign Ecmxx6 = (Adjxx6 | Mo3jw6);
assign Mo3jw6 = (Lcmxx6 & Scmxx6);
assign Scmxx6 = (Zcmxx6 & Gdmxx6);
assign Gdmxx6 = (Ndmxx6 & Udmxx6);
assign Udmxx6 = (Bemxx6 & Iemxx6);
assign Iemxx6 = (~(X6kxx6 & vis_psp_o[8]));
assign Bemxx6 = (~(E7kxx6 & vis_msp_o[8]));
assign Ndmxx6 = (Pemxx6 & Wemxx6);
assign Wemxx6 = (~(Lfjxx6 & Pic7z6[8]));
assign Pemxx6 = (~(Sfjxx6 & vis_r12_o[8]));
assign Zcmxx6 = (Dfmxx6 & Kfmxx6);
assign Kfmxx6 = (Rfmxx6 & Yfmxx6);
assign Yfmxx6 = (~(Ngjxx6 & vis_r11_o[8]));
assign Rfmxx6 = (~(Ugjxx6 & vis_r10_o[8]));
assign Dfmxx6 = (Fgmxx6 & Mgmxx6);
assign Mgmxx6 = (~(Kijxx6 & vis_r7_o[8]));
assign Fgmxx6 = (~(Rijxx6 & vis_r9_o[8]));
assign Lcmxx6 = (Tgmxx6 & Ahmxx6);
assign Ahmxx6 = (Hhmxx6 & Ohmxx6);
assign Ohmxx6 = (Vhmxx6 & Cimxx6);
assign Cimxx6 = (~(Phjxx6 & vis_r8_o[8]));
assign Vhmxx6 = (~(Okjxx6 & vis_r6_o[8]));
assign Hhmxx6 = (Jimxx6 & Qimxx6);
assign Qimxx6 = (~(Vkjxx6 & vis_r5_o[8]));
assign Jimxx6 = (~(Qljxx6 & vis_r4_o[8]));
assign Tgmxx6 = (Ximxx6 & Ejmxx6);
assign Ejmxx6 = (Ljmxx6 & Sjmxx6);
assign Sjmxx6 = (~(Xljxx6 & vis_r3_o[8]));
assign Ljmxx6 = (~(Nnjxx6 & vis_r0_o[8]));
assign Ximxx6 = (Zjmxx6 & Gkmxx6);
assign Gkmxx6 = (~(Unjxx6 & vis_r2_o[8]));
assign Zjmxx6 = (~(Smjxx6 & vis_r1_o[8]));
assign W7mxx6 = (Nkmxx6 & Ukmxx6);
assign Ukmxx6 = (~(K1i7z6[8] & Zs4ov6));
assign Nkmxx6 = (Blmxx6 & Ilmxx6);
assign Ilmxx6 = (~(Xzjxx6 & vis_pc_o[8]));
assign Blmxx6 = (~(S8jxx6 & Cmm7z6[8]));
assign Nas7v6 = (~(Plmxx6 & Wlmxx6));
assign Wlmxx6 = (Dmmxx6 & Kmmxx6);
assign Kmmxx6 = (~(Xzjxx6 & vis_pc_o[9]));
assign Dmmxx6 = (Rmmxx6 & Ymmxx6);
assign Ymmxx6 = (~(U9jxx6 & L7jnv6));
assign L7jnv6 = (~(Fnmxx6 & Mnmxx6));
assign Mnmxx6 = (Tnmxx6 & Aomxx6);
assign Aomxx6 = (~(Aamxx6 & Ex77x6));
assign Tnmxx6 = (Homxx6 & Oomxx6);
assign Oomxx6 = (~(Vamxx6 & Ab67x6));
assign Homxx6 = (~(Cbmxx6 & Ob67x6));
assign Fnmxx6 = (Jbmxx6 & Vomxx6);
assign Vomxx6 = (~(Xbmxx6 & Vv77x6));
assign Rmmxx6 = (Adjxx6 | L79jw6);
assign L79jw6 = (Cpmxx6 & Jpmxx6);
assign Jpmxx6 = (Qpmxx6 & Xpmxx6);
assign Xpmxx6 = (Eqmxx6 & Lqmxx6);
assign Lqmxx6 = (Sqmxx6 & Zqmxx6);
assign Zqmxx6 = (~(X6kxx6 & vis_psp_o[9]));
assign Sqmxx6 = (~(E7kxx6 & vis_msp_o[9]));
assign Eqmxx6 = (Grmxx6 & Nrmxx6);
assign Nrmxx6 = (~(Lfjxx6 & Pic7z6[9]));
assign Grmxx6 = (~(Sfjxx6 & vis_r12_o[9]));
assign Qpmxx6 = (Urmxx6 & Bsmxx6);
assign Bsmxx6 = (Ismxx6 & Psmxx6);
assign Psmxx6 = (~(Ngjxx6 & vis_r11_o[9]));
assign Ismxx6 = (~(Ugjxx6 & vis_r10_o[9]));
assign Urmxx6 = (Wsmxx6 & Dtmxx6);
assign Dtmxx6 = (~(Kijxx6 & vis_r7_o[9]));
assign Wsmxx6 = (~(Rijxx6 & vis_r9_o[9]));
assign Cpmxx6 = (Ktmxx6 & Rtmxx6);
assign Rtmxx6 = (Ytmxx6 & Fumxx6);
assign Fumxx6 = (Mumxx6 & Tumxx6);
assign Tumxx6 = (~(Phjxx6 & vis_r8_o[9]));
assign Mumxx6 = (~(Okjxx6 & vis_r6_o[9]));
assign Ytmxx6 = (Avmxx6 & Hvmxx6);
assign Hvmxx6 = (~(Vkjxx6 & vis_r5_o[9]));
assign Avmxx6 = (~(Qljxx6 & vis_r4_o[9]));
assign Ktmxx6 = (Ovmxx6 & Vvmxx6);
assign Vvmxx6 = (Cwmxx6 & Jwmxx6);
assign Jwmxx6 = (~(Xljxx6 & vis_r3_o[9]));
assign Cwmxx6 = (~(Nnjxx6 & vis_r0_o[9]));
assign Ovmxx6 = (Qwmxx6 & Xwmxx6);
assign Xwmxx6 = (~(Unjxx6 & vis_r2_o[9]));
assign Qwmxx6 = (~(Smjxx6 & vis_r1_o[9]));
assign Plmxx6 = (Exmxx6 & Lxmxx6);
assign Lxmxx6 = (~(S8jxx6 & Cmm7z6[9]));
assign Exmxx6 = (~(K1i7z6[9] & Zs4ov6));
assign Gas7v6 = (~(Sxmxx6 & Zxmxx6));
assign Zxmxx6 = (Gymxx6 & Nymxx6);
assign Nymxx6 = (~(U9jxx6 & Glknv6));
assign Glknv6 = (~(Uymxx6 & Bzmxx6));
assign Bzmxx6 = (Izmxx6 & Pzmxx6);
assign Pzmxx6 = (~(Aamxx6 & Icfov6));
assign Izmxx6 = (Wzmxx6 & D0nxx6);
assign D0nxx6 = (~(Kdfov6 & Vamxx6));
assign Wzmxx6 = (~(Ddfov6 & Cbmxx6));
assign Uymxx6 = (Jbmxx6 & K0nxx6);
assign K0nxx6 = (~(Xbmxx6 & Bcfov6));
assign Gymxx6 = (R0nxx6 & Wgkxx6);
assign R0nxx6 = (Adjxx6 | Sc4jw6);
assign Sc4jw6 = (Y0nxx6 & F1nxx6);
assign F1nxx6 = (M1nxx6 & T1nxx6);
assign T1nxx6 = (A2nxx6 & H2nxx6);
assign H2nxx6 = (O2nxx6 & V2nxx6);
assign V2nxx6 = (~(X6kxx6 & vis_psp_o[10]));
assign O2nxx6 = (~(E7kxx6 & vis_msp_o[10]));
assign A2nxx6 = (C3nxx6 & J3nxx6);
assign J3nxx6 = (~(Lfjxx6 & Pic7z6[10]));
assign C3nxx6 = (~(Sfjxx6 & vis_r12_o[10]));
assign M1nxx6 = (Q3nxx6 & X3nxx6);
assign X3nxx6 = (E4nxx6 & L4nxx6);
assign L4nxx6 = (~(Ngjxx6 & vis_r11_o[10]));
assign E4nxx6 = (~(Ugjxx6 & vis_r10_o[10]));
assign Q3nxx6 = (S4nxx6 & Z4nxx6);
assign Z4nxx6 = (~(Kijxx6 & vis_r7_o[10]));
assign S4nxx6 = (~(Rijxx6 & vis_r9_o[10]));
assign Y0nxx6 = (G5nxx6 & N5nxx6);
assign N5nxx6 = (U5nxx6 & B6nxx6);
assign B6nxx6 = (I6nxx6 & P6nxx6);
assign P6nxx6 = (~(Phjxx6 & vis_r8_o[10]));
assign I6nxx6 = (~(Okjxx6 & vis_r6_o[10]));
assign U5nxx6 = (W6nxx6 & D7nxx6);
assign D7nxx6 = (~(Vkjxx6 & vis_r5_o[10]));
assign W6nxx6 = (~(Qljxx6 & vis_r4_o[10]));
assign G5nxx6 = (K7nxx6 & R7nxx6);
assign R7nxx6 = (Y7nxx6 & F8nxx6);
assign F8nxx6 = (~(Xljxx6 & vis_r3_o[10]));
assign Y7nxx6 = (~(Nnjxx6 & vis_r0_o[10]));
assign K7nxx6 = (M8nxx6 & T8nxx6);
assign T8nxx6 = (~(Unjxx6 & vis_r2_o[10]));
assign M8nxx6 = (~(Smjxx6 & vis_r1_o[10]));
assign Sxmxx6 = (A9nxx6 & H9nxx6);
assign H9nxx6 = (~(K1i7z6[10] & Zs4ov6));
assign A9nxx6 = (O9nxx6 & V9nxx6);
assign V9nxx6 = (~(Xzjxx6 & vis_pc_o[10]));
assign O9nxx6 = (~(S8jxx6 & Cmm7z6[10]));
assign Z9s7v6 = (~(Canxx6 & Janxx6));
assign Janxx6 = (Qanxx6 & Xanxx6);
assign Xanxx6 = (~(U9jxx6 & Jjknv6));
assign Jjknv6 = (~(Ebnxx6 & Lbnxx6));
assign Lbnxx6 = (Sbnxx6 & Zbnxx6);
assign Zbnxx6 = (~(Mmlov6 & Aamxx6));
assign Sbnxx6 = (Gcnxx6 & Ncnxx6);
assign Ncnxx6 = (~(Onlov6 & Vamxx6));
assign Gcnxx6 = (~(Hnlov6 & Cbmxx6));
assign Ebnxx6 = (Jbmxx6 & Ucnxx6);
assign Ucnxx6 = (~(Fmlov6 & Xbmxx6));
assign Qanxx6 = (Bdnxx6 & Wgkxx6);
assign Bdnxx6 = (Adjxx6 | Lyajw6);
assign Lyajw6 = (Idnxx6 & Pdnxx6);
assign Pdnxx6 = (Wdnxx6 & Denxx6);
assign Denxx6 = (Kenxx6 & Renxx6);
assign Renxx6 = (Yenxx6 & Ffnxx6);
assign Ffnxx6 = (~(X6kxx6 & vis_psp_o[11]));
assign Yenxx6 = (~(E7kxx6 & vis_msp_o[11]));
assign Kenxx6 = (Mfnxx6 & Tfnxx6);
assign Tfnxx6 = (~(Lfjxx6 & Pic7z6[11]));
assign Mfnxx6 = (~(Sfjxx6 & vis_r12_o[11]));
assign Wdnxx6 = (Agnxx6 & Hgnxx6);
assign Hgnxx6 = (Ognxx6 & Vgnxx6);
assign Vgnxx6 = (~(Ngjxx6 & vis_r11_o[11]));
assign Ognxx6 = (~(Ugjxx6 & vis_r10_o[11]));
assign Agnxx6 = (Chnxx6 & Jhnxx6);
assign Jhnxx6 = (~(Kijxx6 & vis_r7_o[11]));
assign Chnxx6 = (~(Rijxx6 & vis_r9_o[11]));
assign Idnxx6 = (Qhnxx6 & Xhnxx6);
assign Xhnxx6 = (Einxx6 & Linxx6);
assign Linxx6 = (Sinxx6 & Zinxx6);
assign Zinxx6 = (~(Phjxx6 & vis_r8_o[11]));
assign Sinxx6 = (~(Okjxx6 & vis_r6_o[11]));
assign Einxx6 = (Gjnxx6 & Njnxx6);
assign Njnxx6 = (~(Vkjxx6 & vis_r5_o[11]));
assign Gjnxx6 = (~(Qljxx6 & vis_r4_o[11]));
assign Qhnxx6 = (Ujnxx6 & Bknxx6);
assign Bknxx6 = (Iknxx6 & Pknxx6);
assign Pknxx6 = (~(Xljxx6 & vis_r3_o[11]));
assign Iknxx6 = (~(Nnjxx6 & vis_r0_o[11]));
assign Ujnxx6 = (Wknxx6 & Dlnxx6);
assign Dlnxx6 = (~(Unjxx6 & vis_r2_o[11]));
assign Wknxx6 = (~(Smjxx6 & vis_r1_o[11]));
assign Canxx6 = (Klnxx6 & Rlnxx6);
assign Rlnxx6 = (~(K1i7z6[11] & Zs4ov6));
assign Klnxx6 = (Ylnxx6 & Fmnxx6);
assign Fmnxx6 = (~(Xzjxx6 & vis_pc_o[11]));
assign Ylnxx6 = (~(S8jxx6 & Cmm7z6[11]));
assign S9s7v6 = (~(Mmnxx6 & Tmnxx6));
assign Tmnxx6 = (Annxx6 & Hnnxx6);
assign Hnnxx6 = (~(Xzjxx6 & vis_pc_o[12]));
assign Annxx6 = (Onnxx6 & Vnnxx6);
assign Vnnxx6 = (~(U9jxx6 & Thknv6));
assign Thknv6 = (~(Conxx6 & Jonxx6));
assign Jonxx6 = (Qonxx6 & Xonxx6);
assign Xonxx6 = (~(Cb77x6 & Aamxx6));
assign Qonxx6 = (Epnxx6 & Lpnxx6);
assign Lpnxx6 = (~(Tw57x6 & Vamxx6));
assign Epnxx6 = (~(Ax57x6 & Cbmxx6));
assign Conxx6 = (Jbmxx6 & Spnxx6);
assign Spnxx6 = (~(T977x6 & Xbmxx6));
assign Onnxx6 = (Adjxx6 | Tmg6x6);
assign Tmg6x6 = (Zpnxx6 & Gqnxx6);
assign Gqnxx6 = (Nqnxx6 & Uqnxx6);
assign Uqnxx6 = (Brnxx6 & Irnxx6);
assign Irnxx6 = (Prnxx6 & Wrnxx6);
assign Wrnxx6 = (~(X6kxx6 & vis_psp_o[12]));
assign Prnxx6 = (~(E7kxx6 & vis_msp_o[12]));
assign Brnxx6 = (Dsnxx6 & Ksnxx6);
assign Ksnxx6 = (~(Lfjxx6 & Pic7z6[12]));
assign Dsnxx6 = (~(Sfjxx6 & vis_r12_o[12]));
assign Nqnxx6 = (Rsnxx6 & Ysnxx6);
assign Ysnxx6 = (Ftnxx6 & Mtnxx6);
assign Mtnxx6 = (~(Ngjxx6 & vis_r11_o[12]));
assign Ftnxx6 = (~(Ugjxx6 & vis_r10_o[12]));
assign Rsnxx6 = (Ttnxx6 & Aunxx6);
assign Aunxx6 = (~(Kijxx6 & vis_r7_o[12]));
assign Ttnxx6 = (~(Rijxx6 & vis_r9_o[12]));
assign Zpnxx6 = (Hunxx6 & Ounxx6);
assign Ounxx6 = (Vunxx6 & Cvnxx6);
assign Cvnxx6 = (Jvnxx6 & Qvnxx6);
assign Qvnxx6 = (~(Phjxx6 & vis_r8_o[12]));
assign Jvnxx6 = (~(Okjxx6 & vis_r6_o[12]));
assign Vunxx6 = (Xvnxx6 & Ewnxx6);
assign Ewnxx6 = (~(Vkjxx6 & vis_r5_o[12]));
assign Xvnxx6 = (~(Qljxx6 & vis_r4_o[12]));
assign Hunxx6 = (Lwnxx6 & Swnxx6);
assign Swnxx6 = (Zwnxx6 & Gxnxx6);
assign Gxnxx6 = (~(Xljxx6 & vis_r3_o[12]));
assign Zwnxx6 = (~(Nnjxx6 & vis_r0_o[12]));
assign Lwnxx6 = (Nxnxx6 & Uxnxx6);
assign Uxnxx6 = (~(Unjxx6 & vis_r2_o[12]));
assign Nxnxx6 = (~(Smjxx6 & vis_r1_o[12]));
assign Mmnxx6 = (Bynxx6 & Iynxx6);
assign Iynxx6 = (~(S8jxx6 & Cmm7z6[12]));
assign Bynxx6 = (~(K1i7z6[12] & Zs4ov6));
assign L9s7v6 = (~(Pynxx6 & Wynxx6));
assign Wynxx6 = (Dznxx6 & Kznxx6);
assign Kznxx6 = (~(U9jxx6 & Dgknv6));
assign Dgknv6 = (~(Rznxx6 & Yznxx6));
assign Yznxx6 = (F0oxx6 & M0oxx6);
assign M0oxx6 = (~(C477x6 & Aamxx6));
assign F0oxx6 = (T0oxx6 & A1oxx6);
assign A1oxx6 = (~(Qr57x6 & Vamxx6));
assign T0oxx6 = (~(Xr57x6 & Cbmxx6));
assign Rznxx6 = (Jbmxx6 & H1oxx6);
assign H1oxx6 = (~(T277x6 & Xbmxx6));
assign Dznxx6 = (O1oxx6 & Wgkxx6);
assign O1oxx6 = (Adjxx6 | Z7k6x6);
assign Z7k6x6 = (V1oxx6 & C2oxx6);
assign C2oxx6 = (J2oxx6 & Q2oxx6);
assign Q2oxx6 = (X2oxx6 & E3oxx6);
assign E3oxx6 = (L3oxx6 & S3oxx6);
assign S3oxx6 = (~(X6kxx6 & vis_psp_o[13]));
assign L3oxx6 = (~(E7kxx6 & vis_msp_o[13]));
assign X2oxx6 = (Z3oxx6 & G4oxx6);
assign G4oxx6 = (~(Lfjxx6 & Pic7z6[13]));
assign Z3oxx6 = (~(Sfjxx6 & vis_r12_o[13]));
assign J2oxx6 = (N4oxx6 & U4oxx6);
assign U4oxx6 = (B5oxx6 & I5oxx6);
assign I5oxx6 = (~(Ngjxx6 & vis_r11_o[13]));
assign B5oxx6 = (~(Ugjxx6 & vis_r10_o[13]));
assign N4oxx6 = (P5oxx6 & W5oxx6);
assign W5oxx6 = (~(Kijxx6 & vis_r7_o[13]));
assign P5oxx6 = (~(Rijxx6 & vis_r9_o[13]));
assign V1oxx6 = (D6oxx6 & K6oxx6);
assign K6oxx6 = (R6oxx6 & Y6oxx6);
assign Y6oxx6 = (F7oxx6 & M7oxx6);
assign M7oxx6 = (~(Phjxx6 & vis_r8_o[13]));
assign F7oxx6 = (~(Okjxx6 & vis_r6_o[13]));
assign R6oxx6 = (T7oxx6 & A8oxx6);
assign A8oxx6 = (~(Vkjxx6 & vis_r5_o[13]));
assign T7oxx6 = (~(Qljxx6 & vis_r4_o[13]));
assign D6oxx6 = (H8oxx6 & O8oxx6);
assign O8oxx6 = (V8oxx6 & C9oxx6);
assign C9oxx6 = (~(Xljxx6 & vis_r3_o[13]));
assign V8oxx6 = (~(Nnjxx6 & vis_r0_o[13]));
assign H8oxx6 = (J9oxx6 & Q9oxx6);
assign Q9oxx6 = (~(Unjxx6 & vis_r2_o[13]));
assign J9oxx6 = (~(Smjxx6 & vis_r1_o[13]));
assign Pynxx6 = (X9oxx6 & Eaoxx6);
assign Eaoxx6 = (~(K1i7z6[13] & Zs4ov6));
assign X9oxx6 = (Laoxx6 & Saoxx6);
assign Saoxx6 = (~(Xzjxx6 & vis_pc_o[13]));
assign Laoxx6 = (~(S8jxx6 & Cmm7z6[13]));
assign E9s7v6 = (~(Zaoxx6 & Gboxx6));
assign Gboxx6 = (Nboxx6 & Uboxx6);
assign Uboxx6 = (~(U9jxx6 & Neknv6));
assign Neknv6 = (~(Bcoxx6 & Icoxx6));
assign Icoxx6 = (Pcoxx6 & Wcoxx6);
assign Wcoxx6 = (~(Cx67x6 & Aamxx6));
assign Pcoxx6 = (Ddoxx6 & Kdoxx6);
assign Kdoxx6 = (~(Nm57x6 & Vamxx6));
assign Ddoxx6 = (~(Um57x6 & Cbmxx6));
assign Bcoxx6 = (Jbmxx6 & Rdoxx6);
assign Rdoxx6 = (~(Tv67x6 & Xbmxx6));
assign Nboxx6 = (Ydoxx6 & Wgkxx6);
assign Ydoxx6 = (Adjxx6 | Vvm6x6);
assign Vvm6x6 = (Feoxx6 & Meoxx6);
assign Meoxx6 = (Teoxx6 & Afoxx6);
assign Afoxx6 = (Hfoxx6 & Ofoxx6);
assign Ofoxx6 = (Vfoxx6 & Cgoxx6);
assign Cgoxx6 = (~(X6kxx6 & vis_psp_o[14]));
assign Vfoxx6 = (~(E7kxx6 & vis_msp_o[14]));
assign Hfoxx6 = (Jgoxx6 & Qgoxx6);
assign Qgoxx6 = (~(Lfjxx6 & Pic7z6[14]));
assign Jgoxx6 = (~(Sfjxx6 & vis_r12_o[14]));
assign Teoxx6 = (Xgoxx6 & Ehoxx6);
assign Ehoxx6 = (Lhoxx6 & Shoxx6);
assign Shoxx6 = (~(Ngjxx6 & vis_r11_o[14]));
assign Lhoxx6 = (~(Ugjxx6 & vis_r10_o[14]));
assign Xgoxx6 = (Zhoxx6 & Gioxx6);
assign Gioxx6 = (~(Kijxx6 & vis_r7_o[14]));
assign Zhoxx6 = (~(Rijxx6 & vis_r9_o[14]));
assign Feoxx6 = (Nioxx6 & Uioxx6);
assign Uioxx6 = (Bjoxx6 & Ijoxx6);
assign Ijoxx6 = (Pjoxx6 & Wjoxx6);
assign Wjoxx6 = (~(Phjxx6 & vis_r8_o[14]));
assign Pjoxx6 = (~(Okjxx6 & vis_r6_o[14]));
assign Bjoxx6 = (Dkoxx6 & Kkoxx6);
assign Kkoxx6 = (~(Vkjxx6 & vis_r5_o[14]));
assign Dkoxx6 = (~(Qljxx6 & vis_r4_o[14]));
assign Nioxx6 = (Rkoxx6 & Ykoxx6);
assign Ykoxx6 = (Floxx6 & Mloxx6);
assign Mloxx6 = (~(Xljxx6 & vis_r3_o[14]));
assign Floxx6 = (~(Nnjxx6 & vis_r0_o[14]));
assign Rkoxx6 = (Tloxx6 & Amoxx6);
assign Amoxx6 = (~(Unjxx6 & vis_r2_o[14]));
assign Tloxx6 = (~(Smjxx6 & vis_r1_o[14]));
assign Zaoxx6 = (Hmoxx6 & Omoxx6);
assign Omoxx6 = (~(K1i7z6[14] & Zs4ov6));
assign Hmoxx6 = (Vmoxx6 & Cnoxx6);
assign Cnoxx6 = (~(Xzjxx6 & vis_pc_o[14]));
assign Vmoxx6 = (~(S8jxx6 & Cmm7z6[14]));
assign X8s7v6 = (~(Jnoxx6 & Qnoxx6));
assign Qnoxx6 = (Xnoxx6 & Eooxx6);
assign Eooxx6 = (~(U9jxx6 & Xcknv6));
assign Xcknv6 = (~(Looxx6 & Sooxx6));
assign Sooxx6 = (Zooxx6 & Gpoxx6);
assign Gpoxx6 = (~(Aamxx6 & Hp67x6));
assign Aamxx6 = (~(Npoxx6 & Upoxx6));
assign Upoxx6 = (~(Yc9ov6 & Bqoxx6));
assign Zooxx6 = (Iqoxx6 & Pqoxx6);
assign Pqoxx6 = (~(Vamxx6 & Dh57x6));
assign Vamxx6 = (~(Wqoxx6 & Droxx6));
assign Droxx6 = (~(Md9ov6 & Bqoxx6));
assign Iqoxx6 = (~(Cbmxx6 & Rh57x6));
assign Cbmxx6 = (~(Kroxx6 & Rroxx6));
assign Rroxx6 = (~(Cf9ov6 & Bqoxx6));
assign Looxx6 = (Jbmxx6 & Yroxx6);
assign Yroxx6 = (~(Xbmxx6 & Kn67x6));
assign Xbmxx6 = (~(Fsoxx6 & Msoxx6));
assign Msoxx6 = (~(Oe9ov6 & Bqoxx6));
assign Xnoxx6 = (Tsoxx6 & Wgkxx6);
assign Tsoxx6 = (Adjxx6 | C35jw6);
assign C35jw6 = (Atoxx6 & Htoxx6);
assign Htoxx6 = (Otoxx6 & Vtoxx6);
assign Vtoxx6 = (Cuoxx6 & Juoxx6);
assign Juoxx6 = (Quoxx6 & Xuoxx6);
assign Xuoxx6 = (~(X6kxx6 & vis_psp_o[15]));
assign Quoxx6 = (~(E7kxx6 & vis_msp_o[15]));
assign Cuoxx6 = (Evoxx6 & Lvoxx6);
assign Lvoxx6 = (~(Lfjxx6 & Pic7z6[15]));
assign Evoxx6 = (~(Sfjxx6 & vis_r12_o[15]));
assign Otoxx6 = (Svoxx6 & Zvoxx6);
assign Zvoxx6 = (Gwoxx6 & Nwoxx6);
assign Nwoxx6 = (~(Ngjxx6 & vis_r11_o[15]));
assign Gwoxx6 = (~(Ugjxx6 & vis_r10_o[15]));
assign Svoxx6 = (Uwoxx6 & Bxoxx6);
assign Bxoxx6 = (~(Kijxx6 & vis_r7_o[15]));
assign Uwoxx6 = (~(Rijxx6 & vis_r9_o[15]));
assign Atoxx6 = (Ixoxx6 & Pxoxx6);
assign Pxoxx6 = (Wxoxx6 & Dyoxx6);
assign Dyoxx6 = (Kyoxx6 & Ryoxx6);
assign Ryoxx6 = (~(Phjxx6 & vis_r8_o[15]));
assign Kyoxx6 = (~(Okjxx6 & vis_r6_o[15]));
assign Wxoxx6 = (Yyoxx6 & Fzoxx6);
assign Fzoxx6 = (~(Vkjxx6 & vis_r5_o[15]));
assign Yyoxx6 = (~(Qljxx6 & vis_r4_o[15]));
assign Ixoxx6 = (Mzoxx6 & Tzoxx6);
assign Tzoxx6 = (A0pxx6 & H0pxx6);
assign H0pxx6 = (~(Xljxx6 & vis_r3_o[15]));
assign A0pxx6 = (~(Nnjxx6 & vis_r0_o[15]));
assign Mzoxx6 = (O0pxx6 & V0pxx6);
assign V0pxx6 = (~(Unjxx6 & vis_r2_o[15]));
assign O0pxx6 = (~(Smjxx6 & vis_r1_o[15]));
assign Jnoxx6 = (C1pxx6 & J1pxx6);
assign J1pxx6 = (~(K1i7z6[15] & Zs4ov6));
assign C1pxx6 = (Q1pxx6 & X1pxx6);
assign X1pxx6 = (~(Xzjxx6 & vis_pc_o[15]));
assign Q1pxx6 = (~(S8jxx6 & Cmm7z6[15]));
assign Q8s7v6 = (~(E2pxx6 & L2pxx6));
assign L2pxx6 = (S2pxx6 & Z2pxx6);
assign Z2pxx6 = (~(Xzjxx6 & vis_pc_o[16]));
assign S2pxx6 = (G3pxx6 & N3pxx6);
assign N3pxx6 = (~(U9jxx6 & Hbknv6));
assign Hbknv6 = (~(U3pxx6 & B4pxx6));
assign B4pxx6 = (I4pxx6 & P4pxx6);
assign P4pxx6 = (Vwlxx6 | W4pxx6);
assign I4pxx6 = (D5pxx6 & K5pxx6);
assign K5pxx6 = (Xxlxx6 | Z487x6);
assign D5pxx6 = (Wtlxx6 | G587x6);
assign U3pxx6 = (R5pxx6 & Y5pxx6);
assign Y5pxx6 = (Fvlxx6 | F6pxx6);
assign G3pxx6 = (Adjxx6 | Kb8jw6);
assign Kb8jw6 = (M6pxx6 & T6pxx6);
assign T6pxx6 = (A7pxx6 & H7pxx6);
assign H7pxx6 = (O7pxx6 & V7pxx6);
assign V7pxx6 = (C8pxx6 & J8pxx6);
assign J8pxx6 = (~(X6kxx6 & vis_psp_o[16]));
assign C8pxx6 = (~(E7kxx6 & vis_msp_o[16]));
assign O7pxx6 = (Q8pxx6 & X8pxx6);
assign X8pxx6 = (~(Lfjxx6 & Pic7z6[16]));
assign Q8pxx6 = (~(Sfjxx6 & vis_r12_o[16]));
assign A7pxx6 = (E9pxx6 & L9pxx6);
assign L9pxx6 = (S9pxx6 & Z9pxx6);
assign Z9pxx6 = (~(Ngjxx6 & vis_r11_o[16]));
assign S9pxx6 = (~(Ugjxx6 & vis_r10_o[16]));
assign E9pxx6 = (Gapxx6 & Napxx6);
assign Napxx6 = (~(Kijxx6 & vis_r7_o[16]));
assign Gapxx6 = (~(Rijxx6 & vis_r9_o[16]));
assign M6pxx6 = (Uapxx6 & Bbpxx6);
assign Bbpxx6 = (Ibpxx6 & Pbpxx6);
assign Pbpxx6 = (Wbpxx6 & Dcpxx6);
assign Dcpxx6 = (~(Phjxx6 & vis_r8_o[16]));
assign Wbpxx6 = (~(Okjxx6 & vis_r6_o[16]));
assign Ibpxx6 = (Kcpxx6 & Rcpxx6);
assign Rcpxx6 = (~(Vkjxx6 & vis_r5_o[16]));
assign Kcpxx6 = (~(Qljxx6 & vis_r4_o[16]));
assign Uapxx6 = (Ycpxx6 & Fdpxx6);
assign Fdpxx6 = (Mdpxx6 & Tdpxx6);
assign Tdpxx6 = (~(Xljxx6 & vis_r3_o[16]));
assign Mdpxx6 = (~(Nnjxx6 & vis_r0_o[16]));
assign Ycpxx6 = (Aepxx6 & Hepxx6);
assign Hepxx6 = (~(Unjxx6 & vis_r2_o[16]));
assign Aepxx6 = (~(Smjxx6 & vis_r1_o[16]));
assign E2pxx6 = (Oepxx6 & Vepxx6);
assign Vepxx6 = (~(S8jxx6 & Cmm7z6[16]));
assign Oepxx6 = (~(K1i7z6[16] & Zs4ov6));
assign J8s7v6 = (~(Cfpxx6 & Jfpxx6));
assign Jfpxx6 = (Qfpxx6 & Xfpxx6);
assign Xfpxx6 = (~(Xzjxx6 & vis_pc_o[17]));
assign Qfpxx6 = (Egpxx6 & Lgpxx6);
assign Lgpxx6 = (~(U9jxx6 & R9knv6));
assign R9knv6 = (~(Sgpxx6 & Zgpxx6));
assign Zgpxx6 = (Ghpxx6 & Nhpxx6);
assign Nhpxx6 = (Vwlxx6 | Cu97x6);
assign Ghpxx6 = (Uhpxx6 & Bipxx6);
assign Bipxx6 = (Xxlxx6 | Iipxx6);
assign Uhpxx6 = (Wtlxx6 | Pipxx6);
assign Sgpxx6 = (R5pxx6 & Wipxx6);
assign Wipxx6 = (Fvlxx6 | Ju97x6);
assign Egpxx6 = (Adjxx6 | R2ajw6);
assign R2ajw6 = (Djpxx6 & Kjpxx6);
assign Kjpxx6 = (Rjpxx6 & Yjpxx6);
assign Yjpxx6 = (Fkpxx6 & Mkpxx6);
assign Mkpxx6 = (Tkpxx6 & Alpxx6);
assign Alpxx6 = (~(X6kxx6 & vis_psp_o[17]));
assign Tkpxx6 = (~(E7kxx6 & vis_msp_o[17]));
assign Fkpxx6 = (Hlpxx6 & Olpxx6);
assign Olpxx6 = (~(Lfjxx6 & Pic7z6[17]));
assign Hlpxx6 = (~(Sfjxx6 & vis_r12_o[17]));
assign Rjpxx6 = (Vlpxx6 & Cmpxx6);
assign Cmpxx6 = (Jmpxx6 & Qmpxx6);
assign Qmpxx6 = (~(Ngjxx6 & vis_r11_o[17]));
assign Jmpxx6 = (~(Ugjxx6 & vis_r10_o[17]));
assign Vlpxx6 = (Xmpxx6 & Enpxx6);
assign Enpxx6 = (~(Kijxx6 & vis_r7_o[17]));
assign Xmpxx6 = (~(Rijxx6 & vis_r9_o[17]));
assign Djpxx6 = (Lnpxx6 & Snpxx6);
assign Snpxx6 = (Znpxx6 & Gopxx6);
assign Gopxx6 = (Nopxx6 & Uopxx6);
assign Uopxx6 = (~(Phjxx6 & vis_r8_o[17]));
assign Nopxx6 = (~(Okjxx6 & vis_r6_o[17]));
assign Znpxx6 = (Bppxx6 & Ippxx6);
assign Ippxx6 = (~(Vkjxx6 & vis_r5_o[17]));
assign Bppxx6 = (~(Qljxx6 & vis_r4_o[17]));
assign Lnpxx6 = (Pppxx6 & Wppxx6);
assign Wppxx6 = (Dqpxx6 & Kqpxx6);
assign Kqpxx6 = (~(Xljxx6 & vis_r3_o[17]));
assign Dqpxx6 = (~(Nnjxx6 & vis_r0_o[17]));
assign Pppxx6 = (Rqpxx6 & Yqpxx6);
assign Yqpxx6 = (~(Unjxx6 & vis_r2_o[17]));
assign Rqpxx6 = (~(Smjxx6 & vis_r1_o[17]));
assign Cfpxx6 = (Frpxx6 & Mrpxx6);
assign Mrpxx6 = (~(S8jxx6 & Cmm7z6[17]));
assign Frpxx6 = (~(K1i7z6[17] & Zs4ov6));
assign C8s7v6 = (~(Trpxx6 & Aspxx6));
assign Aspxx6 = (Hspxx6 & Ospxx6);
assign Ospxx6 = (~(Xzjxx6 & vis_pc_o[18]));
assign Hspxx6 = (Vspxx6 & Ctpxx6);
assign Ctpxx6 = (~(U9jxx6 & B8knv6));
assign B8knv6 = (~(Jtpxx6 & Qtpxx6));
assign Qtpxx6 = (Xtpxx6 & Eupxx6);
assign Eupxx6 = (Vwlxx6 | Xg97x6);
assign Xtpxx6 = (Lupxx6 & Supxx6);
assign Supxx6 = (Xxlxx6 | Eh97x6);
assign Lupxx6 = (Wtlxx6 | Lh97x6);
assign Jtpxx6 = (R5pxx6 & Zupxx6);
assign Zupxx6 = (Fvlxx6 | Qg97x6);
assign Vspxx6 = (Adjxx6 | Br5jw6);
assign Br5jw6 = (Gvpxx6 & Nvpxx6);
assign Nvpxx6 = (Uvpxx6 & Bwpxx6);
assign Bwpxx6 = (Iwpxx6 & Pwpxx6);
assign Pwpxx6 = (Wwpxx6 & Dxpxx6);
assign Dxpxx6 = (~(X6kxx6 & vis_psp_o[18]));
assign Wwpxx6 = (~(E7kxx6 & vis_msp_o[18]));
assign Iwpxx6 = (Kxpxx6 & Rxpxx6);
assign Rxpxx6 = (~(Lfjxx6 & Pic7z6[18]));
assign Kxpxx6 = (~(Sfjxx6 & vis_r12_o[18]));
assign Uvpxx6 = (Yxpxx6 & Fypxx6);
assign Fypxx6 = (Mypxx6 & Typxx6);
assign Typxx6 = (~(Ngjxx6 & vis_r11_o[18]));
assign Mypxx6 = (~(Ugjxx6 & vis_r10_o[18]));
assign Yxpxx6 = (Azpxx6 & Hzpxx6);
assign Hzpxx6 = (~(Kijxx6 & vis_r7_o[18]));
assign Azpxx6 = (~(Rijxx6 & vis_r9_o[18]));
assign Gvpxx6 = (Ozpxx6 & Vzpxx6);
assign Vzpxx6 = (C0qxx6 & J0qxx6);
assign J0qxx6 = (Q0qxx6 & X0qxx6);
assign X0qxx6 = (~(Phjxx6 & vis_r8_o[18]));
assign Q0qxx6 = (~(Okjxx6 & vis_r6_o[18]));
assign C0qxx6 = (E1qxx6 & L1qxx6);
assign L1qxx6 = (~(Vkjxx6 & vis_r5_o[18]));
assign E1qxx6 = (~(Qljxx6 & vis_r4_o[18]));
assign Ozpxx6 = (S1qxx6 & Z1qxx6);
assign Z1qxx6 = (G2qxx6 & N2qxx6);
assign N2qxx6 = (~(Xljxx6 & vis_r3_o[18]));
assign G2qxx6 = (~(Nnjxx6 & vis_r0_o[18]));
assign S1qxx6 = (U2qxx6 & B3qxx6);
assign B3qxx6 = (~(Unjxx6 & vis_r2_o[18]));
assign U2qxx6 = (~(Smjxx6 & vis_r1_o[18]));
assign Trpxx6 = (I3qxx6 & P3qxx6);
assign P3qxx6 = (~(S8jxx6 & Cmm7z6[18]));
assign I3qxx6 = (~(K1i7z6[18] & Zs4ov6));
assign V7s7v6 = (~(W3qxx6 & D4qxx6));
assign D4qxx6 = (K4qxx6 & R4qxx6);
assign R4qxx6 = (~(Xzjxx6 & vis_pc_o[19]));
assign K4qxx6 = (Y4qxx6 & F5qxx6);
assign F5qxx6 = (~(U9jxx6 & L6knv6));
assign L6knv6 = (~(M5qxx6 & T5qxx6));
assign T5qxx6 = (A6qxx6 & H6qxx6);
assign H6qxx6 = (Vwlxx6 | Sa97x6);
assign A6qxx6 = (O6qxx6 & V6qxx6);
assign V6qxx6 = (Xxlxx6 | M797x6);
assign O6qxx6 = (Wtlxx6 | T797x6);
assign M5qxx6 = (R5pxx6 & C7qxx6);
assign C7qxx6 = (Fvlxx6 | Za97x6);
assign Y4qxx6 = (Adjxx6 | Rtbjw6);
assign Rtbjw6 = (J7qxx6 & Q7qxx6);
assign Q7qxx6 = (X7qxx6 & E8qxx6);
assign E8qxx6 = (L8qxx6 & S8qxx6);
assign S8qxx6 = (Z8qxx6 & G9qxx6);
assign G9qxx6 = (~(X6kxx6 & vis_psp_o[19]));
assign Z8qxx6 = (~(E7kxx6 & vis_msp_o[19]));
assign L8qxx6 = (N9qxx6 & U9qxx6);
assign U9qxx6 = (~(Lfjxx6 & Pic7z6[19]));
assign N9qxx6 = (~(Sfjxx6 & vis_r12_o[19]));
assign X7qxx6 = (Baqxx6 & Iaqxx6);
assign Iaqxx6 = (Paqxx6 & Waqxx6);
assign Waqxx6 = (~(Ngjxx6 & vis_r11_o[19]));
assign Paqxx6 = (~(Ugjxx6 & vis_r10_o[19]));
assign Baqxx6 = (Dbqxx6 & Kbqxx6);
assign Kbqxx6 = (~(Kijxx6 & vis_r7_o[19]));
assign Dbqxx6 = (~(Rijxx6 & vis_r9_o[19]));
assign J7qxx6 = (Rbqxx6 & Ybqxx6);
assign Ybqxx6 = (Fcqxx6 & Mcqxx6);
assign Mcqxx6 = (Tcqxx6 & Adqxx6);
assign Adqxx6 = (~(Phjxx6 & vis_r8_o[19]));
assign Tcqxx6 = (~(Okjxx6 & vis_r6_o[19]));
assign Fcqxx6 = (Hdqxx6 & Odqxx6);
assign Odqxx6 = (~(Vkjxx6 & vis_r5_o[19]));
assign Hdqxx6 = (~(Qljxx6 & vis_r4_o[19]));
assign Rbqxx6 = (Vdqxx6 & Ceqxx6);
assign Ceqxx6 = (Jeqxx6 & Qeqxx6);
assign Qeqxx6 = (~(Xljxx6 & vis_r3_o[19]));
assign Jeqxx6 = (~(Nnjxx6 & vis_r0_o[19]));
assign Vdqxx6 = (Xeqxx6 & Efqxx6);
assign Efqxx6 = (~(Unjxx6 & vis_r2_o[19]));
assign Xeqxx6 = (~(Smjxx6 & vis_r1_o[19]));
assign W3qxx6 = (Lfqxx6 & Sfqxx6);
assign Sfqxx6 = (~(S8jxx6 & Cmm7z6[19]));
assign Lfqxx6 = (~(K1i7z6[19] & Zs4ov6));
assign O7s7v6 = (~(Zfqxx6 & Ggqxx6));
assign Ggqxx6 = (Ngqxx6 & Ugqxx6);
assign Ugqxx6 = (~(Xzjxx6 & vis_pc_o[20]));
assign Ngqxx6 = (Bhqxx6 & Ihqxx6);
assign Ihqxx6 = (~(U9jxx6 & R2knv6));
assign R2knv6 = (~(Phqxx6 & Whqxx6));
assign Whqxx6 = (Diqxx6 & Kiqxx6);
assign Kiqxx6 = (Vwlxx6 | O197x6);
assign Diqxx6 = (Riqxx6 & Yiqxx6);
assign Yiqxx6 = (Xxlxx6 | Fjqxx6);
assign Riqxx6 = (Wtlxx6 | Mjqxx6);
assign Phqxx6 = (R5pxx6 & Tjqxx6);
assign Tjqxx6 = (Fvlxx6 | V197x6);
assign Bhqxx6 = (Adjxx6 | Dqp6x6);
assign Dqp6x6 = (Akqxx6 & Hkqxx6);
assign Hkqxx6 = (Okqxx6 & Vkqxx6);
assign Vkqxx6 = (Clqxx6 & Jlqxx6);
assign Jlqxx6 = (Qlqxx6 & Xlqxx6);
assign Xlqxx6 = (~(X6kxx6 & vis_psp_o[20]));
assign Qlqxx6 = (~(E7kxx6 & vis_msp_o[20]));
assign Clqxx6 = (Emqxx6 & Lmqxx6);
assign Lmqxx6 = (~(Lfjxx6 & Pic7z6[20]));
assign Emqxx6 = (~(Sfjxx6 & vis_r12_o[20]));
assign Okqxx6 = (Smqxx6 & Zmqxx6);
assign Zmqxx6 = (Gnqxx6 & Nnqxx6);
assign Nnqxx6 = (~(Ngjxx6 & vis_r11_o[20]));
assign Gnqxx6 = (~(Ugjxx6 & vis_r10_o[20]));
assign Smqxx6 = (Unqxx6 & Boqxx6);
assign Boqxx6 = (~(Kijxx6 & vis_r7_o[20]));
assign Unqxx6 = (~(Rijxx6 & vis_r9_o[20]));
assign Akqxx6 = (Ioqxx6 & Poqxx6);
assign Poqxx6 = (Woqxx6 & Dpqxx6);
assign Dpqxx6 = (Kpqxx6 & Rpqxx6);
assign Rpqxx6 = (~(Phjxx6 & vis_r8_o[20]));
assign Kpqxx6 = (~(Okjxx6 & vis_r6_o[20]));
assign Woqxx6 = (Ypqxx6 & Fqqxx6);
assign Fqqxx6 = (~(Vkjxx6 & vis_r5_o[20]));
assign Ypqxx6 = (~(Qljxx6 & vis_r4_o[20]));
assign Ioqxx6 = (Mqqxx6 & Tqqxx6);
assign Tqqxx6 = (Arqxx6 & Hrqxx6);
assign Hrqxx6 = (~(Xljxx6 & vis_r3_o[20]));
assign Arqxx6 = (~(Nnjxx6 & vis_r0_o[20]));
assign Mqqxx6 = (Orqxx6 & Vrqxx6);
assign Vrqxx6 = (~(Unjxx6 & vis_r2_o[20]));
assign Orqxx6 = (~(Smjxx6 & vis_r1_o[20]));
assign Zfqxx6 = (Csqxx6 & Jsqxx6);
assign Jsqxx6 = (~(S8jxx6 & Cmm7z6[20]));
assign Csqxx6 = (~(K1i7z6[20] & Zs4ov6));
assign H7s7v6 = (~(Qsqxx6 & Xsqxx6));
assign Xsqxx6 = (Etqxx6 & Ltqxx6);
assign Ltqxx6 = (~(Xzjxx6 & vis_pc_o[21]));
assign Etqxx6 = (Stqxx6 & Ztqxx6);
assign Ztqxx6 = (~(U9jxx6 & B1knv6));
assign B1knv6 = (~(Guqxx6 & Nuqxx6));
assign Nuqxx6 = (Uuqxx6 & Bvqxx6);
assign Bvqxx6 = (Vwlxx6 | Mt87x6);
assign Uuqxx6 = (Ivqxx6 & Pvqxx6);
assign Pvqxx6 = (Xxlxx6 | Wvqxx6);
assign Ivqxx6 = (Wtlxx6 | Dwqxx6);
assign Guqxx6 = (R5pxx6 & Kwqxx6);
assign Kwqxx6 = (Fvlxx6 | Tt87x6);
assign Stqxx6 = (Adjxx6 | Fcj6x6);
assign Fcj6x6 = (Rwqxx6 & Ywqxx6);
assign Ywqxx6 = (Fxqxx6 & Mxqxx6);
assign Mxqxx6 = (Txqxx6 & Ayqxx6);
assign Ayqxx6 = (Hyqxx6 & Oyqxx6);
assign Oyqxx6 = (~(X6kxx6 & vis_psp_o[21]));
assign Hyqxx6 = (~(E7kxx6 & vis_msp_o[21]));
assign Txqxx6 = (Vyqxx6 & Czqxx6);
assign Czqxx6 = (~(Lfjxx6 & Pic7z6[21]));
assign Vyqxx6 = (~(Sfjxx6 & vis_r12_o[21]));
assign Fxqxx6 = (Jzqxx6 & Qzqxx6);
assign Qzqxx6 = (Xzqxx6 & E0rxx6);
assign E0rxx6 = (~(Ngjxx6 & vis_r11_o[21]));
assign Xzqxx6 = (~(Ugjxx6 & vis_r10_o[21]));
assign Jzqxx6 = (L0rxx6 & S0rxx6);
assign S0rxx6 = (~(Kijxx6 & vis_r7_o[21]));
assign L0rxx6 = (~(Rijxx6 & vis_r9_o[21]));
assign Rwqxx6 = (Z0rxx6 & G1rxx6);
assign G1rxx6 = (N1rxx6 & U1rxx6);
assign U1rxx6 = (B2rxx6 & I2rxx6);
assign I2rxx6 = (~(Phjxx6 & vis_r8_o[21]));
assign B2rxx6 = (~(Okjxx6 & vis_r6_o[21]));
assign N1rxx6 = (P2rxx6 & W2rxx6);
assign W2rxx6 = (~(Vkjxx6 & vis_r5_o[21]));
assign P2rxx6 = (~(Qljxx6 & vis_r4_o[21]));
assign Z0rxx6 = (D3rxx6 & K3rxx6);
assign K3rxx6 = (R3rxx6 & Y3rxx6);
assign Y3rxx6 = (~(Xljxx6 & vis_r3_o[21]));
assign R3rxx6 = (~(Nnjxx6 & vis_r0_o[21]));
assign D3rxx6 = (F4rxx6 & M4rxx6);
assign M4rxx6 = (~(Unjxx6 & vis_r2_o[21]));
assign F4rxx6 = (~(Smjxx6 & vis_r1_o[21]));
assign Qsqxx6 = (T4rxx6 & A5rxx6);
assign A5rxx6 = (~(S8jxx6 & Cmm7z6[21]));
assign T4rxx6 = (~(K1i7z6[21] & Zs4ov6));
assign A7s7v6 = (~(H5rxx6 & O5rxx6));
assign O5rxx6 = (V5rxx6 & C6rxx6);
assign C6rxx6 = (~(Xzjxx6 & vis_pc_o[22]));
assign V5rxx6 = (J6rxx6 & Q6rxx6);
assign Q6rxx6 = (~(U9jxx6 & Lzjnv6));
assign Lzjnv6 = (~(X6rxx6 & E7rxx6));
assign E7rxx6 = (L7rxx6 & S7rxx6);
assign S7rxx6 = (Vwlxx6 | Kl87x6);
assign L7rxx6 = (Z7rxx6 & G8rxx6);
assign G8rxx6 = (Xxlxx6 | N8rxx6);
assign Z7rxx6 = (Wtlxx6 | U8rxx6);
assign X6rxx6 = (R5pxx6 & B9rxx6);
assign B9rxx6 = (Fvlxx6 | Rl87x6);
assign J6rxx6 = (Adjxx6 | B0m6x6);
assign B0m6x6 = (I9rxx6 & P9rxx6);
assign P9rxx6 = (W9rxx6 & Darxx6);
assign Darxx6 = (Karxx6 & Rarxx6);
assign Rarxx6 = (Yarxx6 & Fbrxx6);
assign Fbrxx6 = (~(X6kxx6 & vis_psp_o[22]));
assign Yarxx6 = (~(E7kxx6 & vis_msp_o[22]));
assign Karxx6 = (Mbrxx6 & Tbrxx6);
assign Tbrxx6 = (~(Lfjxx6 & Pic7z6[22]));
assign Mbrxx6 = (~(Sfjxx6 & vis_r12_o[22]));
assign W9rxx6 = (Acrxx6 & Hcrxx6);
assign Hcrxx6 = (Ocrxx6 & Vcrxx6);
assign Vcrxx6 = (~(Ngjxx6 & vis_r11_o[22]));
assign Ocrxx6 = (~(Ugjxx6 & vis_r10_o[22]));
assign Acrxx6 = (Cdrxx6 & Jdrxx6);
assign Jdrxx6 = (~(Kijxx6 & vis_r7_o[22]));
assign Cdrxx6 = (~(Rijxx6 & vis_r9_o[22]));
assign I9rxx6 = (Qdrxx6 & Xdrxx6);
assign Xdrxx6 = (Eerxx6 & Lerxx6);
assign Lerxx6 = (Serxx6 & Zerxx6);
assign Zerxx6 = (~(Phjxx6 & vis_r8_o[22]));
assign Serxx6 = (~(Okjxx6 & vis_r6_o[22]));
assign Eerxx6 = (Gfrxx6 & Nfrxx6);
assign Nfrxx6 = (~(Vkjxx6 & vis_r5_o[22]));
assign Gfrxx6 = (~(Qljxx6 & vis_r4_o[22]));
assign Qdrxx6 = (Ufrxx6 & Bgrxx6);
assign Bgrxx6 = (Igrxx6 & Pgrxx6);
assign Pgrxx6 = (~(Xljxx6 & vis_r3_o[22]));
assign Igrxx6 = (~(Nnjxx6 & vis_r0_o[22]));
assign Ufrxx6 = (Wgrxx6 & Dhrxx6);
assign Dhrxx6 = (~(Unjxx6 & vis_r2_o[22]));
assign Wgrxx6 = (~(Smjxx6 & vis_r1_o[22]));
assign H5rxx6 = (Khrxx6 & Rhrxx6);
assign Rhrxx6 = (~(S8jxx6 & Cmm7z6[22]));
assign Khrxx6 = (~(K1i7z6[22] & Zs4ov6));
assign T6s7v6 = (~(Yhrxx6 & Firxx6));
assign Firxx6 = (Mirxx6 & Tirxx6);
assign Tirxx6 = (~(Xzjxx6 & vis_pc_o[23]));
assign Mirxx6 = (Ajrxx6 & Hjrxx6);
assign Hjrxx6 = (~(U9jxx6 & Vxjnv6));
assign Vxjnv6 = (~(Ojrxx6 & Vjrxx6));
assign Vjrxx6 = (Ckrxx6 & Jkrxx6);
assign Jkrxx6 = (Vwlxx6 | Qkrxx6);
assign Vwlxx6 = (~(Oe9ov6 & Edh7z6[1]));
assign Oe9ov6 = (Xgmov6 ? H287x6 : Gaa7x6);
assign Ckrxx6 = (Xkrxx6 & Elrxx6);
assign Elrxx6 = (Xxlxx6 | Llrxx6);
assign Xxlxx6 = (~(Yc9ov6 & Edh7z6[1]));
assign Yc9ov6 = (Xgmov6 ? Gaa7x6 : Av77x6);
assign Xkrxx6 = (Wtlxx6 | Slrxx6);
assign Wtlxx6 = (~(Md9ov6 & Edh7z6[1]));
assign Md9ov6 = (Xgmov6 ? Av77x6 : Dca7x6);
assign Ojrxx6 = (R5pxx6 & Zlrxx6);
assign Zlrxx6 = (Fvlxx6 | Gmrxx6);
assign Fvlxx6 = (~(Cf9ov6 & Edh7z6[1]));
assign Cf9ov6 = (Xgmov6 ? Dca7x6 : H287x6);
assign Ajrxx6 = (Adjxx6 | Quo6x6);
assign Quo6x6 = (Nmrxx6 & Umrxx6);
assign Umrxx6 = (Bnrxx6 & Inrxx6);
assign Inrxx6 = (Pnrxx6 & Wnrxx6);
assign Wnrxx6 = (Dorxx6 & Korxx6);
assign Korxx6 = (~(X6kxx6 & vis_psp_o[23]));
assign Dorxx6 = (~(E7kxx6 & vis_msp_o[23]));
assign Pnrxx6 = (Rorxx6 & Yorxx6);
assign Yorxx6 = (~(Lfjxx6 & Pic7z6[23]));
assign Rorxx6 = (~(Sfjxx6 & vis_r12_o[23]));
assign Bnrxx6 = (Fprxx6 & Mprxx6);
assign Mprxx6 = (Tprxx6 & Aqrxx6);
assign Aqrxx6 = (~(Ngjxx6 & vis_r11_o[23]));
assign Tprxx6 = (~(Ugjxx6 & vis_r10_o[23]));
assign Fprxx6 = (Hqrxx6 & Oqrxx6);
assign Oqrxx6 = (~(Kijxx6 & vis_r7_o[23]));
assign Hqrxx6 = (~(Rijxx6 & vis_r9_o[23]));
assign Nmrxx6 = (Vqrxx6 & Crrxx6);
assign Crrxx6 = (Jrrxx6 & Qrrxx6);
assign Qrrxx6 = (Xrrxx6 & Esrxx6);
assign Esrxx6 = (~(Phjxx6 & vis_r8_o[23]));
assign Xrrxx6 = (~(Okjxx6 & vis_r6_o[23]));
assign Jrrxx6 = (Lsrxx6 & Ssrxx6);
assign Ssrxx6 = (~(Vkjxx6 & vis_r5_o[23]));
assign Lsrxx6 = (~(Qljxx6 & vis_r4_o[23]));
assign Vqrxx6 = (Zsrxx6 & Gtrxx6);
assign Gtrxx6 = (Ntrxx6 & Utrxx6);
assign Utrxx6 = (~(Xljxx6 & vis_r3_o[23]));
assign Ntrxx6 = (~(Nnjxx6 & vis_r0_o[23]));
assign Zsrxx6 = (Burxx6 & Iurxx6);
assign Iurxx6 = (~(Unjxx6 & vis_r2_o[23]));
assign Burxx6 = (~(Smjxx6 & vis_r1_o[23]));
assign Yhrxx6 = (Purxx6 & Wurxx6);
assign Wurxx6 = (~(S8jxx6 & Cmm7z6[23]));
assign Purxx6 = (~(K1i7z6[23] & Zs4ov6));
assign M6s7v6 = (~(Dvrxx6 & Kvrxx6));
assign Kvrxx6 = (Rvrxx6 & Yvrxx6);
assign Yvrxx6 = (~(Xzjxx6 & vis_pc_o[24]));
assign Rvrxx6 = (Fwrxx6 & Mwrxx6);
assign Mwrxx6 = (~(U9jxx6 & Fwjnv6));
assign Fwjnv6 = (~(Twrxx6 & Axrxx6));
assign Axrxx6 = (Hxrxx6 & Oxrxx6);
assign Oxrxx6 = (Kroxx6 | W4pxx6);
assign W4pxx6 = (!Td9ov6);
assign Hxrxx6 = (Vxrxx6 & Cyrxx6);
assign Cyrxx6 = (Fsoxx6 | Z487x6);
assign Z487x6 = (!Jf9ov6);
assign Vxrxx6 = (Npoxx6 | G587x6);
assign G587x6 = (!Ve9ov6);
assign Twrxx6 = (R5pxx6 & Jyrxx6);
assign Jyrxx6 = (Wqoxx6 | F6pxx6);
assign F6pxx6 = (!Fd9ov6);
assign Fwrxx6 = (Adjxx6 | Xf7jw6);
assign Xf7jw6 = (Qyrxx6 & Xyrxx6);
assign Xyrxx6 = (Ezrxx6 & Lzrxx6);
assign Lzrxx6 = (Szrxx6 & Zzrxx6);
assign Zzrxx6 = (G0sxx6 & N0sxx6);
assign N0sxx6 = (~(X6kxx6 & vis_psp_o[24]));
assign G0sxx6 = (~(E7kxx6 & vis_msp_o[24]));
assign Szrxx6 = (U0sxx6 & B1sxx6);
assign B1sxx6 = (~(Lfjxx6 & Pic7z6[24]));
assign U0sxx6 = (~(Sfjxx6 & vis_r12_o[24]));
assign Ezrxx6 = (I1sxx6 & P1sxx6);
assign P1sxx6 = (W1sxx6 & D2sxx6);
assign D2sxx6 = (~(Ngjxx6 & vis_r11_o[24]));
assign W1sxx6 = (~(Ugjxx6 & vis_r10_o[24]));
assign I1sxx6 = (K2sxx6 & R2sxx6);
assign R2sxx6 = (~(Kijxx6 & vis_r7_o[24]));
assign K2sxx6 = (~(Rijxx6 & vis_r9_o[24]));
assign Qyrxx6 = (Y2sxx6 & F3sxx6);
assign F3sxx6 = (M3sxx6 & T3sxx6);
assign T3sxx6 = (A4sxx6 & H4sxx6);
assign H4sxx6 = (~(Phjxx6 & vis_r8_o[24]));
assign A4sxx6 = (~(Okjxx6 & vis_r6_o[24]));
assign M3sxx6 = (O4sxx6 & V4sxx6);
assign V4sxx6 = (~(Vkjxx6 & vis_r5_o[24]));
assign O4sxx6 = (~(Qljxx6 & vis_r4_o[24]));
assign Y2sxx6 = (C5sxx6 & J5sxx6);
assign J5sxx6 = (Q5sxx6 & X5sxx6);
assign X5sxx6 = (~(Xljxx6 & vis_r3_o[24]));
assign Q5sxx6 = (~(Nnjxx6 & vis_r0_o[24]));
assign C5sxx6 = (E6sxx6 & L6sxx6);
assign L6sxx6 = (~(Unjxx6 & vis_r2_o[24]));
assign E6sxx6 = (~(Smjxx6 & vis_r1_o[24]));
assign Dvrxx6 = (S6sxx6 & Z6sxx6);
assign Z6sxx6 = (~(S8jxx6 & Cmm7z6[24]));
assign S6sxx6 = (~(K1i7z6[24] & Zs4ov6));
assign F6s7v6 = (~(G7sxx6 & N7sxx6));
assign N7sxx6 = (U7sxx6 & B8sxx6);
assign B8sxx6 = (~(Xzjxx6 & vis_pc_o[25]));
assign U7sxx6 = (I8sxx6 & P8sxx6);
assign P8sxx6 = (~(U9jxx6 & Pujnv6));
assign Pujnv6 = (~(W8sxx6 & D9sxx6));
assign D9sxx6 = (K9sxx6 & R9sxx6);
assign R9sxx6 = (Kroxx6 | Cu97x6);
assign Cu97x6 = (!Ex77x6);
assign K9sxx6 = (Y9sxx6 & Fasxx6);
assign Fasxx6 = (Fsoxx6 | Iipxx6);
assign Iipxx6 = (!Ab67x6);
assign Y9sxx6 = (Npoxx6 | Pipxx6);
assign Pipxx6 = (!Ob67x6);
assign W8sxx6 = (R5pxx6 & Masxx6);
assign Masxx6 = (Wqoxx6 | Ju97x6);
assign Ju97x6 = (!Vv77x6);
assign I8sxx6 = (Adjxx6 | Dk6jw6);
assign Dk6jw6 = (Tasxx6 & Absxx6);
assign Absxx6 = (Hbsxx6 & Obsxx6);
assign Obsxx6 = (Vbsxx6 & Ccsxx6);
assign Ccsxx6 = (Jcsxx6 & Qcsxx6);
assign Qcsxx6 = (~(X6kxx6 & vis_psp_o[25]));
assign Jcsxx6 = (~(E7kxx6 & vis_msp_o[25]));
assign Vbsxx6 = (Xcsxx6 & Edsxx6);
assign Edsxx6 = (~(Lfjxx6 & Pic7z6[25]));
assign Xcsxx6 = (~(Sfjxx6 & vis_r12_o[25]));
assign Hbsxx6 = (Ldsxx6 & Sdsxx6);
assign Sdsxx6 = (Zdsxx6 & Gesxx6);
assign Gesxx6 = (~(Ngjxx6 & vis_r11_o[25]));
assign Zdsxx6 = (~(Ugjxx6 & vis_r10_o[25]));
assign Ldsxx6 = (Nesxx6 & Uesxx6);
assign Uesxx6 = (~(Kijxx6 & vis_r7_o[25]));
assign Nesxx6 = (~(Rijxx6 & vis_r9_o[25]));
assign Tasxx6 = (Bfsxx6 & Ifsxx6);
assign Ifsxx6 = (Pfsxx6 & Wfsxx6);
assign Wfsxx6 = (Dgsxx6 & Kgsxx6);
assign Kgsxx6 = (~(Phjxx6 & vis_r8_o[25]));
assign Dgsxx6 = (~(Okjxx6 & vis_r6_o[25]));
assign Pfsxx6 = (Rgsxx6 & Ygsxx6);
assign Ygsxx6 = (~(Vkjxx6 & vis_r5_o[25]));
assign Rgsxx6 = (~(Qljxx6 & vis_r4_o[25]));
assign Bfsxx6 = (Fhsxx6 & Mhsxx6);
assign Mhsxx6 = (Thsxx6 & Aisxx6);
assign Aisxx6 = (~(Xljxx6 & vis_r3_o[25]));
assign Thsxx6 = (~(Nnjxx6 & vis_r0_o[25]));
assign Fhsxx6 = (Hisxx6 & Oisxx6);
assign Oisxx6 = (~(Unjxx6 & vis_r2_o[25]));
assign Hisxx6 = (~(Smjxx6 & vis_r1_o[25]));
assign G7sxx6 = (Visxx6 & Cjsxx6);
assign Cjsxx6 = (~(S8jxx6 & Cmm7z6[25]));
assign Visxx6 = (~(K1i7z6[25] & Zs4ov6));
assign Y5s7v6 = (~(Jjsxx6 & Qjsxx6));
assign Qjsxx6 = (Xjsxx6 & Eksxx6);
assign Eksxx6 = (~(Xzjxx6 & vis_pc_o[26]));
assign Xjsxx6 = (Lksxx6 & Sksxx6);
assign Sksxx6 = (~(U9jxx6 & Zsjnv6));
assign Zsjnv6 = (~(Zksxx6 & Glsxx6));
assign Glsxx6 = (Nlsxx6 & Ulsxx6);
assign Ulsxx6 = (Kroxx6 | Xg97x6);
assign Xg97x6 = (!Icfov6);
assign Nlsxx6 = (Bmsxx6 & Imsxx6);
assign Imsxx6 = (Eh97x6 | Fsoxx6);
assign Eh97x6 = (!Kdfov6);
assign Bmsxx6 = (Lh97x6 | Npoxx6);
assign Lh97x6 = (!Ddfov6);
assign Zksxx6 = (R5pxx6 & Pmsxx6);
assign Pmsxx6 = (Wqoxx6 | Qg97x6);
assign Qg97x6 = (!Bcfov6);
assign Lksxx6 = (Adjxx6 | U0s6x6);
assign U0s6x6 = (Wmsxx6 & Dnsxx6);
assign Dnsxx6 = (Knsxx6 & Rnsxx6);
assign Rnsxx6 = (Ynsxx6 & Fosxx6);
assign Fosxx6 = (Mosxx6 & Tosxx6);
assign Tosxx6 = (~(X6kxx6 & vis_psp_o[26]));
assign Mosxx6 = (~(E7kxx6 & vis_msp_o[26]));
assign Ynsxx6 = (Apsxx6 & Hpsxx6);
assign Hpsxx6 = (~(Lfjxx6 & Pic7z6[26]));
assign Apsxx6 = (~(Sfjxx6 & vis_r12_o[26]));
assign Knsxx6 = (Opsxx6 & Vpsxx6);
assign Vpsxx6 = (Cqsxx6 & Jqsxx6);
assign Jqsxx6 = (~(Ngjxx6 & vis_r11_o[26]));
assign Cqsxx6 = (~(Ugjxx6 & vis_r10_o[26]));
assign Opsxx6 = (Qqsxx6 & Xqsxx6);
assign Xqsxx6 = (~(Kijxx6 & vis_r7_o[26]));
assign Qqsxx6 = (~(Rijxx6 & vis_r9_o[26]));
assign Wmsxx6 = (Ersxx6 & Lrsxx6);
assign Lrsxx6 = (Srsxx6 & Zrsxx6);
assign Zrsxx6 = (Gssxx6 & Nssxx6);
assign Nssxx6 = (~(Phjxx6 & vis_r8_o[26]));
assign Gssxx6 = (~(Okjxx6 & vis_r6_o[26]));
assign Srsxx6 = (Vssxx6 & Dtsxx6);
assign Dtsxx6 = (~(Vkjxx6 & vis_r5_o[26]));
assign Vssxx6 = (~(Qljxx6 & vis_r4_o[26]));
assign Ersxx6 = (Ltsxx6 & Ttsxx6);
assign Ttsxx6 = (Busxx6 & Jusxx6);
assign Jusxx6 = (~(Xljxx6 & vis_r3_o[26]));
assign Busxx6 = (~(Nnjxx6 & vis_r0_o[26]));
assign Ltsxx6 = (Rusxx6 & Zusxx6);
assign Zusxx6 = (~(Unjxx6 & vis_r2_o[26]));
assign Rusxx6 = (~(Smjxx6 & vis_r1_o[26]));
assign Jjsxx6 = (Hvsxx6 & Pvsxx6);
assign Pvsxx6 = (~(S8jxx6 & Cmm7z6[26]));
assign Hvsxx6 = (~(K1i7z6[26] & Zs4ov6));
assign R5s7v6 = (~(Xvsxx6 & Fwsxx6));
assign Fwsxx6 = (Nwsxx6 & Vwsxx6);
assign Vwsxx6 = (~(Xzjxx6 & vis_pc_o[27]));
assign Nwsxx6 = (Dxsxx6 & Lxsxx6);
assign Lxsxx6 = (~(U9jxx6 & Jrjnv6));
assign Jrjnv6 = (~(Txsxx6 & Bysxx6));
assign Bysxx6 = (Jysxx6 & Rysxx6);
assign Rysxx6 = (Sa97x6 | Kroxx6);
assign Sa97x6 = (!Mmlov6);
assign Jysxx6 = (Zysxx6 & Hzsxx6);
assign Hzsxx6 = (M797x6 | Fsoxx6);
assign M797x6 = (!Onlov6);
assign Zysxx6 = (T797x6 | Npoxx6);
assign T797x6 = (!Hnlov6);
assign Txsxx6 = (R5pxx6 & Pzsxx6);
assign Pzsxx6 = (Za97x6 | Wqoxx6);
assign Za97x6 = (!Fmlov6);
assign Dxsxx6 = (Adjxx6 | Ers6x6);
assign Ers6x6 = (Xzsxx6 & F0txx6);
assign F0txx6 = (N0txx6 & V0txx6);
assign V0txx6 = (D1txx6 & L1txx6);
assign L1txx6 = (T1txx6 & B2txx6);
assign B2txx6 = (~(X6kxx6 & vis_psp_o[27]));
assign T1txx6 = (~(E7kxx6 & vis_msp_o[27]));
assign D1txx6 = (J2txx6 & R2txx6);
assign R2txx6 = (~(Lfjxx6 & Pic7z6[27]));
assign J2txx6 = (~(Sfjxx6 & vis_r12_o[27]));
assign N0txx6 = (Z2txx6 & H3txx6);
assign H3txx6 = (P3txx6 & X3txx6);
assign X3txx6 = (~(Ngjxx6 & vis_r11_o[27]));
assign P3txx6 = (~(Ugjxx6 & vis_r10_o[27]));
assign Z2txx6 = (F4txx6 & N4txx6);
assign N4txx6 = (~(Kijxx6 & vis_r7_o[27]));
assign F4txx6 = (~(Rijxx6 & vis_r9_o[27]));
assign Xzsxx6 = (V4txx6 & D5txx6);
assign D5txx6 = (L5txx6 & T5txx6);
assign T5txx6 = (B6txx6 & J6txx6);
assign J6txx6 = (~(Phjxx6 & vis_r8_o[27]));
assign B6txx6 = (~(Okjxx6 & vis_r6_o[27]));
assign L5txx6 = (R6txx6 & Z6txx6);
assign Z6txx6 = (~(Vkjxx6 & vis_r5_o[27]));
assign R6txx6 = (~(Qljxx6 & vis_r4_o[27]));
assign V4txx6 = (H7txx6 & P7txx6);
assign P7txx6 = (X7txx6 & F8txx6);
assign F8txx6 = (~(Xljxx6 & vis_r3_o[27]));
assign X7txx6 = (~(Nnjxx6 & vis_r0_o[27]));
assign H7txx6 = (N8txx6 & V8txx6);
assign V8txx6 = (~(Unjxx6 & vis_r2_o[27]));
assign N8txx6 = (~(Smjxx6 & vis_r1_o[27]));
assign Xvsxx6 = (D9txx6 & L9txx6);
assign L9txx6 = (~(S8jxx6 & Cmm7z6[27]));
assign D9txx6 = (~(K1i7z6[27] & Zs4ov6));
assign K5s7v6 = (~(T9txx6 & Batxx6));
assign Batxx6 = (Jatxx6 & Ratxx6);
assign Ratxx6 = (~(Xzjxx6 & vis_pc_o[28]));
assign Jatxx6 = (Zatxx6 & Hbtxx6);
assign Hbtxx6 = (~(U9jxx6 & Tpjnv6));
assign Tpjnv6 = (~(Pbtxx6 & Xbtxx6));
assign Xbtxx6 = (Fctxx6 & Nctxx6);
assign Nctxx6 = (O197x6 | Kroxx6);
assign O197x6 = (!Cb77x6);
assign Fctxx6 = (Vctxx6 & Ddtxx6);
assign Ddtxx6 = (Fjqxx6 | Fsoxx6);
assign Fjqxx6 = (!Tw57x6);
assign Vctxx6 = (Mjqxx6 | Npoxx6);
assign Mjqxx6 = (!Ax57x6);
assign Pbtxx6 = (R5pxx6 & Ldtxx6);
assign Ldtxx6 = (V197x6 | Wqoxx6);
assign V197x6 = (!T977x6);
assign Zatxx6 = (Adjxx6 | Zct6x6);
assign Zct6x6 = (Tdtxx6 & Betxx6);
assign Betxx6 = (Jetxx6 & Retxx6);
assign Retxx6 = (Zetxx6 & Hftxx6);
assign Hftxx6 = (Pftxx6 & Xftxx6);
assign Xftxx6 = (~(X6kxx6 & vis_psp_o[28]));
assign Pftxx6 = (~(E7kxx6 & vis_msp_o[28]));
assign Zetxx6 = (Fgtxx6 & Ngtxx6);
assign Ngtxx6 = (~(Lfjxx6 & Pic7z6[28]));
assign Fgtxx6 = (~(Sfjxx6 & vis_r12_o[28]));
assign Jetxx6 = (Vgtxx6 & Dhtxx6);
assign Dhtxx6 = (Lhtxx6 & Thtxx6);
assign Thtxx6 = (~(Ngjxx6 & vis_r11_o[28]));
assign Lhtxx6 = (~(Ugjxx6 & vis_r10_o[28]));
assign Vgtxx6 = (Bitxx6 & Jitxx6);
assign Jitxx6 = (~(Kijxx6 & vis_r7_o[28]));
assign Bitxx6 = (~(Rijxx6 & vis_r9_o[28]));
assign Tdtxx6 = (Ritxx6 & Zitxx6);
assign Zitxx6 = (Hjtxx6 & Pjtxx6);
assign Pjtxx6 = (Xjtxx6 & Fktxx6);
assign Fktxx6 = (~(Phjxx6 & vis_r8_o[28]));
assign Xjtxx6 = (~(Okjxx6 & vis_r6_o[28]));
assign Hjtxx6 = (Nktxx6 & Vktxx6);
assign Vktxx6 = (~(Vkjxx6 & vis_r5_o[28]));
assign Nktxx6 = (~(Qljxx6 & vis_r4_o[28]));
assign Ritxx6 = (Dltxx6 & Lltxx6);
assign Lltxx6 = (Tltxx6 & Bmtxx6);
assign Bmtxx6 = (~(Xljxx6 & vis_r3_o[28]));
assign Tltxx6 = (~(Nnjxx6 & vis_r0_o[28]));
assign Dltxx6 = (Jmtxx6 & Rmtxx6);
assign Rmtxx6 = (~(Unjxx6 & vis_r2_o[28]));
assign Jmtxx6 = (~(Smjxx6 & vis_r1_o[28]));
assign T9txx6 = (Zmtxx6 & Hntxx6);
assign Hntxx6 = (~(S8jxx6 & Cmm7z6[28]));
assign Zmtxx6 = (~(K1i7z6[28] & Zs4ov6));
assign D5s7v6 = (~(Pntxx6 & Xntxx6));
assign Xntxx6 = (Fotxx6 & Notxx6);
assign Notxx6 = (~(U9jxx6 & Dojnv6));
assign Dojnv6 = (~(Votxx6 & Dptxx6));
assign Dptxx6 = (Lptxx6 & Tptxx6);
assign Tptxx6 = (Mt87x6 | Kroxx6);
assign Mt87x6 = (!C477x6);
assign Lptxx6 = (Bqtxx6 & Jqtxx6);
assign Jqtxx6 = (Wvqxx6 | Fsoxx6);
assign Wvqxx6 = (!Qr57x6);
assign Bqtxx6 = (Dwqxx6 | Npoxx6);
assign Dwqxx6 = (!Xr57x6);
assign Votxx6 = (R5pxx6 & Rqtxx6);
assign Rqtxx6 = (Tt87x6 | Wqoxx6);
assign Tt87x6 = (!T277x6);
assign Fotxx6 = (Zqtxx6 & Wgkxx6);
assign Zqtxx6 = (Adjxx6 | Cybov6);
assign Cybov6 = (Hrtxx6 & Prtxx6);
assign Prtxx6 = (Xrtxx6 & Fstxx6);
assign Fstxx6 = (Nstxx6 & Vstxx6);
assign Vstxx6 = (Dttxx6 & Lttxx6);
assign Lttxx6 = (~(X6kxx6 & vis_psp_o[29]));
assign Dttxx6 = (~(E7kxx6 & vis_msp_o[29]));
assign Nstxx6 = (Tttxx6 & Butxx6);
assign Butxx6 = (~(Lfjxx6 & Pic7z6[29]));
assign Tttxx6 = (~(Sfjxx6 & vis_r12_o[29]));
assign Xrtxx6 = (Jutxx6 & Rutxx6);
assign Rutxx6 = (Zutxx6 & Hvtxx6);
assign Hvtxx6 = (~(Ngjxx6 & vis_r11_o[29]));
assign Zutxx6 = (~(Ugjxx6 & vis_r10_o[29]));
assign Jutxx6 = (Pvtxx6 & Xvtxx6);
assign Xvtxx6 = (~(Kijxx6 & vis_r7_o[29]));
assign Pvtxx6 = (~(Rijxx6 & vis_r9_o[29]));
assign Hrtxx6 = (Fwtxx6 & Nwtxx6);
assign Nwtxx6 = (Vwtxx6 & Dxtxx6);
assign Dxtxx6 = (Lxtxx6 & Txtxx6);
assign Txtxx6 = (~(Phjxx6 & vis_r8_o[29]));
assign Lxtxx6 = (~(Okjxx6 & vis_r6_o[29]));
assign Vwtxx6 = (Bytxx6 & Jytxx6);
assign Jytxx6 = (~(Vkjxx6 & vis_r5_o[29]));
assign Bytxx6 = (~(Qljxx6 & vis_r4_o[29]));
assign Fwtxx6 = (Rytxx6 & Zytxx6);
assign Zytxx6 = (Hztxx6 & Pztxx6);
assign Pztxx6 = (~(Xljxx6 & vis_r3_o[29]));
assign Hztxx6 = (~(Nnjxx6 & vis_r0_o[29]));
assign Rytxx6 = (Xztxx6 & F0uxx6);
assign F0uxx6 = (~(Unjxx6 & vis_r2_o[29]));
assign Xztxx6 = (~(Smjxx6 & vis_r1_o[29]));
assign Pntxx6 = (N0uxx6 & V0uxx6);
assign V0uxx6 = (~(K1i7z6[29] & Zs4ov6));
assign N0uxx6 = (D1uxx6 & L1uxx6);
assign L1uxx6 = (~(Xzjxx6 & vis_pc_o[29]));
assign D1uxx6 = (~(S8jxx6 & Cmm7z6[29]));
assign W4s7v6 = (~(T1uxx6 & B2uxx6));
assign B2uxx6 = (J2uxx6 & R2uxx6);
assign R2uxx6 = (~(U9jxx6 & Xkjnv6));
assign Xkjnv6 = (~(Z2uxx6 & H3uxx6));
assign H3uxx6 = (P3uxx6 & X3uxx6);
assign X3uxx6 = (Kl87x6 | Kroxx6);
assign Kl87x6 = (!Cx67x6);
assign P3uxx6 = (F4uxx6 & N4uxx6);
assign N4uxx6 = (N8rxx6 | Fsoxx6);
assign N8rxx6 = (!Nm57x6);
assign F4uxx6 = (U8rxx6 | Npoxx6);
assign U8rxx6 = (!Um57x6);
assign Z2uxx6 = (R5pxx6 & V4uxx6);
assign V4uxx6 = (Rl87x6 | Wqoxx6);
assign Rl87x6 = (!Tv67x6);
assign J2uxx6 = (D5uxx6 & Wgkxx6);
assign D5uxx6 = (Adjxx6 | F1u6x6);
assign F1u6x6 = (L5uxx6 & T5uxx6);
assign T5uxx6 = (B6uxx6 & J6uxx6);
assign J6uxx6 = (R6uxx6 & Z6uxx6);
assign Z6uxx6 = (H7uxx6 & P7uxx6);
assign P7uxx6 = (~(X6kxx6 & vis_psp_o[30]));
assign H7uxx6 = (~(E7kxx6 & vis_msp_o[30]));
assign R6uxx6 = (X7uxx6 & F8uxx6);
assign F8uxx6 = (~(Lfjxx6 & Pic7z6[30]));
assign X7uxx6 = (~(Sfjxx6 & vis_r12_o[30]));
assign B6uxx6 = (N8uxx6 & V8uxx6);
assign V8uxx6 = (D9uxx6 & L9uxx6);
assign L9uxx6 = (~(Ngjxx6 & vis_r11_o[30]));
assign D9uxx6 = (~(Ugjxx6 & vis_r10_o[30]));
assign N8uxx6 = (T9uxx6 & Bauxx6);
assign Bauxx6 = (~(Kijxx6 & vis_r7_o[30]));
assign T9uxx6 = (~(Rijxx6 & vis_r9_o[30]));
assign L5uxx6 = (Jauxx6 & Rauxx6);
assign Rauxx6 = (Zauxx6 & Hbuxx6);
assign Hbuxx6 = (Pbuxx6 & Xbuxx6);
assign Xbuxx6 = (~(Phjxx6 & vis_r8_o[30]));
assign Pbuxx6 = (~(Okjxx6 & vis_r6_o[30]));
assign Zauxx6 = (Fcuxx6 & Ncuxx6);
assign Ncuxx6 = (~(Vkjxx6 & vis_r5_o[30]));
assign Fcuxx6 = (~(Qljxx6 & vis_r4_o[30]));
assign Jauxx6 = (Vcuxx6 & Dduxx6);
assign Dduxx6 = (Lduxx6 & Tduxx6);
assign Tduxx6 = (~(Xljxx6 & vis_r3_o[30]));
assign Lduxx6 = (~(Nnjxx6 & vis_r0_o[30]));
assign Vcuxx6 = (Beuxx6 & Jeuxx6);
assign Jeuxx6 = (~(Unjxx6 & vis_r2_o[30]));
assign Beuxx6 = (~(Smjxx6 & vis_r1_o[30]));
assign T1uxx6 = (Reuxx6 & Zeuxx6);
assign Zeuxx6 = (~(K1i7z6[30] & Zs4ov6));
assign Reuxx6 = (Hfuxx6 & Pfuxx6);
assign Pfuxx6 = (~(Xzjxx6 & vis_pc_o[30]));
assign Hfuxx6 = (~(S8jxx6 & Cmm7z6[30]));
assign P4s7v6 = (~(Xfuxx6 & Fguxx6));
assign Fguxx6 = (Nguxx6 & Vguxx6);
assign Vguxx6 = (~(Xzjxx6 & vis_pc_o[31]));
assign Xzjxx6 = (Dhuxx6 & Lhuxx6);
assign Dhuxx6 = (~(A2u6x6 | Thuxx6));
assign A2u6x6 = (!R0u6x6);
assign Nguxx6 = (Biuxx6 & Wgkxx6);
assign Wgkxx6 = (~(Jiuxx6 & Hyhhw6));
assign Jiuxx6 = (Riuxx6 & Vqihw6);
assign Biuxx6 = (Adjxx6 | B1cov6);
assign B1cov6 = (Ziuxx6 & Hjuxx6);
assign Hjuxx6 = (Pjuxx6 & Xjuxx6);
assign Xjuxx6 = (Fkuxx6 & Nkuxx6);
assign Nkuxx6 = (Vkuxx6 & Dluxx6);
assign Dluxx6 = (~(X6kxx6 & vis_psp_o[31]));
assign X6kxx6 = (~(Lluxx6 | Ix27x6));
assign Vkuxx6 = (~(E7kxx6 & vis_msp_o[31]));
assign E7kxx6 = (~(Tluxx6 | Lluxx6));
assign Fkuxx6 = (Bmuxx6 & Jmuxx6);
assign Jmuxx6 = (~(Lfjxx6 & Pic7z6[31]));
assign Lfjxx6 = (Rmuxx6 & Zmuxx6);
assign Bmuxx6 = (~(Sfjxx6 & vis_r12_o[31]));
assign Sfjxx6 = (Hnuxx6 & Zmuxx6);
assign Pjuxx6 = (Pnuxx6 & Xnuxx6);
assign Xnuxx6 = (Fouxx6 & Nouxx6);
assign Nouxx6 = (~(Ngjxx6 & vis_r11_o[31]));
assign Ngjxx6 = (Vouxx6 & Dpuxx6);
assign Fouxx6 = (~(Ugjxx6 & vis_r10_o[31]));
assign Ugjxx6 = (Vouxx6 & Zmuxx6);
assign Pnuxx6 = (Lpuxx6 & Tpuxx6);
assign Tpuxx6 = (~(Kijxx6 & vis_r7_o[31]));
assign Kijxx6 = (Rmuxx6 & Bquxx6);
assign Lpuxx6 = (~(Rijxx6 & vis_r9_o[31]));
assign Rijxx6 = (Dpuxx6 & Jquxx6);
assign Ziuxx6 = (Rquxx6 & Zquxx6);
assign Zquxx6 = (Hruxx6 & Pruxx6);
assign Pruxx6 = (Xruxx6 & Fsuxx6);
assign Fsuxx6 = (~(Phjxx6 & vis_r8_o[31]));
assign Phjxx6 = (Jquxx6 & Zmuxx6);
assign Zmuxx6 = (~(Xgfhw6 | Nsuxx6));
assign Xruxx6 = (~(Okjxx6 & vis_r6_o[31]));
assign Okjxx6 = (Rmuxx6 & Vsuxx6);
assign Rmuxx6 = (Tluxx6 & Bjfhw6);
assign Hruxx6 = (Dtuxx6 & Ltuxx6);
assign Ltuxx6 = (~(Vkjxx6 & vis_r5_o[31]));
assign Vkjxx6 = (Hnuxx6 & Bquxx6);
assign Dtuxx6 = (~(Qljxx6 & vis_r4_o[31]));
assign Qljxx6 = (Hnuxx6 & Vsuxx6);
assign Hnuxx6 = (Ix27x6 & Bjfhw6);
assign Ix27x6 = (!Tluxx6);
assign Rquxx6 = (Ttuxx6 & Buuxx6);
assign Buuxx6 = (Juuxx6 & Ruuxx6);
assign Ruuxx6 = (~(Xljxx6 & vis_r3_o[31]));
assign Xljxx6 = (Vouxx6 & Bquxx6);
assign Juuxx6 = (~(Nnjxx6 & vis_r0_o[31]));
assign Nnjxx6 = (Vsuxx6 & Jquxx6);
assign Ttuxx6 = (Zuuxx6 & Hvuxx6);
assign Hvuxx6 = (~(Unjxx6 & vis_r2_o[31]));
assign Unjxx6 = (Vouxx6 & Vsuxx6);
assign Vsuxx6 = (~(Uifhw6 | Xgfhw6));
assign Vouxx6 = (Pvuxx6 & Tluxx6);
assign Zuuxx6 = (~(Smjxx6 & vis_r1_o[31]));
assign Smjxx6 = (Jquxx6 & Bquxx6);
assign Bquxx6 = (~(Uifhw6 | Xvuxx6));
assign Jquxx6 = (~(Bjfhw6 | Tluxx6));
assign Tluxx6 = (~(Vrjxx6 & Fwuxx6));
assign Fwuxx6 = (~(Csjxx6 & Tqq6x6));
assign Tqq6x6 = (~(Nwuxx6 & Vwuxx6));
assign Vwuxx6 = (~(Dxuxx6 & Lxuxx6));
assign Dxuxx6 = (F02nv6 ? Qij7z6[1] : Ovbdt6);
assign Nwuxx6 = (Lxuxx6 | Mz27x6);
assign Mz27x6 = (~(Txuxx6 & Byuxx6));
assign Byuxx6 = (~(Jyuxx6 & Ad9iw6));
assign Jyuxx6 = (~(Hd9iw6 | Q0wnv6));
assign Txuxx6 = (Ryuxx6 | Jjbdt6);
assign Ryuxx6 = (~(Ad9iw6 | Hd9iw6));
assign Hd9iw6 = (Zyuxx6 & Hzuxx6);
assign Hzuxx6 = (Pzuxx6 & Xzuxx6);
assign Xzuxx6 = (~(Tx1jw6 | Qm0jw6));
assign Pzuxx6 = (~(Jti6x6 | Ddo6x6));
assign Zyuxx6 = (F0vxx6 & N0vxx6);
assign N0vxx6 = (~(Nob7z6[1] & Rslov6));
assign F0vxx6 = (V0vxx6 & D1vxx6);
assign D1vxx6 = (~(Rslov6 & L1vxx6));
assign L1vxx6 = (~(T1vxx6 & Flliw6));
assign T1vxx6 = (Gpliw6 & Xxjov6);
assign V0vxx6 = (~(Nob7z6[4] & Rslov6));
assign Lxuxx6 = (~(B2vxx6 & Yy27x6));
assign Yy27x6 = (~(J2vxx6 & Qij7z6[4]));
assign J2vxx6 = (R2vxx6 & F02nv6);
assign B2vxx6 = (~(Z2vxx6 & H3vxx6));
assign H3vxx6 = (P3vxx6 & W6u6x6);
assign Z2vxx6 = (X3vxx6 & Ansov6);
assign Ansov6 = (F4vxx6 & Jgtov6);
assign Adjxx6 = (~(N4vxx6 & Lhuxx6));
assign N4vxx6 = (~(Thuxx6 | R0u6x6));
assign R0u6x6 = (~(Lluxx6 | Vrjxx6));
assign Lluxx6 = (!Csjxx6);
assign Csjxx6 = (Dpuxx6 & Bjfhw6);
assign Dpuxx6 = (Uifhw6 & Xgfhw6);
assign Xfuxx6 = (V4vxx6 & D5vxx6);
assign D5vxx6 = (~(K1i7z6[31] & Zs4ov6));
assign V4vxx6 = (L5vxx6 & T5vxx6);
assign T5vxx6 = (~(U9jxx6 & Hjjnv6));
assign Hjjnv6 = (~(B6vxx6 & J6vxx6));
assign J6vxx6 = (R6vxx6 & Z6vxx6);
assign Z6vxx6 = (Kroxx6 | Qkrxx6);
assign Qkrxx6 = (!Hp67x6);
assign Kroxx6 = (H7vxx6 & P7vxx6);
assign H7vxx6 = (X7vxx6 | Xgmov6);
assign R6vxx6 = (F8vxx6 & N8vxx6);
assign N8vxx6 = (Fsoxx6 | Llrxx6);
assign Llrxx6 = (!Dh57x6);
assign Fsoxx6 = (V8vxx6 & D9vxx6);
assign V8vxx6 = (~(L9vxx6 & Xgmov6));
assign F8vxx6 = (Npoxx6 | Slrxx6);
assign Slrxx6 = (!Rh57x6);
assign Npoxx6 = (T9vxx6 & Bavxx6);
assign T9vxx6 = (~(L9vxx6 & No7et6));
assign B6vxx6 = (R5pxx6 & Javxx6);
assign Javxx6 = (Wqoxx6 | Gmrxx6);
assign Gmrxx6 = (!Kn67x6);
assign Wqoxx6 = (Ravxx6 & Zavxx6);
assign Ravxx6 = (X7vxx6 | No7et6);
assign R5pxx6 = (Hbvxx6 & Pbvxx6);
assign Pbvxx6 = (Xbvxx6 & Fcvxx6);
assign Fcvxx6 = (~(Rh57x6 & Ncvxx6));
assign Ncvxx6 = (~(Vcvxx6 & Ddvxx6));
assign Ddvxx6 = (~(Ldvxx6 & Vt2et6));
assign Ldvxx6 = (Itlxx6 & H287x6);
assign Vcvxx6 = (Tdvxx6 | Aea7x6);
assign Aea7x6 = (!Dca7x6);
assign Xbvxx6 = (Bevxx6 & Jevxx6);
assign Jevxx6 = (~(Dh57x6 & Revxx6));
assign Revxx6 = (~(Zevxx6 & Hfvxx6));
assign Hfvxx6 = (~(Pfvxx6 & Vt2et6));
assign Pfvxx6 = (Itlxx6 & Dca7x6);
assign Zevxx6 = (Tdvxx6 | Yca7x6);
assign Yca7x6 = (!Av77x6);
assign Bevxx6 = (~(Kn67x6 & Xfvxx6));
assign Xfvxx6 = (~(Fgvxx6 & Ngvxx6));
assign Ngvxx6 = (~(Vgvxx6 & Vt2et6));
assign Vgvxx6 = (Itlxx6 & Gaa7x6);
assign Fgvxx6 = (Tdvxx6 | Iba7x6);
assign Iba7x6 = (!H287x6);
assign Hbvxx6 = (Jbmxx6 & Dhvxx6);
assign Dhvxx6 = (~(Hp67x6 & Lhvxx6));
assign Lhvxx6 = (~(Thvxx6 & Bivxx6));
assign Bivxx6 = (~(Jivxx6 & Vt2et6));
assign Jivxx6 = (Itlxx6 & Av77x6);
assign Itlxx6 = (Bqoxx6 & No7et6);
assign Thvxx6 = (Tdvxx6 | Tda7x6);
assign Tda7x6 = (!Gaa7x6);
assign Tdvxx6 = (~(Rivxx6 & Vt2et6));
assign Rivxx6 = (Bqoxx6 & Xgmov6);
assign Jbmxx6 = (Zivxx6 & Hjvxx6);
assign Hjvxx6 = (Pjvxx6 & Xjvxx6);
assign Xjvxx6 = (~(Fkvxx6 & Nkvxx6));
assign Fkvxx6 = (Av77x6 & Hp67x6);
assign Pjvxx6 = (~(Vkvxx6 & Nkvxx6));
assign Vkvxx6 = (Dca7x6 & Dh57x6);
assign Zivxx6 = (Dlvxx6 & Llvxx6);
assign Llvxx6 = (~(Tlvxx6 & Nkvxx6));
assign Tlvxx6 = (H287x6 & Rh57x6);
assign Dlvxx6 = (~(Bmvxx6 & Nkvxx6));
assign Nkvxx6 = (Vt2et6 & Eylxx6);
assign Bmvxx6 = (Gaa7x6 & Kn67x6);
assign U9jxx6 = (Thuxx6 & Lhuxx6);
assign Lhuxx6 = (Hyhhw6 & Jmvxx6);
assign Jmvxx6 = (~(Rmvxx6 & Zmvxx6));
assign Zmvxx6 = (Hnvxx6 & Pnvxx6);
assign Pnvxx6 = (Fiihw6 & Vkhhw6);
assign Hnvxx6 = (B3hhw6 & Vjihw6);
assign Vjihw6 = (~(Ggoov6 & Mpihw6));
assign B3hhw6 = (~(Xnvxx6 & Dioov6));
assign Xnvxx6 = (Dwb7z6[5] & Aqihw6);
assign Rmvxx6 = (Lmhhw6 & Fovxx6);
assign Fovxx6 = (Hkhhw6 & Novxx6);
assign Novxx6 = (~(Clhhw6 & Vovxx6));
assign Hkhhw6 = (Dpvxx6 & Lpvxx6);
assign Lpvxx6 = (I1d7x6 & U3a7x6);
assign Dpvxx6 = (K2d7x6 & Iqmov6);
assign K2d7x6 = (Tpvxx6 | Bqvxx6);
assign Lmhhw6 = (~(Jqvxx6 | Jkihw6));
assign Jkihw6 = (!G9hhw6);
assign G9hhw6 = (Rqvxx6 & Zqvxx6);
assign Zqvxx6 = (Hrvxx6 & Prvxx6);
assign Prvxx6 = (Kb9iw6 & I3wnv6);
assign I3wnv6 = (!Atmov6);
assign Hrvxx6 = (Xrvxx6 & Mq9iw6);
assign Xrvxx6 = (~(Rb9iw6 & Dwb7z6[1]));
assign Rqvxx6 = (Fsvxx6 & Nsvxx6);
assign Fsvxx6 = (Vsvxx6 & Dtvxx6);
assign Dtvxx6 = (~(Ltvxx6 & Luvnv6));
assign Vsvxx6 = (~(Ttvxx6 & Bhoov6));
assign Ttvxx6 = (Nvvnv6 & Buvxx6);
assign Jqvxx6 = (~(Juvxx6 & Ruvxx6));
assign Juvxx6 = (~(Tnzdt6 & Zuvxx6));
assign Zuvxx6 = (~(Hvvxx6 & Pvvxx6));
assign Pvvxx6 = (~(S0bov6 | Q0hhw6));
assign S0bov6 = (!Rhphw6);
assign Hvvxx6 = (Xvvxx6 & Fwvxx6);
assign Thuxx6 = (Nwvxx6 & Vwvxx6);
assign Vwvxx6 = (Hcihw6 & Dxvxx6);
assign Dxvxx6 = (Pvuxx6 ^ Qdihw6);
assign Pvuxx6 = (!Bjfhw6);
assign Bjfhw6 = (~(Lxvxx6 & Txvxx6));
assign Txvxx6 = (Byvxx6 & Jyvxx6);
assign Jyvxx6 = (~(Ryvxx6 & Oac7z6[2]));
assign Byvxx6 = (~(X3vxx6 & Rrfhw6));
assign Lxvxx6 = (Zyvxx6 & Hzvxx6);
assign Hzvxx6 = (~(Pzvxx6 & Xzvxx6));
assign Xzvxx6 = (~(F0wxx6 & N0wxx6));
assign N0wxx6 = (V0wxx6 & D1wxx6);
assign D1wxx6 = (~(G3nov6 & L1wxx6));
assign G3nov6 = (~(T1wxx6 & B2wxx6));
assign T1wxx6 = (J2wxx6 & R2wxx6);
assign R2wxx6 = (~(Z2wxx6 & H3wxx6));
assign H3wxx6 = (~(P3wxx6 | X3wxx6));
assign Z2wxx6 = (F4wxx6 & N4wxx6);
assign V0wxx6 = (V4wxx6 & D5wxx6);
assign D5wxx6 = (~(L5wxx6 & Kpaov6));
assign V4wxx6 = (~(Ntg7z6[2] & T5wxx6));
assign F0wxx6 = (B6wxx6 & J6wxx6);
assign B6wxx6 = (R6wxx6 & Z6wxx6);
assign Z6wxx6 = (~(H7wxx6 & Qij7z6[2]));
assign R6wxx6 = (~(U2wnv6 & Pxg7z6[2]));
assign Zyvxx6 = (~(P7wxx6 & Xwe7z6[2]));
assign Hcihw6 = (X7wxx6 & Qg2nv6);
assign Nwvxx6 = (F8wxx6 & N8wxx6);
assign N8wxx6 = (~(Ijfhw6 ^ Vcihw6));
assign Ijfhw6 = (!Vrjxx6);
assign Vrjxx6 = (V8wxx6 & D9wxx6);
assign D9wxx6 = (L9wxx6 & T9wxx6);
assign T9wxx6 = (~(Pzvxx6 & Bawxx6));
assign Bawxx6 = (~(Jawxx6 & Rawxx6));
assign Rawxx6 = (Zawxx6 & Hbwxx6);
assign Hbwxx6 = (Pbwxx6 & Eminv6);
assign Pbwxx6 = (~(Xbwxx6 & Ckihw6));
assign Xbwxx6 = (Cwlnv6 & Fcwxx6);
assign Fcwxx6 = (~(Xkr8v6 & Ncwxx6));
assign Ncwxx6 = (~(Xdphw6 & H7nov6));
assign Zawxx6 = (Vcwxx6 & Ddwxx6);
assign Ddwxx6 = (~(Ldwxx6 & H7wxx6));
assign Ldwxx6 = (Qij7z6[1] & Tdwxx6);
assign Vcwxx6 = (~(Bewxx6 & Lxydt6));
assign Bewxx6 = (~(Jewxx6 & Rewxx6));
assign Rewxx6 = (~(Zewxx6 & Q0wnv6));
assign Zewxx6 = (Clhhw6 & H7nov6);
assign H7nov6 = (~(Hfwxx6 & Pfwxx6));
assign Pfwxx6 = (Xfwxx6 & Fgwxx6);
assign Fgwxx6 = (~(Ngwxx6 & Vgwxx6));
assign Ngwxx6 = (~(Dhwxx6 | Lhwxx6));
assign Xfwxx6 = (Thwxx6 & Biwxx6);
assign Thwxx6 = (~(Jiwxx6 & Riwxx6));
assign Riwxx6 = (Ziwxx6 & Hjwxx6);
assign Jiwxx6 = (Pjwxx6 & Xjwxx6);
assign Hfwxx6 = (B2wxx6 & Fkwxx6);
assign Fkwxx6 = (~(F4wxx6 & Nkwxx6));
assign Nkwxx6 = (~(Vkwxx6 & N4wxx6));
assign B2wxx6 = (Dlwxx6 & Llwxx6);
assign Llwxx6 = (~(Xjwxx6 & Tlwxx6));
assign Jewxx6 = (~(Ntg7z6[1] & Ot97x6));
assign Jawxx6 = (Bmwxx6 & Jmwxx6);
assign Jmwxx6 = (~(Rmwxx6 & Dwb7z6[5]));
assign Bmwxx6 = (Zmwxx6 & Hnwxx6);
assign Hnwxx6 = (~(Pnwxx6 & Qg2nv6));
assign Pnwxx6 = (~(Xnwxx6 & Fowxx6));
assign Fowxx6 = (Nowxx6 & Vowxx6);
assign Vowxx6 = (~(Ntg7z6[1] & Tka7x6));
assign Nowxx6 = (Xma7x6 & Rhphw6);
assign Rhphw6 = (~(Dpwxx6 & Dioov6));
assign Dpwxx6 = (Lpwxx6 & Luvnv6);
assign Xnwxx6 = (Tpwxx6 & Bqwxx6);
assign Bqwxx6 = (~(Ywaov6 & Vqihw6));
assign Tpwxx6 = (~(U2wnv6 & Pxg7z6[1]));
assign Zmwxx6 = (~(Rioov6 & Xumov6));
assign L9wxx6 = (~(P7wxx6 & Xwe7z6[1]));
assign V8wxx6 = (Jqwxx6 & Rqwxx6);
assign Rqwxx6 = (~(X3vxx6 & Sofhw6));
assign Jqwxx6 = (~(Ryvxx6 & Oac7z6[1]));
assign F8wxx6 = (Zqwxx6 & Hrwxx6);
assign Hrwxx6 = (Xvuxx6 ^ Seihw6);
assign Xvuxx6 = (!Xgfhw6);
assign Xgfhw6 = (~(Prwxx6 & Xrwxx6));
assign Xrwxx6 = (Fswxx6 & Nswxx6);
assign Nswxx6 = (~(Pzvxx6 & Vswxx6));
assign Vswxx6 = (~(Dtwxx6 & Ltwxx6));
assign Ltwxx6 = (Ttwxx6 & Buwxx6);
assign Buwxx6 = (~(L1wxx6 & Ixmov6));
assign Ixmov6 = (~(Juwxx6 & Ruwxx6));
assign Juwxx6 = (Zuwxx6 & Hvwxx6);
assign Hvwxx6 = (~(Pvwxx6 & Xjwxx6));
assign Pvwxx6 = (Xvwxx6 & Fwwxx6);
assign Xvwxx6 = (~(Nwwxx6 & Vwwxx6));
assign Vwwxx6 = (~(Dxwxx6 & Ziwxx6));
assign Zuwxx6 = (~(Lxwxx6 & Txwxx6));
assign Lxwxx6 = (~(Bywxx6 & Jywxx6));
assign Jywxx6 = (~(Rywxx6 & N4wxx6));
assign Rywxx6 = (~(Vkwxx6 & Zywxx6));
assign Zywxx6 = (Hzwxx6 | Pzwxx6);
assign Ttwxx6 = (Xzwxx6 & F0xxx6);
assign F0xxx6 = (~(L5wxx6 & Pxmov6));
assign Xzwxx6 = (~(Ntg7z6[0] & T5wxx6));
assign Dtwxx6 = (N0xxx6 & J6wxx6);
assign N0xxx6 = (V0xxx6 & D1xxx6);
assign D1xxx6 = (~(H7wxx6 & Qij7z6[0]));
assign V0xxx6 = (~(U2wnv6 & Pxg7z6[0]));
assign Fswxx6 = (~(Xwe7z6[0] & P7wxx6));
assign Prwxx6 = (L1xxx6 & T1xxx6);
assign T1xxx6 = (~(X3vxx6 & B2xxx6));
assign L1xxx6 = (~(Ryvxx6 & Oac7z6[0]));
assign Zqwxx6 = (Nsuxx6 ^ Gfihw6);
assign Nsuxx6 = (!Uifhw6);
assign Uifhw6 = (~(J2xxx6 & R2xxx6));
assign R2xxx6 = (Z2xxx6 & H3xxx6);
assign H3xxx6 = (~(Pzvxx6 & P3xxx6));
assign P3xxx6 = (~(X3xxx6 & F4xxx6));
assign F4xxx6 = (N4xxx6 & V4xxx6);
assign V4xxx6 = (~(H0nov6 & L1wxx6));
assign L1wxx6 = (Clhhw6 | Fpphw6);
assign H0nov6 = (~(D5xxx6 & Ruwxx6));
assign Ruwxx6 = (Dlwxx6 & Biwxx6);
assign Biwxx6 = (~(L5xxx6 & T5xxx6));
assign T5xxx6 = (!B6xxx6);
assign Dlwxx6 = (~(J6xxx6 & R6xxx6));
assign J6xxx6 = (~(Z6xxx6 | Dhwxx6));
assign D5xxx6 = (J2wxx6 & H7xxx6);
assign H7xxx6 = (~(P7xxx6 & Xjwxx6));
assign P7xxx6 = (~(Tlwxx6 | X7xxx6));
assign J2wxx6 = (~(F8xxx6 & Z6xxx6));
assign N4xxx6 = (N8xxx6 & V8xxx6);
assign V8xxx6 = (~(L5wxx6 & Xlaov6));
assign L5wxx6 = (Cwlnv6 | Rioov6);
assign N8xxx6 = (~(Ntg7z6[3] & T5wxx6));
assign X3xxx6 = (D9xxx6 & J6wxx6);
assign J6wxx6 = (L9xxx6 & T9xxx6);
assign T9xxx6 = (Baxxx6 & Jaxxx6);
assign Jaxxx6 = (~(Cwlnv6 & Raxxx6));
assign Baxxx6 = (Zaxxx6 & Hbxxx6);
assign Hbxxx6 = (~(Vxphw6 & Aga7z6));
assign Vxphw6 = (~(Vkhhw6 & Twphw6));
assign Zaxxx6 = (~(Tnzdt6 & Pbxxx6));
assign Pbxxx6 = (Tka7x6 | U2wnv6);
assign L9xxx6 = (~(Xbxxx6 | Fcxxx6));
assign Fcxxx6 = (Clhhw6 & K9d7x6);
assign Xbxxx6 = (H7wxx6 ? Qij7z6[4] : Ncxxx6);
assign Ncxxx6 = (Vcxxx6 & Ddxxx6);
assign Ddxxx6 = (Yihhw6 & L5xiw6);
assign L5xiw6 = (!U2wnv6);
assign Vcxxx6 = (Ldxxx6 & Tdxxx6);
assign Ldxxx6 = (!T5wxx6);
assign T5wxx6 = (Tka7x6 | Ot97x6);
assign D9xxx6 = (Bexxx6 & Jexxx6);
assign Jexxx6 = (~(H7wxx6 & Qij7z6[3]));
assign Bexxx6 = (~(U2wnv6 & Pxg7z6[3]));
assign Z2xxx6 = (~(P7wxx6 & Xwe7z6[3]));
assign P7wxx6 = (~(Rexxx6 | Pzvxx6));
assign Rexxx6 = (~(Zexxx6 & Hfxxx6));
assign J2xxx6 = (Pfxxx6 & Xfxxx6);
assign Xfxxx6 = (~(X3vxx6 & Omfhw6));
assign X3vxx6 = (~(Hfxxx6 | Pzvxx6));
assign Pfxxx6 = (~(Ryvxx6 & Oac7z6[3]));
assign Ryvxx6 = (~(Fgxxx6 | Zexxx6));
assign Zexxx6 = (K4aov6 | Ngxxx6);
assign Fgxxx6 = (Pzvxx6 | Bi37x6);
assign Bi37x6 = (!Hfxxx6);
assign Hfxxx6 = (~(Vgxxx6 & Dhxxx6));
assign Dhxxx6 = (~(Qg2nv6 & Lhxxx6));
assign Lhxxx6 = (~(Thxxx6 & Bitiw6));
assign Thxxx6 = (Dxtiw6 & Bixxx6);
assign Bixxx6 = (~(Jixxx6 & Rixxx6));
assign Rixxx6 = (Bdf7z6[0] ? Hjxxx6 : Zixxx6);
assign Hjxxx6 = (Pjxxx6 & Pxfov6);
assign Pjxxx6 = (~(Ghtiw6 | Bdf7z6[3]));
assign Zixxx6 = (M5aov6 & Egtiw6);
assign Egtiw6 = (!Xjxxx6);
assign Jixxx6 = (~(Zgtiw6 | G427x6));
assign Dxtiw6 = (~(Tdtiw6 & Ehgdt6));
assign Vgxxx6 = (~(Yxtiw6 & Mrnov6));
assign Pzvxx6 = (~(Fkxxx6 & Nkxxx6));
assign Nkxxx6 = (Wi37x6 & Wb37x6);
assign Wb37x6 = (~(Raxxx6 & Vkxxx6));
assign Vkxxx6 = (~(Dlxxx6 & Llxxx6));
assign Llxxx6 = (Tlxxx6 & Bmxxx6);
assign Bmxxx6 = (C7jxx6 | Jmxxx6);
assign Tlxxx6 = (Rmxxx6 & Zmxxx6);
assign Zmxxx6 = (~(Nvvnv6 & Hnxxx6));
assign Hnxxx6 = (~(Pnxxx6 & Xnxxx6));
assign Xnxxx6 = (~(Dwb7z6[0] & Sna7x6));
assign Rmxxx6 = (~(Xfa7x6 & Foxxx6));
assign Foxxx6 = (~(Noxxx6 & Voxxx6));
assign Voxxx6 = (~(Doihw6 & Aqihw6));
assign Noxxx6 = (~(Bhoov6 & Bqvxx6));
assign Dlxxx6 = (Dpxxx6 & Lpxxx6);
assign Lpxxx6 = (Dwb7z6[1] ? Bqxxx6 : Tpxxx6);
assign Bqxxx6 = (~(Lpwxx6 & Dwb7z6[3]));
assign Dpxxx6 = (Jqxxx6 & Rqxxx6);
assign Rqxxx6 = (~(Rb9iw6 & Aqihw6));
assign Wi37x6 = (Zqxxx6 & Hrxxx6);
assign Hrxxx6 = (~(Prxxx6 & Xrxxx6));
assign Xrxxx6 = (~(Qij7z6[6] | X4eet6));
assign Prxxx6 = (~(Fsxxx6 | Qij7z6[5]));
assign Zqxxx6 = (~(Rmwxx6 & Lpwxx6));
assign Fkxxx6 = (Dj37x6 & Ib37x6);
assign Ib37x6 = (Nsxxx6 & Vsxxx6);
assign Vsxxx6 = (Dtxxx6 & Ltxxx6);
assign Ltxxx6 = (~(Ttxxx6 & Vglhw6));
assign Ttxxx6 = (~(Qg2nv6 & Buxxx6));
assign Dtxxx6 = (Juxxx6 & Xma7x6);
assign Xma7x6 = (~(Ruxxx6 & Fxaov6));
assign Juxxx6 = (~(Zuxxx6 & Dioov6));
assign Zuxxx6 = (Fxaov6 & Lpwxx6);
assign Nsxxx6 = (Hvxxx6 & Qlinv6);
assign Qlinv6 = (Pvxxx6 & C0b7x6);
assign C0b7x6 = (Gha7x6 | Xvxxx6);
assign Pvxxx6 = (~(Rmwxx6 & Bhoov6));
assign Hvxxx6 = (Fwxxx6 & Nwxxx6);
assign Nwxxx6 = (~(Vwxxx6 & Aga7z6));
assign Vwxxx6 = (~(Dxxxx6 & Tdxxx6));
assign Dxxxx6 = (I1d7x6 & Tpvxx6);
assign Fwxxx6 = (~(L9nov6 & K9d7x6));
assign Dj37x6 = (Lxxxx6 & Txxxx6);
assign Txxxx6 = (~(Ii9ov6 & Byxxx6));
assign Byxxx6 = (Jyxxx6 | Dur7x6);
assign Jyxxx6 = (Hjihw6 & L9nov6);
assign L9nov6 = (!Tdxxx6);
assign Lxxxx6 = (~(Ryxxx6 | Eyknv6));
assign Ryxxx6 = (!Zyxxx6);
assign L5vxx6 = (~(S8jxx6 & Cmm7z6[31]));
assign S8jxx6 = (Hyhhw6 & Hzxxx6);
assign Hzxxx6 = (~(Pzxxx6 & Xzxxx6));
assign Xzxxx6 = (F0yxx6 & N0yxx6);
assign N0yxx6 = (~(Lsphw6 & Clhhw6));
assign F0yxx6 = (V0yxx6 & Qsaov6);
assign V0yxx6 = (~(D1yxx6 & Qg2nv6));
assign D1yxx6 = (Q0hhw6 | D4hhw6);
assign D4hhw6 = (!Fwvxx6);
assign Pzxxx6 = (Wvhhw6 & C8nov6);
assign C8nov6 = (L1yxx6 & T1yxx6);
assign L1yxx6 = (~(Dihhw6 | B2yxx6));
assign Wvhhw6 = (J2yxx6 & R2yxx6);
assign R2yxx6 = (Qxknv6 & Z2yxx6);
assign J2yxx6 = (H3yxx6 & G3a7x6);
assign H3yxx6 = (Xvvxx6 | Tnzdt6);
assign Xvvxx6 = (P3yxx6 & X3yxx6);
assign Hyhhw6 = (!Zs4ov6);
assign Zs4ov6 = (~(Yfadt6 & F4yxx6));
assign F4yxx6 = (~(N4yxx6 & V4yxx6));
assign V4yxx6 = (D5yxx6 & L5yxx6);
assign L5yxx6 = (T5yxx6 & Fwvxx6);
assign Fwvxx6 = (~(B6yxx6 & Xfa7x6));
assign B6yxx6 = (Doihw6 & Fxaov6);
assign T5yxx6 = (~(J6yxx6 & Bhoov6));
assign J6yxx6 = (Vqihw6 & R6yxx6);
assign R6yxx6 = (~(Zna7x6 & Z6yxx6));
assign Z6yxx6 = (~(Tnzdt6 & Dwb7z6[3]));
assign D5yxx6 = (H7yxx6 & P7yxx6);
assign P7yxx6 = (~(D3jnv6 & X7yxx6));
assign D3jnv6 = (O5a7z6 & Aga7z6);
assign H7yxx6 = (~(Tnzdt6 & F8yxx6));
assign F8yxx6 = (~(Mq9iw6 & N8yxx6));
assign N8yxx6 = (~(Rb9iw6 & Fxaov6));
assign Mq9iw6 = (~(V8yxx6 & Fulnv6));
assign V8yxx6 = (Lpwxx6 & Nvvnv6);
assign N4yxx6 = (D9yxx6 & L9yxx6);
assign L9yxx6 = (T9yxx6 & Bayxx6);
assign Bayxx6 = (~(Q0hhw6 & Jayxx6));
assign Jayxx6 = (~(Qg2nv6 & Rayxx6));
assign Rayxx6 = (~(Noa7x6 & Zayxx6));
assign T9yxx6 = (~(Gr2et6 & Hbyxx6));
assign Hbyxx6 = (~(Pbyxx6 & Xbyxx6));
assign Xbyxx6 = (Fcyxx6 & Ncyxx6);
assign Ncyxx6 = (Vcyxx6 & Srknv6);
assign Fcyxx6 = (Ddyxx6 & Ldyxx6);
assign Ldyxx6 = (~(Lpwxx6 & Tdyxx6));
assign Tdyxx6 = (~(Bwvnv6 & Zna7x6));
assign Ddyxx6 = (~(Beyxx6 & Mpihw6));
assign Pbyxx6 = (Jeyxx6 & Reyxx6);
assign Reyxx6 = (P3yxx6 | Olzdt6);
assign Olzdt6 = (Iga7z6 & Qg2nv6);
assign Jeyxx6 = (Kur7x6 & Zeyxx6);
assign Zeyxx6 = (G3a7x6 | Aiadt6);
assign Kur7x6 = (~(Clhhw6 & Hjihw6));
assign D9yxx6 = (Zwehw6 & Hfyxx6);
assign Hfyxx6 = (~(Pfyxx6 & Raxxx6));
assign Raxxx6 = (!Ckihw6);
assign Pfyxx6 = (~(Xfyxx6 & Fgyxx6));
assign Fgyxx6 = (Ngyxx6 & Nsvxx6);
assign Nsvxx6 = (Vgyxx6 & Jqxxx6);
assign Jqxxx6 = (Dhyxx6 & Gpmov6);
assign Vgyxx6 = (Lhyxx6 & Thyxx6);
assign Thyxx6 = (~(Biyxx6 & Bhoov6));
assign Biyxx6 = (Xfa7x6 & Xvxxx6);
assign Lhyxx6 = (~(Ruxxx6 & Mpihw6));
assign Ngyxx6 = (Jiyxx6 & N3a7x6);
assign Jiyxx6 = (Sga7x6 | Jmxxx6);
assign Jmxxx6 = (Riyxx6 & Ziyxx6);
assign Ziyxx6 = (~(Lpwxx6 & Kioov6));
assign Riyxx6 = (~(Bhoov6 & Mpihw6));
assign Xfyxx6 = (~(Hjyxx6 | Pjyxx6));
assign Pjyxx6 = (Fkyxx6 ? Rb9iw6 : Xjyxx6);
assign Xjyxx6 = (Bhoov6 & Nvvnv6);
assign Hjyxx6 = (Kioov6 ? Ggoov6 : Ltvxx6);
assign Zwehw6 = (Esihw6 & U1ihw6);
assign U1ihw6 = (!Kxvnv6);
assign Kxvnv6 = (N3onv6 & Nkyxx6);
assign Esihw6 = (!Irriw6);
assign Irriw6 = (S0ihw6 | Mqhhw6);
assign Mqhhw6 = (N3onv6 & Vkyxx6);
assign S0ihw6 = (Yqvnv6 | Wwvnv6);
assign Wwvnv6 = (Dlyxx6 & N3onv6);
assign Dlyxx6 = (Ryfhw6 & Llyxx6);
assign Yqvnv6 = (N3onv6 & Tlyxx6);
assign I4s7v6 = (~(Bmyxx6 & Jmyxx6));
assign Jmyxx6 = (~(L8wnv6 & Itb7z6[27]));
assign Bmyxx6 = (Rmyxx6 & Zmyxx6);
assign Zmyxx6 = (~(G9wnv6 & Hnyxx6));
assign Hnyxx6 = (~(Pnyxx6 & Xnyxx6));
assign Xnyxx6 = (Foyxx6 & Noyxx6);
assign Noyxx6 = (Wawnv6 | Voyxx6);
assign Foyxx6 = (~(Dtm7z6[3] & Dpyxx6));
assign Pnyxx6 = (Lpyxx6 & Tpyxx6);
assign Tpyxx6 = (~(Dtm7z6[0] & HRDATAD[27]));
assign Lpyxx6 = (~(Dtm7z6[1] & HRDATAS[27]));
assign Rmyxx6 = (~(Fcwnv6 & Mnyhw6));
assign Mnyhw6 = (JTAGNSW ? Aixmz6[27] : Ulxmz6[27]);
assign B4s7v6 = (~(Bqyxx6 & Jqyxx6));
assign Jqyxx6 = (~(L8wnv6 & Itb7z6[28]));
assign Bqyxx6 = (Rqyxx6 & Zqyxx6);
assign Zqyxx6 = (~(G9wnv6 & Hryxx6));
assign Hryxx6 = (~(Pryxx6 & Xryxx6));
assign Xryxx6 = (Fsyxx6 & Nsyxx6);
assign Nsyxx6 = (Wawnv6 | Vsyxx6);
assign Fsyxx6 = (~(Dtm7z6[3] & Dtyxx6));
assign Pryxx6 = (Ltyxx6 & Ttyxx6);
assign Ttyxx6 = (~(Dtm7z6[0] & HRDATAD[28]));
assign Ltyxx6 = (~(Dtm7z6[1] & HRDATAS[28]));
assign Rqyxx6 = (~(Fcwnv6 & Lqyhw6));
assign Lqyhw6 = (JTAGNSW ? Aixmz6[28] : Ulxmz6[28]);
assign U3s7v6 = (~(Buyxx6 & Juyxx6));
assign Juyxx6 = (~(Gsexx6 & Ruyxx6));
assign Ruyxx6 = (~(Zuyxx6 & Hvyxx6));
assign Hvyxx6 = (Pvyxx6 & Xvyxx6);
assign Xvyxx6 = (Fwyxx6 & Nwyxx6);
assign Nwyxx6 = (Vwyxx6 & Dxyxx6);
assign Dxyxx6 = (~(Yuexx6 & Bq0nz6[7]));
assign Vwyxx6 = (Lxyxx6 & Txyxx6);
assign Txyxx6 = (~(Tvexx6 & Fl0nz6[7]));
assign Lxyxx6 = (~(Awexx6 & Jg0nz6[7]));
assign Fwyxx6 = (Byyxx6 & Jyyxx6);
assign Jyyxx6 = (~(Vwexx6 & Nb0nz6[7]));
assign Byyxx6 = (Ryyxx6 & Zyyxx6);
assign Zyyxx6 = (~(Qxexx6 & R60nz6[7]));
assign Ryyxx6 = (~(Xxexx6 & V10nz6[7]));
assign Pvyxx6 = (Hzyxx6 & Pzyxx6);
assign Pzyxx6 = (Xzyxx6 & F0zxx6);
assign F0zxx6 = (~(Gzexx6 & Zwzmz6[7]));
assign Xzyxx6 = (N0zxx6 & V0zxx6);
assign V0zxx6 = (~(B0fxx6 & Dszmz6[7]));
assign N0zxx6 = (~(I0fxx6 & Lo0nz6[7]));
assign Hzyxx6 = (D1zxx6 & L1zxx6);
assign L1zxx6 = (~(D1fxx6 & Pj0nz6[7]));
assign D1zxx6 = (T1zxx6 & B2zxx6);
assign B2zxx6 = (~(Y1fxx6 & Te0nz6[7]));
assign T1zxx6 = (~(F2fxx6 & X90nz6[7]));
assign Zuyxx6 = (J2zxx6 & R2zxx6);
assign R2zxx6 = (Z2zxx6 & H3zxx6);
assign H3zxx6 = (P3zxx6 & X3zxx6);
assign X3zxx6 = (~(C4fxx6 & B50nz6[7]));
assign P3zxx6 = (F4zxx6 & N4zxx6);
assign N4zxx6 = (~(X4fxx6 & F00nz6[7]));
assign F4zxx6 = (~(E5fxx6 & Jvzmz6[7]));
assign Z2zxx6 = (V4zxx6 & D5zxx6);
assign D5zxx6 = (~(Z5fxx6 & Nqzmz6[7]));
assign V4zxx6 = (L5zxx6 & T5zxx6);
assign T5zxx6 = (~(U6fxx6 & Vm0nz6[7]));
assign L5zxx6 = (~(B7fxx6 & Zh0nz6[7]));
assign J2zxx6 = (B6zxx6 & J6zxx6);
assign J6zxx6 = (R6zxx6 & Z6zxx6);
assign Z6zxx6 = (~(K8fxx6 & Dd0nz6[7]));
assign R6zxx6 = (H7zxx6 & P7zxx6);
assign P7zxx6 = (~(F9fxx6 & H80nz6[7]));
assign H7zxx6 = (~(M9fxx6 & L30nz6[7]));
assign B6zxx6 = (X7zxx6 & F8zxx6);
assign F8zxx6 = (~(Xozmz6[7] & Hafxx6));
assign X7zxx6 = (N8zxx6 & V8zxx6);
assign V8zxx6 = (~(Cbfxx6 & Ttzmz6[7]));
assign N8zxx6 = (~(Jbfxx6 & Pyzmz6[7]));
assign Buyxx6 = (Gs5ov6 ? L9zxx6 : D9zxx6);
assign L9zxx6 = (~(T9zxx6 & Bazxx6));
assign Bazxx6 = (~(Uu0nz6[0] | Uu0nz6[2]));
assign T9zxx6 = (~(Jazxx6 | At67v6));
assign D9zxx6 = (!Sj67z6);
assign N3s7v6 = (~(Razxx6 & Zazxx6));
assign Zazxx6 = (~(Gsexx6 & Hbzxx6));
assign Hbzxx6 = (~(Pbzxx6 & Xbzxx6));
assign Xbzxx6 = (Fczxx6 & Nczxx6);
assign Nczxx6 = (Vczxx6 & Ddzxx6);
assign Ddzxx6 = (Ldzxx6 & Tdzxx6);
assign Tdzxx6 = (~(Yuexx6 & Bq0nz6[6]));
assign Ldzxx6 = (Bezxx6 & Jezxx6);
assign Jezxx6 = (~(Tvexx6 & Fl0nz6[6]));
assign Bezxx6 = (~(Awexx6 & Jg0nz6[6]));
assign Vczxx6 = (Rezxx6 & Zezxx6);
assign Zezxx6 = (~(Vwexx6 & Nb0nz6[6]));
assign Rezxx6 = (Hfzxx6 & Pfzxx6);
assign Pfzxx6 = (~(Qxexx6 & R60nz6[6]));
assign Hfzxx6 = (~(Xxexx6 & V10nz6[6]));
assign Fczxx6 = (Xfzxx6 & Fgzxx6);
assign Fgzxx6 = (Ngzxx6 & Vgzxx6);
assign Vgzxx6 = (~(Gzexx6 & Zwzmz6[6]));
assign Ngzxx6 = (Dhzxx6 & Lhzxx6);
assign Lhzxx6 = (~(B0fxx6 & Dszmz6[6]));
assign Dhzxx6 = (~(I0fxx6 & Lo0nz6[6]));
assign Xfzxx6 = (Thzxx6 & Bizxx6);
assign Bizxx6 = (~(D1fxx6 & Pj0nz6[6]));
assign Thzxx6 = (Jizxx6 & Rizxx6);
assign Rizxx6 = (~(Y1fxx6 & Te0nz6[6]));
assign Jizxx6 = (~(F2fxx6 & X90nz6[6]));
assign Pbzxx6 = (Zizxx6 & Hjzxx6);
assign Hjzxx6 = (Pjzxx6 & Xjzxx6);
assign Xjzxx6 = (Fkzxx6 & Nkzxx6);
assign Nkzxx6 = (~(C4fxx6 & B50nz6[6]));
assign Fkzxx6 = (Vkzxx6 & Dlzxx6);
assign Dlzxx6 = (~(X4fxx6 & F00nz6[6]));
assign Vkzxx6 = (~(E5fxx6 & Jvzmz6[6]));
assign Pjzxx6 = (Llzxx6 & Tlzxx6);
assign Tlzxx6 = (~(Z5fxx6 & Nqzmz6[6]));
assign Llzxx6 = (Bmzxx6 & Jmzxx6);
assign Jmzxx6 = (~(U6fxx6 & Vm0nz6[6]));
assign Bmzxx6 = (~(B7fxx6 & Zh0nz6[6]));
assign Zizxx6 = (Rmzxx6 & Zmzxx6);
assign Zmzxx6 = (Hnzxx6 & Pnzxx6);
assign Pnzxx6 = (~(K8fxx6 & Dd0nz6[6]));
assign Hnzxx6 = (Xnzxx6 & Fozxx6);
assign Fozxx6 = (~(F9fxx6 & H80nz6[6]));
assign Xnzxx6 = (~(M9fxx6 & L30nz6[6]));
assign Rmzxx6 = (Nozxx6 & Vozxx6);
assign Vozxx6 = (~(Xozmz6[6] & Hafxx6));
assign Nozxx6 = (Dpzxx6 & Lpzxx6);
assign Lpzxx6 = (~(Cbfxx6 & Ttzmz6[6]));
assign Dpzxx6 = (~(Jbfxx6 & Pyzmz6[6]));
assign Razxx6 = (~(Kj67z6 & Lr5ov6));
assign G3s7v6 = (~(Tpzxx6 & Bqzxx6));
assign Bqzxx6 = (~(Gsexx6 & Jqzxx6));
assign Jqzxx6 = (~(Rqzxx6 & Zqzxx6));
assign Zqzxx6 = (Hrzxx6 & Przxx6);
assign Przxx6 = (Xrzxx6 & Fszxx6);
assign Fszxx6 = (Nszxx6 & Vszxx6);
assign Vszxx6 = (~(Yuexx6 & Bq0nz6[5]));
assign Nszxx6 = (Dtzxx6 & Ltzxx6);
assign Ltzxx6 = (~(Tvexx6 & Fl0nz6[5]));
assign Dtzxx6 = (~(Awexx6 & Jg0nz6[5]));
assign Xrzxx6 = (Ttzxx6 & Buzxx6);
assign Buzxx6 = (~(Vwexx6 & Nb0nz6[5]));
assign Ttzxx6 = (Juzxx6 & Ruzxx6);
assign Ruzxx6 = (~(Qxexx6 & R60nz6[5]));
assign Juzxx6 = (~(Xxexx6 & V10nz6[5]));
assign Hrzxx6 = (Zuzxx6 & Hvzxx6);
assign Hvzxx6 = (Pvzxx6 & Xvzxx6);
assign Xvzxx6 = (~(Gzexx6 & Zwzmz6[5]));
assign Pvzxx6 = (Fwzxx6 & Nwzxx6);
assign Nwzxx6 = (~(B0fxx6 & Dszmz6[5]));
assign Fwzxx6 = (~(I0fxx6 & Lo0nz6[5]));
assign Zuzxx6 = (Vwzxx6 & Dxzxx6);
assign Dxzxx6 = (~(D1fxx6 & Pj0nz6[5]));
assign Vwzxx6 = (Lxzxx6 & Txzxx6);
assign Txzxx6 = (~(Y1fxx6 & Te0nz6[5]));
assign Lxzxx6 = (~(F2fxx6 & X90nz6[5]));
assign Rqzxx6 = (Byzxx6 & Jyzxx6);
assign Jyzxx6 = (Ryzxx6 & Zyzxx6);
assign Zyzxx6 = (Hzzxx6 & Pzzxx6);
assign Pzzxx6 = (~(C4fxx6 & B50nz6[5]));
assign Hzzxx6 = (Xzzxx6 & F00yx6);
assign F00yx6 = (~(X4fxx6 & F00nz6[5]));
assign Xzzxx6 = (~(E5fxx6 & Jvzmz6[5]));
assign Ryzxx6 = (N00yx6 & V00yx6);
assign V00yx6 = (~(Z5fxx6 & Nqzmz6[5]));
assign N00yx6 = (D10yx6 & L10yx6);
assign L10yx6 = (~(U6fxx6 & Vm0nz6[5]));
assign D10yx6 = (~(B7fxx6 & Zh0nz6[5]));
assign Byzxx6 = (T10yx6 & B20yx6);
assign B20yx6 = (J20yx6 & R20yx6);
assign R20yx6 = (~(K8fxx6 & Dd0nz6[5]));
assign J20yx6 = (Z20yx6 & H30yx6);
assign H30yx6 = (~(F9fxx6 & H80nz6[5]));
assign Z20yx6 = (~(M9fxx6 & L30nz6[5]));
assign T10yx6 = (P30yx6 & X30yx6);
assign X30yx6 = (~(Xozmz6[5] & Hafxx6));
assign P30yx6 = (F40yx6 & N40yx6);
assign N40yx6 = (~(Cbfxx6 & Ttzmz6[5]));
assign F40yx6 = (~(Jbfxx6 & Pyzmz6[5]));
assign Tpzxx6 = (~(Cj67z6 & Lr5ov6));
assign Z2s7v6 = (~(V40yx6 & D50yx6));
assign D50yx6 = (~(Gsexx6 & L50yx6));
assign L50yx6 = (~(T50yx6 & B60yx6));
assign B60yx6 = (J60yx6 & R60yx6);
assign R60yx6 = (Z60yx6 & H70yx6);
assign H70yx6 = (P70yx6 & X70yx6);
assign X70yx6 = (~(Yuexx6 & Bq0nz6[4]));
assign P70yx6 = (F80yx6 & N80yx6);
assign N80yx6 = (~(Tvexx6 & Fl0nz6[4]));
assign F80yx6 = (~(Awexx6 & Jg0nz6[4]));
assign Z60yx6 = (V80yx6 & D90yx6);
assign D90yx6 = (~(Vwexx6 & Nb0nz6[4]));
assign V80yx6 = (L90yx6 & T90yx6);
assign T90yx6 = (~(Qxexx6 & R60nz6[4]));
assign L90yx6 = (~(Xxexx6 & V10nz6[4]));
assign J60yx6 = (Ba0yx6 & Ja0yx6);
assign Ja0yx6 = (Ra0yx6 & Za0yx6);
assign Za0yx6 = (~(Gzexx6 & Zwzmz6[4]));
assign Ra0yx6 = (Hb0yx6 & Pb0yx6);
assign Pb0yx6 = (~(B0fxx6 & Dszmz6[4]));
assign Hb0yx6 = (~(I0fxx6 & Lo0nz6[4]));
assign Ba0yx6 = (Xb0yx6 & Fc0yx6);
assign Fc0yx6 = (~(D1fxx6 & Pj0nz6[4]));
assign Xb0yx6 = (Nc0yx6 & Vc0yx6);
assign Vc0yx6 = (~(Y1fxx6 & Te0nz6[4]));
assign Nc0yx6 = (~(F2fxx6 & X90nz6[4]));
assign T50yx6 = (Dd0yx6 & Ld0yx6);
assign Ld0yx6 = (Td0yx6 & Be0yx6);
assign Be0yx6 = (Je0yx6 & Re0yx6);
assign Re0yx6 = (~(C4fxx6 & B50nz6[4]));
assign Je0yx6 = (Ze0yx6 & Hf0yx6);
assign Hf0yx6 = (~(X4fxx6 & F00nz6[4]));
assign Ze0yx6 = (~(E5fxx6 & Jvzmz6[4]));
assign Td0yx6 = (Pf0yx6 & Xf0yx6);
assign Xf0yx6 = (~(Z5fxx6 & Nqzmz6[4]));
assign Pf0yx6 = (Fg0yx6 & Ng0yx6);
assign Ng0yx6 = (~(U6fxx6 & Vm0nz6[4]));
assign Fg0yx6 = (~(B7fxx6 & Zh0nz6[4]));
assign Dd0yx6 = (Vg0yx6 & Dh0yx6);
assign Dh0yx6 = (Lh0yx6 & Th0yx6);
assign Th0yx6 = (~(K8fxx6 & Dd0nz6[4]));
assign Lh0yx6 = (Bi0yx6 & Ji0yx6);
assign Ji0yx6 = (~(F9fxx6 & H80nz6[4]));
assign Bi0yx6 = (~(M9fxx6 & L30nz6[4]));
assign Vg0yx6 = (Ri0yx6 & Zi0yx6);
assign Zi0yx6 = (~(Xozmz6[4] & Hafxx6));
assign Ri0yx6 = (Hj0yx6 & Pj0yx6);
assign Pj0yx6 = (~(Cbfxx6 & Ttzmz6[4]));
assign Hj0yx6 = (~(Jbfxx6 & Pyzmz6[4]));
assign V40yx6 = (~(Ui67z6 & Lr5ov6));
assign S2s7v6 = (~(Xj0yx6 & Fk0yx6));
assign Fk0yx6 = (~(Mi67z6 & Lr5ov6));
assign Xj0yx6 = (Nk0yx6 & Vk0yx6);
assign Nk0yx6 = (~(Gsexx6 & Dl0yx6));
assign Dl0yx6 = (~(Ll0yx6 & Tl0yx6));
assign Tl0yx6 = (Bm0yx6 & Jm0yx6);
assign Jm0yx6 = (Rm0yx6 & Zm0yx6);
assign Zm0yx6 = (Hn0yx6 & Pn0yx6);
assign Pn0yx6 = (~(Yuexx6 & Bq0nz6[3]));
assign Hn0yx6 = (Xn0yx6 & Fo0yx6);
assign Fo0yx6 = (~(Tvexx6 & Fl0nz6[3]));
assign Xn0yx6 = (~(Awexx6 & Jg0nz6[3]));
assign Rm0yx6 = (No0yx6 & Vo0yx6);
assign Vo0yx6 = (~(Vwexx6 & Nb0nz6[3]));
assign No0yx6 = (Dp0yx6 & Lp0yx6);
assign Lp0yx6 = (~(Qxexx6 & R60nz6[3]));
assign Dp0yx6 = (~(Xxexx6 & V10nz6[3]));
assign Bm0yx6 = (Tp0yx6 & Bq0yx6);
assign Bq0yx6 = (Jq0yx6 & Rq0yx6);
assign Rq0yx6 = (~(Gzexx6 & Zwzmz6[3]));
assign Jq0yx6 = (Zq0yx6 & Hr0yx6);
assign Hr0yx6 = (~(B0fxx6 & Dszmz6[3]));
assign Zq0yx6 = (~(I0fxx6 & Lo0nz6[3]));
assign Tp0yx6 = (Pr0yx6 & Xr0yx6);
assign Xr0yx6 = (~(D1fxx6 & Pj0nz6[3]));
assign Pr0yx6 = (Fs0yx6 & Ns0yx6);
assign Ns0yx6 = (~(Y1fxx6 & Te0nz6[3]));
assign Fs0yx6 = (~(F2fxx6 & X90nz6[3]));
assign Ll0yx6 = (Vs0yx6 & Dt0yx6);
assign Dt0yx6 = (Lt0yx6 & Tt0yx6);
assign Tt0yx6 = (Bu0yx6 & Ju0yx6);
assign Ju0yx6 = (~(C4fxx6 & B50nz6[3]));
assign Bu0yx6 = (Ru0yx6 & Zu0yx6);
assign Zu0yx6 = (~(X4fxx6 & F00nz6[3]));
assign Ru0yx6 = (~(E5fxx6 & Jvzmz6[3]));
assign Lt0yx6 = (Hv0yx6 & Pv0yx6);
assign Pv0yx6 = (~(Z5fxx6 & Nqzmz6[3]));
assign Hv0yx6 = (Xv0yx6 & Fw0yx6);
assign Fw0yx6 = (~(U6fxx6 & Vm0nz6[3]));
assign Xv0yx6 = (~(B7fxx6 & Zh0nz6[3]));
assign Vs0yx6 = (Nw0yx6 & Vw0yx6);
assign Vw0yx6 = (Dx0yx6 & Lx0yx6);
assign Lx0yx6 = (~(K8fxx6 & Dd0nz6[3]));
assign Dx0yx6 = (Tx0yx6 & By0yx6);
assign By0yx6 = (~(F9fxx6 & H80nz6[3]));
assign Tx0yx6 = (~(M9fxx6 & L30nz6[3]));
assign Nw0yx6 = (Jy0yx6 & Ry0yx6);
assign Ry0yx6 = (~(Xozmz6[3] & Hafxx6));
assign Jy0yx6 = (Zy0yx6 & Hz0yx6);
assign Hz0yx6 = (~(Cbfxx6 & Ttzmz6[3]));
assign Zy0yx6 = (~(Jbfxx6 & Pyzmz6[3]));
assign L2s7v6 = (~(Pz0yx6 & Xz0yx6));
assign Xz0yx6 = (~(Ei67z6 & Lr5ov6));
assign Pz0yx6 = (F01yx6 & Vk0yx6);
assign Vk0yx6 = (~(N01yx6 & V01yx6));
assign N01yx6 = (!D11yx6);
assign F01yx6 = (~(Gsexx6 & L11yx6));
assign L11yx6 = (~(T11yx6 & B21yx6));
assign B21yx6 = (J21yx6 & R21yx6);
assign R21yx6 = (Z21yx6 & H31yx6);
assign H31yx6 = (P31yx6 & X31yx6);
assign X31yx6 = (~(Yuexx6 & Bq0nz6[2]));
assign P31yx6 = (F41yx6 & N41yx6);
assign N41yx6 = (~(Tvexx6 & Fl0nz6[2]));
assign F41yx6 = (~(Awexx6 & Jg0nz6[2]));
assign Z21yx6 = (V41yx6 & D51yx6);
assign D51yx6 = (~(Vwexx6 & Nb0nz6[2]));
assign V41yx6 = (L51yx6 & T51yx6);
assign T51yx6 = (~(Qxexx6 & R60nz6[2]));
assign L51yx6 = (~(Xxexx6 & V10nz6[2]));
assign J21yx6 = (B61yx6 & J61yx6);
assign J61yx6 = (R61yx6 & Z61yx6);
assign Z61yx6 = (~(Gzexx6 & Zwzmz6[2]));
assign R61yx6 = (H71yx6 & P71yx6);
assign P71yx6 = (~(B0fxx6 & Dszmz6[2]));
assign H71yx6 = (~(I0fxx6 & Lo0nz6[2]));
assign B61yx6 = (X71yx6 & F81yx6);
assign F81yx6 = (~(D1fxx6 & Pj0nz6[2]));
assign X71yx6 = (N81yx6 & V81yx6);
assign V81yx6 = (~(Y1fxx6 & Te0nz6[2]));
assign N81yx6 = (~(F2fxx6 & X90nz6[2]));
assign T11yx6 = (D91yx6 & L91yx6);
assign L91yx6 = (T91yx6 & Ba1yx6);
assign Ba1yx6 = (Ja1yx6 & Ra1yx6);
assign Ra1yx6 = (~(C4fxx6 & B50nz6[2]));
assign Ja1yx6 = (Za1yx6 & Hb1yx6);
assign Hb1yx6 = (~(X4fxx6 & F00nz6[2]));
assign Za1yx6 = (~(E5fxx6 & Jvzmz6[2]));
assign T91yx6 = (Pb1yx6 & Xb1yx6);
assign Xb1yx6 = (~(Z5fxx6 & Nqzmz6[2]));
assign Pb1yx6 = (Fc1yx6 & Nc1yx6);
assign Nc1yx6 = (~(U6fxx6 & Vm0nz6[2]));
assign Fc1yx6 = (~(B7fxx6 & Zh0nz6[2]));
assign D91yx6 = (Vc1yx6 & Dd1yx6);
assign Dd1yx6 = (Ld1yx6 & Td1yx6);
assign Td1yx6 = (~(K8fxx6 & Dd0nz6[2]));
assign Ld1yx6 = (Be1yx6 & Je1yx6);
assign Je1yx6 = (~(F9fxx6 & H80nz6[2]));
assign Be1yx6 = (~(M9fxx6 & L30nz6[2]));
assign Vc1yx6 = (Re1yx6 & Ze1yx6);
assign Ze1yx6 = (~(Xozmz6[2] & Hafxx6));
assign Re1yx6 = (Hf1yx6 & Pf1yx6);
assign Pf1yx6 = (~(Cbfxx6 & Ttzmz6[2]));
assign Hf1yx6 = (~(Jbfxx6 & Pyzmz6[2]));
assign E2s7v6 = (~(Xf1yx6 & Fg1yx6));
assign Fg1yx6 = (~(Gsexx6 & Ng1yx6));
assign Ng1yx6 = (~(Vg1yx6 & Dh1yx6));
assign Dh1yx6 = (Lh1yx6 & Th1yx6);
assign Th1yx6 = (Bi1yx6 & Ji1yx6);
assign Ji1yx6 = (Ri1yx6 & Zi1yx6);
assign Zi1yx6 = (~(Yuexx6 & Bq0nz6[1]));
assign Yuexx6 = (~(Hj1yx6 | Jxrnv6));
assign Ri1yx6 = (Pj1yx6 & Xj1yx6);
assign Xj1yx6 = (~(Tvexx6 & Fl0nz6[1]));
assign Tvexx6 = (~(Fk1yx6 | Jxrnv6));
assign Pj1yx6 = (~(Awexx6 & Jg0nz6[1]));
assign Awexx6 = (~(Hj1yx6 | Xxrnv6));
assign Bi1yx6 = (Nk1yx6 & Vk1yx6);
assign Vk1yx6 = (~(Vwexx6 & Nb0nz6[1]));
assign Vwexx6 = (~(Fk1yx6 | Xxrnv6));
assign Nk1yx6 = (Dl1yx6 & Ll1yx6);
assign Ll1yx6 = (~(Qxexx6 & R60nz6[1]));
assign Qxexx6 = (~(Hj1yx6 | Eyrnv6));
assign Dl1yx6 = (~(Xxexx6 & V10nz6[1]));
assign Xxexx6 = (~(Fk1yx6 | Eyrnv6));
assign Lh1yx6 = (Tl1yx6 & Bm1yx6);
assign Bm1yx6 = (Jm1yx6 & Rm1yx6);
assign Rm1yx6 = (~(Gzexx6 & Zwzmz6[1]));
assign Gzexx6 = (~(Hj1yx6 | Srcov6));
assign Hj1yx6 = (~(Zm1yx6 & Lyrnv6));
assign Jm1yx6 = (Hn1yx6 & Pn1yx6);
assign Pn1yx6 = (~(B0fxx6 & Dszmz6[1]));
assign B0fxx6 = (~(Fk1yx6 | Srcov6));
assign Fk1yx6 = (~(Zm1yx6 & E5d7v6));
assign Zm1yx6 = (Cxrnv6 & Owrnv6);
assign Hn1yx6 = (~(I0fxx6 & Lo0nz6[1]));
assign I0fxx6 = (~(Xn1yx6 | Jxrnv6));
assign Tl1yx6 = (Fo1yx6 & No1yx6);
assign No1yx6 = (~(D1fxx6 & Pj0nz6[1]));
assign D1fxx6 = (~(Vo1yx6 | Jxrnv6));
assign Fo1yx6 = (Dp1yx6 & Lp1yx6);
assign Lp1yx6 = (~(Y1fxx6 & Te0nz6[1]));
assign Y1fxx6 = (~(Xn1yx6 | Xxrnv6));
assign Dp1yx6 = (~(F2fxx6 & X90nz6[1]));
assign F2fxx6 = (~(Vo1yx6 | Xxrnv6));
assign Vg1yx6 = (Tp1yx6 & Bq1yx6);
assign Bq1yx6 = (Jq1yx6 & Rq1yx6);
assign Rq1yx6 = (Zq1yx6 & Hr1yx6);
assign Hr1yx6 = (~(C4fxx6 & B50nz6[1]));
assign C4fxx6 = (~(Xn1yx6 | Eyrnv6));
assign Zq1yx6 = (Pr1yx6 & Xr1yx6);
assign Xr1yx6 = (~(X4fxx6 & F00nz6[1]));
assign X4fxx6 = (~(Vo1yx6 | Eyrnv6));
assign Pr1yx6 = (~(E5fxx6 & Jvzmz6[1]));
assign E5fxx6 = (~(Xn1yx6 | Srcov6));
assign Xn1yx6 = (~(Fs1yx6 & Rr0nz6[0]));
assign Fs1yx6 = (Lyrnv6 & Owrnv6);
assign Jq1yx6 = (Ns1yx6 & Vs1yx6);
assign Vs1yx6 = (~(Z5fxx6 & Nqzmz6[1]));
assign Z5fxx6 = (~(Vo1yx6 | Srcov6));
assign Vo1yx6 = (~(Dt1yx6 & E5d7v6));
assign Dt1yx6 = (Rr0nz6[0] & Owrnv6);
assign Owrnv6 = (!Rr0nz6[1]);
assign Ns1yx6 = (Lt1yx6 & Tt1yx6);
assign Tt1yx6 = (~(U6fxx6 & Vm0nz6[1]));
assign U6fxx6 = (~(Bu1yx6 | Jxrnv6));
assign Lt1yx6 = (~(B7fxx6 & Zh0nz6[1]));
assign B7fxx6 = (~(Ju1yx6 | Jxrnv6));
assign Jxrnv6 = (~(Ercov6 & Qqcov6));
assign Tp1yx6 = (Ru1yx6 & Zu1yx6);
assign Zu1yx6 = (Hv1yx6 & Pv1yx6);
assign Pv1yx6 = (~(K8fxx6 & Dd0nz6[1]));
assign K8fxx6 = (~(Bu1yx6 | Xxrnv6));
assign Hv1yx6 = (Xv1yx6 & Fw1yx6);
assign Fw1yx6 = (~(F9fxx6 & H80nz6[1]));
assign F9fxx6 = (~(Xxrnv6 | Ju1yx6));
assign Xxrnv6 = (~(Hw0nz6[1] & Ercov6));
assign Xv1yx6 = (~(M9fxx6 & L30nz6[1]));
assign M9fxx6 = (~(Bu1yx6 | Eyrnv6));
assign Ru1yx6 = (Nw1yx6 & Vw1yx6);
assign Vw1yx6 = (~(Xozmz6[1] & Hafxx6));
assign Nw1yx6 = (Dx1yx6 & Lx1yx6);
assign Lx1yx6 = (~(Cbfxx6 & Ttzmz6[1]));
assign Cbfxx6 = (~(Bu1yx6 | Srcov6));
assign Bu1yx6 = (~(Tx1yx6 & Rr0nz6[1]));
assign Tx1yx6 = (Lyrnv6 & Cxrnv6);
assign Lyrnv6 = (!E5d7v6);
assign Dx1yx6 = (~(Jbfxx6 & Pyzmz6[1]));
assign Jbfxx6 = (~(Ju1yx6 | Eyrnv6));
assign Eyrnv6 = (Ercov6 | Hw0nz6[1]);
assign Gsexx6 = (V01yx6 & D11yx6);
assign V01yx6 = (By1yx6 & Gs5ov6);
assign By1yx6 = (~(H3dov6 | At67v6));
assign Xf1yx6 = (~(Wh67z6 & Lr5ov6));
assign X1s7v6 = (Ry1yx6 ? Jy1yx6 : Bv1nz6[1]);
assign Jy1yx6 = (~(Zy1yx6 & Hz1yx6));
assign Hz1yx6 = (~(Wh67z6 & Cc5ov6));
assign Q1s7v6 = (Pz1yx6 ? Ak67z6 : Au1nz6[0]);
assign J1s7v6 = (Pz1yx6 ? Sj67z6 : Au1nz6[7]);
assign C1s7v6 = (Pz1yx6 ? Kj67z6 : Au1nz6[6]);
assign V0s7v6 = (Pz1yx6 ? Cj67z6 : Au1nz6[5]);
assign O0s7v6 = (Pz1yx6 ? Ui67z6 : Au1nz6[4]);
assign H0s7v6 = (Pz1yx6 ? Mi67z6 : Au1nz6[3]);
assign A0s7v6 = (Pz1yx6 ? Ei67z6 : Au1nz6[2]);
assign Tzr7v6 = (Pz1yx6 ? Wh67z6 : Au1nz6[1]);
assign Pz1yx6 = (Xz1yx6 & F02yx6);
assign Xz1yx6 = (~(N02yx6 | V02yx6));
assign Mzr7v6 = (D12yx6 ? Ak67z6 : Zs1nz6[0]);
assign Fzr7v6 = (D12yx6 ? Sj67z6 : Zs1nz6[7]);
assign Yyr7v6 = (D12yx6 ? Kj67z6 : Zs1nz6[6]);
assign Ryr7v6 = (D12yx6 ? Cj67z6 : Zs1nz6[5]);
assign Kyr7v6 = (D12yx6 ? Ui67z6 : Zs1nz6[4]);
assign Dyr7v6 = (D12yx6 ? Mi67z6 : Zs1nz6[3]);
assign Wxr7v6 = (D12yx6 ? Ei67z6 : Zs1nz6[2]);
assign Pxr7v6 = (D12yx6 ? Wh67z6 : Zs1nz6[1]);
assign D12yx6 = (L12yx6 & V02yx6);
assign L12yx6 = (~(T12yx6 | N02yx6));
assign Ixr7v6 = (B22yx6 ? Ak67z6 : Yr1nz6[0]);
assign Bxr7v6 = (B22yx6 ? Sj67z6 : Yr1nz6[7]);
assign Uwr7v6 = (B22yx6 ? Kj67z6 : Yr1nz6[6]);
assign Nwr7v6 = (B22yx6 ? Cj67z6 : Yr1nz6[5]);
assign Gwr7v6 = (B22yx6 ? Ui67z6 : Yr1nz6[4]);
assign Zvr7v6 = (B22yx6 ? Mi67z6 : Yr1nz6[3]);
assign Svr7v6 = (B22yx6 ? Ei67z6 : Yr1nz6[2]);
assign Lvr7v6 = (B22yx6 ? Wh67z6 : Yr1nz6[1]);
assign B22yx6 = (J22yx6 & N02yx6);
assign J22yx6 = (F02yx6 & R22yx6);
assign R22yx6 = (!V02yx6);
assign Evr7v6 = (~(Z22yx6 & H32yx6));
assign H32yx6 = (P32yx6 | X32yx6);
assign P32yx6 = (!F42yx6);
assign Z22yx6 = (~(Ja1nz6[2] & T12yx6));
assign Xur7v6 = (~(N42yx6 & V42yx6));
assign V42yx6 = (~(F42yx6 & D52yx6));
assign D52yx6 = (Zy1yx6 ^ X32yx6);
assign X32yx6 = (Ja1nz6[2] ? T52yx6 : L52yx6);
assign T52yx6 = (N02yx6 & B62yx6);
assign L52yx6 = (~(N02yx6 & V02yx6));
assign N42yx6 = (~(Ja1nz6[1] & T12yx6));
assign Qur7v6 = (~(J62yx6 & R62yx6));
assign R62yx6 = (~(F42yx6 & Z62yx6));
assign Z62yx6 = (Zy1yx6 ^ B62yx6);
assign Zy1yx6 = (~(H72yx6 & P72yx6));
assign H72yx6 = (V02yx6 ^ N02yx6);
assign F42yx6 = (~(T12yx6 | Hae7v6));
assign J62yx6 = (~(Ja1nz6[0] & T12yx6));
assign Jur7v6 = (Ry1yx6 ? X72yx6 : Bv1nz6[0]);
assign X72yx6 = (~(B62yx6 & F82yx6));
assign F82yx6 = (~(Ak67z6 & Cc5ov6));
assign B62yx6 = (V02yx6 | N82yx6);
assign Cur7v6 = (Ry1yx6 ? Sj67z6 : Xq1nz6[7]);
assign Vtr7v6 = (Ry1yx6 ? Kj67z6 : Xq1nz6[6]);
assign Otr7v6 = (Ry1yx6 ? Cj67z6 : Xq1nz6[5]);
assign Htr7v6 = (Ry1yx6 ? Ui67z6 : Xq1nz6[4]);
assign Atr7v6 = (Ry1yx6 ? Mi67z6 : Xq1nz6[3]);
assign Tsr7v6 = (Ry1yx6 ? Ei67z6 : Xq1nz6[2]);
assign Ry1yx6 = (F02yx6 & V82yx6);
assign V82yx6 = (~(Cc5ov6 & D92yx6));
assign D92yx6 = (~(L92yx6 & T92yx6));
assign F02yx6 = (!T12yx6);
assign T12yx6 = (~(Dniiw6 & Ba2yx6));
assign Ba2yx6 = (~(P72yx6 & Ja2yx6));
assign Ja2yx6 = (~(Ra2yx6 & W197z6));
assign Ra2yx6 = (~(Za2yx6 | Eee7v6));
assign Msr7v6 = (Xb2yx6 ? Pb2yx6 : Hb2yx6);
assign Fsr7v6 = (Ah2nz6[2] ? Nc2yx6 : Fc2yx6);
assign Nc2yx6 = (Vc2yx6 | Dd2yx6);
assign Dd2yx6 = (~(Ld2yx6 | Ah2nz6[1]));
assign Fc2yx6 = (Td2yx6 & Ah2nz6[1]);
assign Yrr7v6 = (Xb2yx6 ? Mwf7v6 : Be2yx6);
assign Rrr7v6 = (Nl1nz6[0] & Je2yx6);
assign Je2yx6 = (~(Re2yx6 & Ze2yx6));
assign Ze2yx6 = (~(Ctf7v6 & Hf2yx6));
assign Hf2yx6 = (!Vuf7v6);
assign Re2yx6 = (~(Pf2yx6 | Xf2yx6));
assign Pf2yx6 = (~(Pb2yx6 | Mwf7v6));
assign Krr7v6 = (!Fg2yx6);
assign Fg2yx6 = (Ah2nz6[0] ? Vg2yx6 : Ng2yx6);
assign Ng2yx6 = (~(Dh2yx6 & Vg2yx6));
assign Drr7v6 = (Ah2nz6[1] ? Vc2yx6 : Td2yx6);
assign Vc2yx6 = (~(Vg2yx6 & Lh2yx6));
assign Lh2yx6 = (Ld2yx6 | Ah2nz6[0]);
assign Td2yx6 = (Th2yx6 & Ah2nz6[0]);
assign Th2yx6 = (Dh2yx6 & Vg2yx6);
assign Vg2yx6 = (~(Bi2yx6 & Ji2yx6));
assign Ji2yx6 = (Ri2yx6 | Pb2yx6);
assign Bi2yx6 = (~(Nl1nz6[0] & V91nv6));
assign Dh2yx6 = (!Ld2yx6);
assign Wqr7v6 = (Xb2yx6 ? M2e7v6 : Zi2yx6);
assign Xb2yx6 = (Hj2yx6 & Pj2yx6);
assign Pj2yx6 = (~(Xj2yx6 & Fk2yx6));
assign Fk2yx6 = (~(Nk2yx6 & Twhiw6));
assign Nk2yx6 = (~(Vuf7v6 & Vk2yx6));
assign Vk2yx6 = (~(Qk77z6 & Dl2yx6));
assign Xj2yx6 = (Ll2yx6 & Tl2yx6);
assign Ll2yx6 = (~(Bm2yx6 & Pb2yx6));
assign Bm2yx6 = (~(Jm2yx6 & Nl1nz6[1]));
assign Jm2yx6 = (~(Rm2yx6 | Nl1nz6[0]));
assign Hj2yx6 = (Zm2yx6 & Ri2yx6);
assign Ri2yx6 = (~(Mwf7v6 & Xf2yx6));
assign Zm2yx6 = (Nl1nz6[1] | Hn2yx6);
assign Hn2yx6 = (Pn2yx6 & Xn2yx6);
assign Xn2yx6 = (~(Fo2yx6 & No2yx6));
assign No2yx6 = (Vo2yx6 & Dp2yx6);
assign Vo2yx6 = (~(Kf2nz6[1] | Kf2nz6[2]));
assign Fo2yx6 = (Lp2yx6 & Dl2yx6);
assign Lp2yx6 = (~(Ld2yx6 | Xf2yx6));
assign Pn2yx6 = (~(Tp2yx6 & Bq2yx6));
assign Bq2yx6 = (Jq2yx6 & Ah2nz6[0]);
assign Jq2yx6 = (Nl1nz6[0] & V91nv6);
assign Tp2yx6 = (Ah2nz6[2] & Ah2nz6[1]);
assign Zi2yx6 = (~(Hb2yx6 | Be2yx6));
assign Be2yx6 = (~(Rq2yx6 & Zq2yx6));
assign Zq2yx6 = (Qk77z6 | Dl2yx6);
assign Rq2yx6 = (~(Tl2yx6 & Twhiw6));
assign Hb2yx6 = (~(Hr2yx6 & Pr2yx6));
assign Pr2yx6 = (~(Tl2yx6 & Xr2yx6));
assign Xr2yx6 = (~(Qk77z6 & Twhiw6));
assign Hr2yx6 = (!Fs2yx6);
assign Pqr7v6 = (Ns2yx6 ^ Vs2yx6);
assign Iqr7v6 = (Eb1nv6 ^ Dt2yx6);
assign Bqr7v6 = (Ec2nz6[2] ^ Lt2yx6);
assign Upr7v6 = (Ec2nz6[3] ^ Tt2yx6);
assign Tt2yx6 = (Lt2yx6 & Ec2nz6[2]);
assign Lt2yx6 = (~(Dt2yx6 | Eb1nv6));
assign Npr7v6 = (Vs2yx6 ? Dxe7v6 : Bu2yx6);
assign Gpr7v6 = (~(Ju2yx6 & Ru2yx6));
assign Ru2yx6 = (~(B5e7v6 & M8e7v6));
assign Zor7v6 = (~(Zu2yx6 & Hv2yx6));
assign Hv2yx6 = (~(Pv2yx6 & Xv2yx6));
assign Sor7v6 = (Pv2yx6 ? R0f7v6 : Xv2yx6);
assign Lor7v6 = (~(Fw2yx6 & Nw2yx6));
assign Nw2yx6 = (Vw2yx6 | Dxe7v6);
assign Vw2yx6 = (~(Kve7v6 | Dx2yx6));
assign Dx2yx6 = (~(Lx2yx6 | Vs2yx6));
assign Fw2yx6 = (~(Kve7v6 & Vs2yx6));
assign Eor7v6 = (T32nz6[0] ? By2yx6 : Tx2yx6);
assign Xnr7v6 = (T32nz6[1] ? Ry2yx6 : Jy2yx6);
assign Qnr7v6 = (!Zy2yx6);
assign Zy2yx6 = (T32nz6[2] ? Pz2yx6 : Hz2yx6);
assign Hz2yx6 = (~(Jy2yx6 & T32nz6[1]));
assign Jnr7v6 = (T32nz6[3] ? F03yx6 : Xz2yx6);
assign F03yx6 = (~(Pz2yx6 & N03yx6));
assign N03yx6 = (T32nz6[2] | Kve7v6);
assign Pz2yx6 = (~(Ry2yx6 | V03yx6));
assign V03yx6 = (~(T32nz6[1] | Kve7v6));
assign Ry2yx6 = (By2yx6 | D13yx6);
assign D13yx6 = (~(T32nz6[0] | Kve7v6));
assign By2yx6 = (Vs2yx6 | L13yx6);
assign L13yx6 = (~(Bu2yx6 | Kve7v6));
assign Xz2yx6 = (T13yx6 & Jy2yx6);
assign Jy2yx6 = (Tx2yx6 & T32nz6[0]);
assign Tx2yx6 = (B23yx6 & Bu2yx6);
assign Bu2yx6 = (!J23yx6);
assign B23yx6 = (~(Vs2yx6 | Kve7v6));
assign Cnr7v6 = (Z23yx6 ? R23yx6 : Yb1nz6[0]);
assign R23yx6 = (~(H33yx6 ^ P33yx6));
assign Vmr7v6 = (Z23yx6 ? X33yx6 : Yb1nz6[1]);
assign X33yx6 = (F43yx6 ^ H33yx6);
assign H33yx6 = (~(N43yx6 ^ P33yx6));
assign Omr7v6 = (Z23yx6 ? F43yx6 : Yb1nz6[2]);
assign Z23yx6 = (V43yx6 & D53yx6);
assign V43yx6 = (~(L53yx6 & T53yx6));
assign T53yx6 = (~(B63yx6 & V91nv6));
assign F43yx6 = (~(J63yx6 ^ Yb1nz6[2]));
assign J63yx6 = (~(R63yx6 & P33yx6));
assign P33yx6 = (Z63yx6 | H73yx6);
assign Hmr7v6 = (P73yx6 & Ci6ft6);
assign P73yx6 = (X73yx6 & F83yx6);
assign F83yx6 = (Ak6ft6 | Og6ft6);
assign X73yx6 = (~(N83yx6 & V83yx6));
assign V83yx6 = (D93yx6 & L93yx6);
assign L93yx6 = (T93yx6 & Ba3yx6);
assign Ba3yx6 = (N02yx6 ^ Ja3yx6);
assign N02yx6 = (Hae7v6 ? Bv1nz6[1] : T92yx6);
assign T93yx6 = (~(V02yx6 ^ Ra3yx6));
assign V02yx6 = (Hae7v6 ? Bv1nz6[0] : L92yx6);
assign D93yx6 = (Za3yx6 & Hb3yx6);
assign Hb3yx6 = (~(Ul5ov6 ^ Pb3yx6));
assign Za3yx6 = (Nl5ov6 ^ Xb3yx6);
assign N83yx6 = (Fc3yx6 & Nc3yx6);
assign Nc3yx6 = (~(Lj1nz6[2] ^ Ja1nz6[2]));
assign Fc3yx6 = (Vc3yx6 & Hbe7v6);
assign Vc3yx6 = (~(Hi1nz6[2] ^ U81nz6[2]));
assign Amr7v6 = (Ab5ov6 ? Dd3yx6 : Pp1nz6[0]);
assign Dd3yx6 = (~(Ld5ov6 & Ld3yx6));
assign Ld3yx6 = (~(Zd5ov6 & Cc5ov6));
assign Zd5ov6 = (~(Td3yx6 & Be3yx6));
assign Be3yx6 = (~(V7xmz6[0] & Pf5ov6));
assign Td3yx6 = (I347v6 ? Re3yx6 : Je3yx6);
assign Re3yx6 = (Ze3yx6 & Hf3yx6);
assign Hf3yx6 = (Pf3yx6 & Xf3yx6);
assign Xf3yx6 = (~(Mh5ov6 & Vcxmz6[21]));
assign Pf3yx6 = (~(Vcxmz6[0] & Gjfnv6));
assign Ze3yx6 = (Fg3yx6 & Ng3yx6);
assign Ng3yx6 = (~(Hi5ov6 & Vcxmz6[14]));
assign Fg3yx6 = (~(Oi5ov6 & Vcxmz6[7]));
assign Je3yx6 = (Vg3yx6 & Dh3yx6);
assign Dh3yx6 = (Lh3yx6 & Th3yx6);
assign Th3yx6 = (~(Mh5ov6 & Vcxmz6[47]));
assign Lh3yx6 = (~(Gjfnv6 & Vcxmz6[26]));
assign Vg3yx6 = (Bi3yx6 & Ji3yx6);
assign Ji3yx6 = (~(Hi5ov6 & Vcxmz6[40]));
assign Bi3yx6 = (~(Oi5ov6 & Vcxmz6[33]));
assign Ld5ov6 = (Ul5ov6 | Ri3yx6);
assign Tlr7v6 = (~(Zi3yx6 & Hj3yx6));
assign Hj3yx6 = (~(Kwvmz6[1] & Pj3yx6));
assign Mlr7v6 = (~(Xj3yx6 & Fk3yx6));
assign Fk3yx6 = (~(Kwvmz6[2] & Pj3yx6));
assign Flr7v6 = (~(Nk3yx6 & Vk3yx6));
assign Vk3yx6 = (~(Kwvmz6[3] & Pj3yx6));
assign Ykr7v6 = (~(Dl3yx6 & Ll3yx6));
assign Ll3yx6 = (~(Kwvmz6[4] & Pj3yx6));
assign Rkr7v6 = (~(Tl3yx6 & Bm3yx6));
assign Bm3yx6 = (~(Kwvmz6[0] & Pj3yx6));
assign Kkr7v6 = (Jm3yx6 ^ Rm3yx6);
assign Dkr7v6 = (~(Zm3yx6 ^ Hn3yx6));
assign Hn3yx6 = (~(Rm3yx6 | Jm3yx6));
assign Jm3yx6 = (Pn3yx6 & Xn3yx6);
assign Xn3yx6 = (Zi3yx6 | Fo3yx6);
assign Wjr7v6 = (No3yx6 ? Jt37v6 : Fo3yx6);
assign Pjr7v6 = (Ci6ft6 & Vo3yx6);
assign Vo3yx6 = (~(Og6ft6 & Dp3yx6));
assign Dp3yx6 = (Lp3yx6 | Ak6ft6);
assign Lp3yx6 = (~(Tp3yx6 | Id6ft6));
assign Ijr7v6 = (~(Bq3yx6 & Jq3yx6));
assign Jq3yx6 = (Rq3yx6 | Zq3yx6);
assign Bq3yx6 = (~(Hr3yx6 & Vis7z6[5]));
assign Bjr7v6 = (Vis7z6[4] ? Xr3yx6 : Pr3yx6);
assign Xr3yx6 = (~(Fs3yx6 & Ns3yx6));
assign Ns3yx6 = (~(Vs3yx6 & Dt3yx6));
assign Pr3yx6 = (Vs3yx6 & Lt3yx6);
assign Uir7v6 = (Tt3yx6 ? Vs3yx6 : Hr3yx6);
assign Nir7v6 = (Ru3yx6 ? Ju3yx6 : Bu3yx6);
assign Ru3yx6 = (!Vis7z6[1]);
assign Ju3yx6 = (Vs3yx6 & Vis7z6[0]);
assign Bu3yx6 = (~(Zu3yx6 & Hv3yx6));
assign Hv3yx6 = (~(Vs3yx6 & Tt3yx6));
assign Tt3yx6 = (!Vis7z6[0]);
assign Gir7v6 = (~(Pv3yx6 & Xv3yx6));
assign Xv3yx6 = (~(Vs3yx6 & Fw3yx6));
assign Fw3yx6 = (Vis7z6[2] ^ Nw3yx6);
assign Nw3yx6 = (Vis7z6[1] & Vis7z6[0]);
assign Pv3yx6 = (~(Hr3yx6 & Vis7z6[2]));
assign Zhr7v6 = (!Vw3yx6);
assign Vw3yx6 = (Vis7z6[3] ? Fs3yx6 : Dx3yx6);
assign Fs3yx6 = (Zu3yx6 & Lx3yx6);
assign Lx3yx6 = (~(Vs3yx6 & Tx3yx6));
assign Dx3yx6 = (Rq3yx6 | Tx3yx6);
assign Rq3yx6 = (!Vs3yx6);
assign Vs3yx6 = (By3yx6 & Jy3yx6);
assign Jy3yx6 = (~(Ry3yx6 | Zy3yx6));
assign By3yx6 = (~(Hz3yx6 | Hr3yx6));
assign Hr3yx6 = (!Zu3yx6);
assign Zu3yx6 = (~(Pz3yx6 & Xz3yx6));
assign Pz3yx6 = (~(Hz3yx6 | Zy3yx6));
assign Shr7v6 = (~(F04yx6 & N04yx6));
assign N04yx6 = (~(Sl37v6 & V04yx6));
assign F04yx6 = (~(D14yx6 & P7s7z6[8]));
assign Lhr7v6 = (~(L14yx6 & T14yx6));
assign T14yx6 = (~(Iw27v6 & V04yx6));
assign L14yx6 = (~(P7s7z6[30] & D14yx6));
assign Ehr7v6 = (E46ft6 ? J24yx6 : B24yx6);
assign B24yx6 = (R24yx6 & Z24yx6);
assign R24yx6 = (~(H34yx6 & P34yx6));
assign P34yx6 = (~(X34yx6 & F44yx6));
assign F44yx6 = (N44yx6 & V44yx6);
assign V44yx6 = (D54yx6 & L54yx6);
assign D54yx6 = (~(P7s7z6[26] | P7s7z6[8]));
assign X34yx6 = (T54yx6 & B64yx6);
assign B64yx6 = (~(J64yx6 | P7s7z6[17]));
assign J64yx6 = (P7s7z6[18] | P7s7z6[20]);
assign T54yx6 = (R64yx6 & Z64yx6);
assign H34yx6 = (~(Fho7v6 & H74yx6));
assign H74yx6 = (~(P74yx6 & X74yx6));
assign X74yx6 = (F84yx6 & N84yx6);
assign N84yx6 = (~(P7s7z6[8] | P7s7z6[9]));
assign P74yx6 = (V84yx6 & D94yx6);
assign V84yx6 = (~(L94yx6 | P7s7z6[10]));
assign Xgr7v6 = (~(T94yx6 & Ba4yx6));
assign Ba4yx6 = (~(Lk37v6 & V04yx6));
assign T94yx6 = (~(D14yx6 & P7s7z6[9]));
assign Qgr7v6 = (~(Ja4yx6 & Ra4yx6));
assign Ra4yx6 = (~(Ej37v6 & V04yx6));
assign Ja4yx6 = (~(D14yx6 & P7s7z6[10]));
assign Jgr7v6 = (~(Za4yx6 & Hb4yx6));
assign Hb4yx6 = (~(Xh37v6 & V04yx6));
assign Za4yx6 = (~(P7s7z6[11] & D14yx6));
assign Cgr7v6 = (~(Pb4yx6 & Xb4yx6));
assign Xb4yx6 = (~(Qg37v6 & V04yx6));
assign Pb4yx6 = (~(P7s7z6[12] & D14yx6));
assign Vfr7v6 = (~(Fc4yx6 & Nc4yx6));
assign Nc4yx6 = (~(Jf37v6 & V04yx6));
assign Fc4yx6 = (~(P7s7z6[13] & D14yx6));
assign Ofr7v6 = (~(Vc4yx6 & Dd4yx6));
assign Dd4yx6 = (~(Ce37v6 & V04yx6));
assign Vc4yx6 = (~(P7s7z6[14] & D14yx6));
assign Hfr7v6 = (~(Ld4yx6 & Td4yx6));
assign Td4yx6 = (~(Vc37v6 & V04yx6));
assign Ld4yx6 = (~(P7s7z6[16] & D14yx6));
assign Afr7v6 = (~(Be4yx6 & Je4yx6));
assign Je4yx6 = (~(Ob37v6 & V04yx6));
assign Be4yx6 = (~(P7s7z6[17] & D14yx6));
assign Ter7v6 = (~(Re4yx6 & Ze4yx6));
assign Ze4yx6 = (~(Ha37v6 & V04yx6));
assign Re4yx6 = (~(P7s7z6[18] & D14yx6));
assign Mer7v6 = (~(Hf4yx6 & Pf4yx6));
assign Pf4yx6 = (~(A937v6 & V04yx6));
assign Hf4yx6 = (~(P7s7z6[19] & D14yx6));
assign Fer7v6 = (~(Xf4yx6 & Fg4yx6));
assign Fg4yx6 = (~(T737v6 & V04yx6));
assign Xf4yx6 = (~(P7s7z6[20] & D14yx6));
assign Ydr7v6 = (~(Ng4yx6 & Vg4yx6));
assign Vg4yx6 = (~(M637v6 & V04yx6));
assign Ng4yx6 = (~(P7s7z6[21] & D14yx6));
assign Rdr7v6 = (~(Dh4yx6 & Lh4yx6));
assign Lh4yx6 = (~(F537v6 & V04yx6));
assign Dh4yx6 = (~(P7s7z6[22] & D14yx6));
assign Kdr7v6 = (~(Th4yx6 & Bi4yx6));
assign Bi4yx6 = (~(Y337v6 & V04yx6));
assign Th4yx6 = (~(P7s7z6[24] & D14yx6));
assign Ddr7v6 = (~(Ji4yx6 & Ri4yx6));
assign Ri4yx6 = (~(R237v6 & V04yx6));
assign Ji4yx6 = (~(P7s7z6[25] & D14yx6));
assign Wcr7v6 = (~(Zi4yx6 & Hj4yx6));
assign Hj4yx6 = (~(K137v6 & V04yx6));
assign Zi4yx6 = (~(P7s7z6[26] & D14yx6));
assign Pcr7v6 = (~(Pj4yx6 & Xj4yx6));
assign Xj4yx6 = (~(D037v6 & V04yx6));
assign Pj4yx6 = (~(P7s7z6[27] & D14yx6));
assign Icr7v6 = (~(Fk4yx6 & Nk4yx6));
assign Nk4yx6 = (~(Wy27v6 & V04yx6));
assign Fk4yx6 = (~(P7s7z6[28] & D14yx6));
assign Bcr7v6 = (~(Vk4yx6 & Dl4yx6));
assign Dl4yx6 = (~(Px27v6 & V04yx6));
assign V04yx6 = (J24yx6 & Ll4yx6);
assign Ll4yx6 = (!D14yx6);
assign Vk4yx6 = (~(P7s7z6[29] & D14yx6));
assign D14yx6 = (J24yx6 & Tl4yx6);
assign Tl4yx6 = (~(Bm4yx6 & Ldo7v6));
assign Ubr7v6 = (~(Jm4yx6 & Rm4yx6));
assign Rm4yx6 = (~(Zm4yx6 & E46ft6));
assign Zm4yx6 = (Hn4yx6 & Eifnv6);
assign Jm4yx6 = (~(Nu27v6 & J24yx6));
assign Nbr7v6 = (~(Pn4yx6 & Xn4yx6));
assign Xn4yx6 = (~(Ur37v6 & Fo4yx6));
assign Pn4yx6 = (~(Txadt6 & X66ft6));
assign Gbr7v6 = (~(No4yx6 ^ Vo4yx6));
assign Vo4yx6 = (Lp4yx6 ? No4yx6 : Dp4yx6);
assign Zar7v6 = (Tp4yx6 ? X9s7z6[1] : Zas7z6[1]);
assign Sar7v6 = (Tp4yx6 ? X9s7z6[3] : Or27v6);
assign Lar7v6 = (Tp4yx6 ? X9s7z6[4] : Hq27v6);
assign Ear7v6 = (Tp4yx6 ? X9s7z6[5] : Ap27v6);
assign X9r7v6 = (Tp4yx6 ? X9s7z6[6] : Tn27v6);
assign Q9r7v6 = (Tp4yx6 ? X9s7z6[7] : Mm27v6);
assign J9r7v6 = (Tp4yx6 ? X9s7z6[8] : U42nv6);
assign C9r7v6 = (Tp4yx6 ? X9s7z6[9] : B52nv6);
assign V8r7v6 = (Tp4yx6 ? X9s7z6[10] : I52nv6);
assign O8r7v6 = (Tp4yx6 ? X9s7z6[11] : P52nv6);
assign H8r7v6 = (Tp4yx6 ? X9s7z6[12] : W52nv6);
assign A8r7v6 = (Tp4yx6 ? X9s7z6[13] : D62nv6);
assign T7r7v6 = (Tp4yx6 ? X9s7z6[14] : K62nv6);
assign M7r7v6 = (Tp4yx6 ? X9s7z6[15] : R62nv6);
assign F7r7v6 = (Tp4yx6 ? X9s7z6[16] : U47iw6);
assign Y6r7v6 = (Tp4yx6 ? X9s7z6[17] : J27iw6);
assign R6r7v6 = (Tp4yx6 ? X9s7z6[18] : H17iw6);
assign K6r7v6 = (Tp4yx6 ? X9s7z6[19] : Dz6iw6);
assign D6r7v6 = (Tp4yx6 ? X9s7z6[20] : Emhov6);
assign W5r7v6 = (Tp4yx6 ? X9s7z6[21] : Guhov6);
assign P5r7v6 = (Tp4yx6 ? X9s7z6[22] : Bk6iw6);
assign I5r7v6 = (Tp4yx6 ? X9s7z6[23] : Z0iov6);
assign B5r7v6 = (Tp4yx6 ? X9s7z6[24] : Is5iw6);
assign U4r7v6 = (Tp4yx6 ? X9s7z6[25] : Gr5iw6);
assign N4r7v6 = (Tp4yx6 ? X9s7z6[26] : Jp5iw6);
assign G4r7v6 = (Tp4yx6 ? X9s7z6[27] : Mn5iw6);
assign Z3r7v6 = (Tp4yx6 ? X9s7z6[28] : Bl5iw6);
assign S3r7v6 = (Tp4yx6 ? X9s7z6[29] : Ej5iw6);
assign L3r7v6 = (Tp4yx6 ? X9s7z6[30] : D85iw6);
assign E3r7v6 = (Tp4yx6 ? X9s7z6[31] : Cx4iw6);
assign X2r7v6 = (Tp4yx6 ? X9s7z6[32] : Wf4iw6);
assign Q2r7v6 = (Tp4yx6 ? X9s7z6[33] : Iklov6);
assign J2r7v6 = (Tp4yx6 ? X9s7z6[34] : E64iw6);
assign Tp4yx6 = (!Bq4yx6);
assign C2r7v6 = (Bq4yx6 ? H44iw6 : X9s7z6[35]);
assign V1r7v6 = (Bq4yx6 ? W14iw6 : X9s7z6[36]);
assign O1r7v6 = (Bq4yx6 ? Zz3iw6 : X9s7z6[37]);
assign H1r7v6 = (Bq4yx6 ? Ro3iw6 : X9s7z6[38]);
assign A1r7v6 = (Bq4yx6 ? X0hov6 : X9s7z6[39]);
assign T0r7v6 = (Bq4yx6 ? Zas7z6[0] : X9s7z6[0]);
assign M0r7v6 = (Lp4yx6 ? Rq4yx6 : Jq4yx6);
assign Rq4yx6 = (~(No4yx6 | Dp4yx6));
assign Jq4yx6 = (Zas7z6[2] & Zq4yx6);
assign Zq4yx6 = (~(Orhov6 & Hr4yx6));
assign Orhov6 = (!U42nv6);
assign F0r7v6 = (Bq4yx6 ? Zas7z6[2] : Tl6ft6);
assign Bq4yx6 = (Lp4yx6 & Pr4yx6);
assign Lp4yx6 = (Xr4yx6 & Fs4yx6);
assign Fs4yx6 = (Ci27v6 & Ns4yx6);
assign Ns4yx6 = (~(Vs4yx6 & C397z6));
assign Vs4yx6 = (Mm27v6 ? Lt4yx6 : Dt4yx6);
assign Lt4yx6 = (Tt4yx6 ? Scs7z6[2] : Scs7z6[3]);
assign Dt4yx6 = (Tt4yx6 ? Scs7z6[0] : Scs7z6[1]);
assign Xr4yx6 = (Rj27v6 & Fl27v6);
assign Yzq7v6 = (~(Bu4yx6 & Ju4yx6));
assign Ju4yx6 = (~(Xwadt6 & Ru4yx6));
assign Ru4yx6 = (~(Zu4yx6 & K4a8x6));
assign Bu4yx6 = (K4a8x6 | Nw5ft6);
assign K4a8x6 = (!T5a8x6);
assign Rzq7v6 = (Hv4yx6 & Xwadt6);
assign Hv4yx6 = (Pv4yx6 & Xv4yx6);
assign Pv4yx6 = (T5a8x6 | Nw5ft6);
assign T5a8x6 = (~(Fw4yx6 & Nw4yx6));
assign Nw4yx6 = (Az98x6 & S1a8x6);
assign S1a8x6 = (~(D9r7x6 & Vw4yx6));
assign Vw4yx6 = (~(O75ft6 & Jc4iw6));
assign D9r7x6 = (Dx4yx6 & Kjo7x6);
assign Kjo7x6 = (!N2a8x6);
assign Dx4yx6 = (~(Lx4yx6 & Tx4yx6));
assign Tx4yx6 = (~(Hmp7z6[1] & By4yx6));
assign Lx4yx6 = (Jy4yx6 & Ry4yx6);
assign Ry4yx6 = (~(Dm2ft6 & Fko7x6));
assign Fko7x6 = (~(Mko7x6 & Veo7x6));
assign Jy4yx6 = (Veo7x6 | Zy4yx6);
assign Az98x6 = (~(S2fiw6 & Hz4yx6));
assign Hz4yx6 = (~(Fy4ft6 & Jc4iw6));
assign S2fiw6 = (Pz4yx6 & V0fiw6);
assign Pz4yx6 = (~(Xz4yx6 & F05yx6));
assign F05yx6 = (~(Hyp7z6[1] & E2fiw6));
assign Xz4yx6 = (N05yx6 & V05yx6);
assign V05yx6 = (L2fiw6 | X1fiw6);
assign L2fiw6 = (!Gs2ft6);
assign N05yx6 = (~(D15yx6 & Hyp7z6[0]));
assign Fw4yx6 = (E99ov6 & Q8o7x6);
assign Q8o7x6 = (~(L15yx6 & Y5o7x6));
assign L15yx6 = (T15yx6 & O7o7x6);
assign O7o7x6 = (~(B25yx6 & J25yx6));
assign J25yx6 = (~(I7p7z6[1] & R25yx6));
assign B25yx6 = (Z25yx6 & H35yx6);
assign H35yx6 = (~(M12ft6 & A7o7x6));
assign A7o7x6 = (R25yx6 | P35yx6);
assign Z25yx6 = (~(P35yx6 & I7p7z6[0]));
assign T15yx6 = (~(Um4ft6 & Jc4iw6));
assign E99ov6 = (~(Yx98x6 & X35yx6));
assign X35yx6 = (~(Mi5ft6 & Jc4iw6));
assign Yx98x6 = (F45yx6 & Ryeiw6);
assign Ryeiw6 = (!Wxeiw6);
assign F45yx6 = (~(N45yx6 & V45yx6));
assign V45yx6 = (~(Sgp7z6[1] & Tzeiw6));
assign N45yx6 = (D55yx6 & L55yx6);
assign L55yx6 = (~(Ei2ft6 & Mzeiw6));
assign Mzeiw6 = (Tzeiw6 | T55yx6);
assign D55yx6 = (~(T55yx6 & Sgp7z6[0]));
assign T55yx6 = (!F6fiw6);
assign Kzq7v6 = (~(B65yx6 & J65yx6));
assign J65yx6 = (~(Uur7z6[1] & R65yx6));
assign R65yx6 = (Z65yx6 | H75yx6);
assign B65yx6 = (Lhliw6 | Uur7z6[0]);
assign Dzq7v6 = (P75yx6 & Uur7z6[1]);
assign P75yx6 = (X75yx6 & Z65yx6);
assign Z65yx6 = (~(Zu4yx6 & F85yx6));
assign X75yx6 = (Uur7z6[0] | H75yx6);
assign H75yx6 = (!Lhliw6);
assign Wyq7v6 = (~(N85yx6 & V85yx6));
assign V85yx6 = (~(Hsr7z6[1] & D95yx6));
assign D95yx6 = (L95yx6 | T95yx6);
assign N85yx6 = (Inhiw6 | Hsr7z6[0]);
assign Pyq7v6 = (Ba5yx6 & Hsr7z6[1]);
assign Ba5yx6 = (Ja5yx6 & L95yx6);
assign L95yx6 = (~(Zu4yx6 & Ra5yx6));
assign Ja5yx6 = (Hsr7z6[0] | T95yx6);
assign T95yx6 = (!Inhiw6);
assign Inhiw6 = (~(Za5yx6 & Xkhiw6));
assign Za5yx6 = (Khhiw6 & Xkq7z6[12]);
assign Iyq7v6 = (~(Hb5yx6 & Pb5yx6));
assign Pb5yx6 = (~(Xb5yx6 & Fc5yx6));
assign Xb5yx6 = (~(C4s7z6[0] & Nc5yx6));
assign Byq7v6 = (Vc5yx6 & Dd5yx6);
assign Dd5yx6 = (~(Ld5yx6 & Td5yx6));
assign Td5yx6 = (!C4s7z6[0]);
assign Ld5yx6 = (!Fc5yx6);
assign Vc5yx6 = (!Hb5yx6);
assign Uxq7v6 = (~(Be5yx6 & Je5yx6));
assign Je5yx6 = (~(V1s7z6[0] & Re5yx6));
assign Nxq7v6 = (~(Ze5yx6 & Hf5yx6));
assign Hf5yx6 = (~(V1s7z6[1] & Re5yx6));
assign Gxq7v6 = (~(Pf5yx6 & Xf5yx6));
assign Xf5yx6 = (~(V1s7z6[2] & Re5yx6));
assign Zwq7v6 = (~(Fg5yx6 & Ng5yx6));
assign Ng5yx6 = (~(V1s7z6[3] & Re5yx6));
assign Swq7v6 = (~(Vg5yx6 & Dh5yx6));
assign Dh5yx6 = (~(V1s7z6[4] & Re5yx6));
assign Lwq7v6 = (~(Lh5yx6 & Th5yx6));
assign Th5yx6 = (~(V1s7z6[5] & Re5yx6));
assign Re5yx6 = (~(Bi5yx6 & Ji5yx6));
assign Ji5yx6 = (~(C4s7z6[0] & Ri5yx6));
assign Bi5yx6 = (Hb5yx6 & Fc5yx6);
assign Fc5yx6 = (~(Zi5yx6 & Hj5yx6));
assign Hj5yx6 = (Pj5yx6 & Lh5yx6);
assign Pj5yx6 = (Vg5yx6 & Fg5yx6);
assign Fg5yx6 = (~(Xj5yx6 & Fk5yx6));
assign Fk5yx6 = (Nk5yx6 & Pdq7z6[5]);
assign Nk5yx6 = (Pdq7z6[6] & Pdq7z6[7]);
assign Xj5yx6 = (Mja8x6 & Efa8x6);
assign Efa8x6 = (Vk5yx6 & Yba8x6);
assign Yba8x6 = (Paa8x6 & Pdq7z6[2]);
assign Paa8x6 = (Pdq7z6[1] & Pdq7z6[0]);
assign Vk5yx6 = (Pdq7z6[3] & Pdq7z6[4]);
assign Mja8x6 = (~(Dl5yx6 | Ll5yx6));
assign Dl5yx6 = (~(Hka8x6 & Pbadt6));
assign Hka8x6 = (Xkq7z6[20] & HTMDHBURST[0]);
assign Vg5yx6 = (~(Tl5yx6 & Bm5yx6));
assign Bm5yx6 = (Jm5yx6 & Tbq7z6[5]);
assign Jm5yx6 = (Tbq7z6[6] & Tbq7z6[7]);
assign Tl5yx6 = (Csgiw6 & Nngiw6);
assign Nngiw6 = (Rm5yx6 & Hkgiw6);
assign Hkgiw6 = (Yigiw6 & Tbq7z6[2]);
assign Yigiw6 = (Tbq7z6[1] & Tbq7z6[0]);
assign Rm5yx6 = (Tbq7z6[3] & Tbq7z6[4]);
assign Csgiw6 = (Zm5yx6 & Hn5yx6);
assign Zm5yx6 = (Xkq7z6[21] & Knbdt6);
assign Zi5yx6 = (Pn5yx6 & Be5yx6);
assign Be5yx6 = (~(Xn5yx6 & Fo5yx6));
assign Fo5yx6 = (No5yx6 & Cjq7z6[5]);
assign No5yx6 = (Cjq7z6[6] & Cjq7z6[7]);
assign Xn5yx6 = (Aya8x6 & Sta8x6);
assign Sta8x6 = (Vo5yx6 & Mqa8x6);
assign Mqa8x6 = (Dpa8x6 & Cjq7z6[2]);
assign Dpa8x6 = (Cjq7z6[1] & Cjq7z6[0]);
assign Vo5yx6 = (Cjq7z6[3] & Cjq7z6[4]);
assign Aya8x6 = (Dp5yx6 & Vya8x6);
assign Vya8x6 = (Xkq7z6[17] & HTMDHBURST[0]);
assign Dp5yx6 = (~(Ll5yx6 | Pbadt6));
assign Ll5yx6 = (~(Lp5yx6 & Tp5yx6));
assign Tp5yx6 = (Wfo7v6 & Tlmov6);
assign Lp5yx6 = (Oaadt6 & Bq5yx6);
assign Pn5yx6 = (Ze5yx6 & Pf5yx6);
assign Pf5yx6 = (~(Jq5yx6 & Rq5yx6));
assign Rq5yx6 = (Zq5yx6 & Kfq7z6[5]);
assign Zq5yx6 = (Kfq7z6[6] & Kfq7z6[7]);
assign Jq5yx6 = (L7hiw6 & W2hiw6);
assign W2hiw6 = (Hr5yx6 & Qzgiw6);
assign Qzgiw6 = (Hygiw6 & Kfq7z6[2]);
assign Hygiw6 = (Kfq7z6[1] & Kfq7z6[0]);
assign Hr5yx6 = (Kfq7z6[3] & Kfq7z6[4]);
assign L7hiw6 = (Pr5yx6 & Xkq7z6[19]);
assign Pr5yx6 = (HTMDHBURST[0] & Bnhiw6);
assign Ze5yx6 = (~(Xr5yx6 & Fs5yx6));
assign Fs5yx6 = (Ns5yx6 & Hhq7z6[5]);
assign Ns5yx6 = (Hhq7z6[6] & Hhq7z6[7]);
assign Xr5yx6 = (~(Rdliw6 | O8liw6));
assign O8liw6 = (~(Vs5yx6 & I5liw6));
assign I5liw6 = (S3liw6 & Hhq7z6[2]);
assign S3liw6 = (Hhq7z6[1] & Hhq7z6[0]);
assign Vs5yx6 = (Hhq7z6[3] & Hhq7z6[4]);
assign Rdliw6 = (~(Dt5yx6 & Lt5yx6));
assign Lt5yx6 = (Tt5yx6 & HTMDHBURST[0]);
assign Tt5yx6 = (~(Tlmov6 | Oaadt6));
assign Dt5yx6 = (Xkq7z6[18] & Bq5yx6);
assign Hb5yx6 = (~(C4s7z6[1] & Bu5yx6));
assign Bu5yx6 = (~(Zu4yx6 & Ju5yx6));
assign Lh5yx6 = (~(Ru5yx6 & Xkhiw6));
assign Xkhiw6 = (Zu5yx6 & Hv5yx6);
assign Hv5yx6 = (Pv5yx6 & Xv5yx6);
assign Xv5yx6 = (Xkq7z6[12] | Xkq7z6[22]);
assign Pv5yx6 = (Gy2ft6 ^ Fw5yx6);
assign Zu5yx6 = (~(Nw5yx6 | Vw5yx6));
assign Ru5yx6 = (Khhiw6 & Gmhiw6);
assign Gmhiw6 = (!Xkq7z6[12]);
assign Khhiw6 = (Dx5yx6 & Lx5yx6);
assign Lx5yx6 = (~(W3q7z6[2] | W3q7z6[3]));
assign Dx5yx6 = (~(W3q7z6[0] | W3q7z6[1]));
assign Ewq7v6 = (~(Tx5yx6 & By5yx6));
assign By5yx6 = (~(Ixr7z6[1] & Jy5yx6));
assign Jy5yx6 = (Ry5yx6 | Alo7x6);
assign Tx5yx6 = (Xy4ov6 | Ixr7z6[0]);
assign Xy4ov6 = (!Alo7x6);
assign Xvq7v6 = (~(Lz4ov6 & Zy5yx6));
assign Zy5yx6 = (~(Y4wmz6[0] & Hz5yx6));
assign Qvq7v6 = (Pz5yx6 ? Ez4ov6 : Gyvmz6[7]);
assign Ez4ov6 = (~(Xz5yx6 & F06yx6));
assign F06yx6 = (N06yx6 & V06yx6);
assign V06yx6 = (~(Iuvmz6[8] & D16yx6));
assign N06yx6 = (L16yx6 & T16yx6);
assign T16yx6 = (~(Iuvmz6[7] & B26yx6));
assign L16yx6 = (~(Iuvmz6[6] & J26yx6));
assign Xz5yx6 = (R26yx6 & Z26yx6);
assign Z26yx6 = (~(Iuvmz6[5] & H36yx6));
assign R26yx6 = (~(Iuvmz6[4] & P36yx6));
assign Jvq7v6 = (Y4wmz6[1] ^ Pz5yx6);
assign Cvq7v6 = (F46yx6 ? X36yx6 : D047v6);
assign X36yx6 = (!N46yx6);
assign Vuq7v6 = (V46yx6 ^ D56yx6);
assign Ouq7v6 = (~(L56yx6 ^ T56yx6));
assign T56yx6 = (~(D56yx6 | V46yx6));
assign D56yx6 = (~(B66yx6 & N46yx6));
assign B66yx6 = (D047v6 | J66yx6);
assign Huq7v6 = (~(R66yx6 & Z66yx6));
assign Z66yx6 = (H76yx6 | P76yx6);
assign Auq7v6 = (~(K5xmz6[1] ^ X76yx6));
assign Ttq7v6 = (~(F86yx6 & N86yx6));
assign N86yx6 = (V86yx6 | D96yx6);
assign Mtq7v6 = (Hwwmz6[1] ^ L96yx6);
assign Ftq7v6 = (Ba6yx6 ? Bv37v6 : T96yx6);
assign Ysq7v6 = (Ja6yx6 ^ Ra6yx6);
assign Rsq7v6 = (~(Za6yx6 ^ Hb6yx6));
assign Hb6yx6 = (~(Ra6yx6 | Ja6yx6));
assign Ja6yx6 = (Pb6yx6 & Xb6yx6);
assign Xb6yx6 = (Tl3yx6 | T96yx6);
assign Ksq7v6 = (~(Fc6yx6 & Nc6yx6));
assign Nc6yx6 = (Vc6yx6 | Dd6yx6);
assign Dsq7v6 = (Enwmz6[1] ^ Ld6yx6);
assign Wrq7v6 = (Be6yx6 ? Tw37v6 : Td6yx6);
assign Prq7v6 = (Je6yx6 ^ Re6yx6);
assign Irq7v6 = (~(Ze6yx6 ^ Hf6yx6));
assign Hf6yx6 = (~(Re6yx6 | Je6yx6));
assign Je6yx6 = (Pf6yx6 & Xf6yx6);
assign Xf6yx6 = (Dl3yx6 | Td6yx6);
assign Brq7v6 = (~(Fg6yx6 & Ng6yx6));
assign Ng6yx6 = (Vg6yx6 | Dh6yx6);
assign Uqq7v6 = (Bewmz6[1] ^ Lh6yx6);
assign Nqq7v6 = (Bi6yx6 ? Ly37v6 : Th6yx6);
assign Th6yx6 = (!Ji6yx6);
assign Gqq7v6 = (Ri6yx6 ^ Zi6yx6);
assign Zpq7v6 = (~(Hj6yx6 ^ Pj6yx6));
assign Pj6yx6 = (~(Zi6yx6 | Ri6yx6));
assign Ri6yx6 = (Xj6yx6 & Fk6yx6);
assign Fk6yx6 = (~(Nk6yx6 & Ji6yx6));
assign Spq7v6 = (Lh6yx6 ? Vk6yx6 : J7wmz6[7]);
assign Lpq7v6 = (Fg6yx6 ? N9wmz6[7] : Vk6yx6);
assign Vk6yx6 = (~(Dl6yx6 & Ll6yx6));
assign Ll6yx6 = (Tl6yx6 & Bm6yx6);
assign Bm6yx6 = (~(Iuvmz6[4] & D16yx6));
assign Tl6yx6 = (Jm6yx6 & Rm6yx6);
assign Rm6yx6 = (~(Iuvmz6[8] & B26yx6));
assign Jm6yx6 = (~(Iuvmz6[7] & J26yx6));
assign Dl6yx6 = (Zm6yx6 & Hn6yx6);
assign Hn6yx6 = (~(Iuvmz6[6] & H36yx6));
assign Zm6yx6 = (~(Iuvmz6[5] & P36yx6));
assign Epq7v6 = (~(Pn6yx6 & Xn6yx6));
assign Xn6yx6 = (~(Bi6yx6 & Sqvmz6[7]));
assign Pn6yx6 = (Fo6yx6 & No6yx6);
assign No6yx6 = (~(Vo6yx6 & J7wmz6[7]));
assign Fo6yx6 = (~(Dp6yx6 & N9wmz6[7]));
assign Xoq7v6 = (Ld6yx6 ? Lp6yx6 : Mgwmz6[7]);
assign Qoq7v6 = (Fc6yx6 ? Qiwmz6[7] : Lp6yx6);
assign Lp6yx6 = (~(Tp6yx6 & Bq6yx6));
assign Bq6yx6 = (Jq6yx6 & Rq6yx6);
assign Rq6yx6 = (~(Iuvmz6[5] & D16yx6));
assign Jq6yx6 = (Zq6yx6 & Hr6yx6);
assign Hr6yx6 = (~(Iuvmz6[4] & B26yx6));
assign Zq6yx6 = (~(Iuvmz6[8] & J26yx6));
assign Tp6yx6 = (Pr6yx6 & Xr6yx6);
assign Xr6yx6 = (~(Iuvmz6[7] & H36yx6));
assign Pr6yx6 = (~(Iuvmz6[6] & P36yx6));
assign Joq7v6 = (~(Fs6yx6 & Ns6yx6));
assign Ns6yx6 = (~(Be6yx6 & Xovmz6[7]));
assign Fs6yx6 = (Vs6yx6 & Dt6yx6);
assign Dt6yx6 = (~(Lt6yx6 & Mgwmz6[7]));
assign Vs6yx6 = (~(Tt6yx6 & Qiwmz6[7]));
assign Coq7v6 = (L96yx6 ? Bu6yx6 : Ppwmz6[7]);
assign Vnq7v6 = (F86yx6 ? Trwmz6[7] : Bu6yx6);
assign Bu6yx6 = (~(Ju6yx6 & Ru6yx6));
assign Ru6yx6 = (Zu6yx6 & Hv6yx6);
assign Hv6yx6 = (~(Iuvmz6[6] & D16yx6));
assign Zu6yx6 = (Pv6yx6 & Xv6yx6);
assign Xv6yx6 = (~(Iuvmz6[5] & B26yx6));
assign Pv6yx6 = (~(Iuvmz6[4] & J26yx6));
assign Ju6yx6 = (Fw6yx6 & Nw6yx6);
assign Nw6yx6 = (~(Iuvmz6[8] & H36yx6));
assign Fw6yx6 = (~(Iuvmz6[7] & P36yx6));
assign Onq7v6 = (~(Vw6yx6 & Dx6yx6));
assign Dx6yx6 = (~(Ba6yx6 & Cnvmz6[7]));
assign Vw6yx6 = (Lx6yx6 & Tx6yx6);
assign Tx6yx6 = (~(By6yx6 & Ppwmz6[7]));
assign Lx6yx6 = (~(Jy6yx6 & Trwmz6[7]));
assign Hnq7v6 = (X76yx6 ? Sywmz6[7] : Ry6yx6);
assign Anq7v6 = (R66yx6 ? W0xmz6[7] : Ry6yx6);
assign Ry6yx6 = (~(Zy6yx6 & Hz6yx6));
assign Hz6yx6 = (Pz6yx6 & Xz6yx6);
assign Xz6yx6 = (~(Iuvmz6[7] & D16yx6));
assign D16yx6 = (~(F07yx6 & N07yx6));
assign N07yx6 = (V07yx6 & D17yx6);
assign D17yx6 = (~(X9s7z6[15] & L17yx6));
assign V07yx6 = (T17yx6 & B27yx6);
assign B27yx6 = (~(J27yx6 & L94yx6));
assign T17yx6 = (~(Gqr7z6[7] & R27yx6));
assign F07yx6 = (Z27yx6 & H37yx6);
assign H37yx6 = (~(Wlr7z6[7] & P37yx6));
assign Z27yx6 = (X37yx6 & F47yx6);
assign F47yx6 = (~(Cor7z6[7] & N47yx6));
assign X37yx6 = (~(Tjr7z6[9] & V47yx6));
assign Pz6yx6 = (D57yx6 & L57yx6);
assign L57yx6 = (~(Iuvmz6[6] & B26yx6));
assign B26yx6 = (~(T57yx6 & B67yx6));
assign B67yx6 = (J67yx6 & R67yx6);
assign R67yx6 = (~(Cor7z6[15] & N47yx6));
assign J67yx6 = (~(Z67yx6 | H77yx6));
assign Z67yx6 = (Gqr7z6[15] & R27yx6);
assign T57yx6 = (P77yx6 & X77yx6);
assign X77yx6 = (~(X9s7z6[23] & L17yx6));
assign P77yx6 = (~(Wlr7z6[15] & P37yx6));
assign D57yx6 = (~(Iuvmz6[5] & J26yx6));
assign J26yx6 = (~(F87yx6 & N87yx6));
assign N87yx6 = (V87yx6 & D97yx6);
assign D97yx6 = (~(Cor7z6[23] & N47yx6));
assign V87yx6 = (~(Gqr7z6[23] & R27yx6));
assign F87yx6 = (L97yx6 & T97yx6);
assign T97yx6 = (~(Wlr7z6[23] & P37yx6));
assign L97yx6 = (~(X9s7z6[31] & L17yx6));
assign Zy6yx6 = (Ba7yx6 & Ja7yx6);
assign Ja7yx6 = (~(Iuvmz6[4] & H36yx6));
assign H36yx6 = (~(Ra7yx6 & Za7yx6));
assign Za7yx6 = (Hb7yx6 & Pb7yx6);
assign Pb7yx6 = (~(Cor7z6[31] & N47yx6));
assign Hb7yx6 = (~(Gqr7z6[31] & R27yx6));
assign Ra7yx6 = (Xb7yx6 & Fc7yx6);
assign Fc7yx6 = (~(Wlr7z6[31] & P37yx6));
assign Xb7yx6 = (~(X9s7z6[39] & L17yx6));
assign Ba7yx6 = (~(Iuvmz6[8] & P36yx6));
assign P36yx6 = (~(Nc7yx6 & Vc7yx6));
assign Vc7yx6 = (Dd7yx6 & Ld7yx6);
assign Nc7yx6 = (~(Td7yx6 | Be7yx6));
assign Td7yx6 = (X9s7z6[7] & L17yx6);
assign Tmq7v6 = (X76yx6 ? Sywmz6[3] : Je7yx6);
assign Mmq7v6 = (R66yx6 ? W0xmz6[3] : Je7yx6);
assign Je7yx6 = (~(Re7yx6 & Ze7yx6));
assign Ze7yx6 = (Hf7yx6 & Pf7yx6);
assign Pf7yx6 = (~(Iuvmz6[8] & Xf7yx6));
assign Hf7yx6 = (Fg7yx6 & Ng7yx6);
assign Ng7yx6 = (~(Iuvmz6[7] & Vg7yx6));
assign Fg7yx6 = (~(Iuvmz6[6] & Dh7yx6));
assign Re7yx6 = (Lh7yx6 & Th7yx6);
assign Th7yx6 = (~(Iuvmz6[5] & Bi7yx6));
assign Lh7yx6 = (~(Iuvmz6[4] & Ji7yx6));
assign Fmq7v6 = (L96yx6 ? Ri7yx6 : Ppwmz6[3]);
assign Ylq7v6 = (F86yx6 ? Trwmz6[3] : Ri7yx6);
assign Ri7yx6 = (~(Zi7yx6 & Hj7yx6));
assign Hj7yx6 = (Pj7yx6 & Xj7yx6);
assign Xj7yx6 = (~(Iuvmz6[7] & Xf7yx6));
assign Pj7yx6 = (Fk7yx6 & Nk7yx6);
assign Nk7yx6 = (~(Iuvmz6[6] & Vg7yx6));
assign Fk7yx6 = (~(Iuvmz6[5] & Dh7yx6));
assign Zi7yx6 = (Vk7yx6 & Dl7yx6);
assign Dl7yx6 = (~(Iuvmz6[4] & Bi7yx6));
assign Vk7yx6 = (~(Iuvmz6[8] & Ji7yx6));
assign Rlq7v6 = (~(Ll7yx6 & Tl7yx6));
assign Tl7yx6 = (~(Ba6yx6 & Cnvmz6[3]));
assign Ll7yx6 = (Bm7yx6 & Jm7yx6);
assign Jm7yx6 = (~(Ppwmz6[3] & By6yx6));
assign Bm7yx6 = (~(Trwmz6[3] & Jy6yx6));
assign Klq7v6 = (Ld6yx6 ? Rm7yx6 : Mgwmz6[3]);
assign Dlq7v6 = (Fc6yx6 ? Qiwmz6[3] : Rm7yx6);
assign Rm7yx6 = (~(Zm7yx6 & Hn7yx6));
assign Hn7yx6 = (Pn7yx6 & Xn7yx6);
assign Xn7yx6 = (~(Iuvmz6[6] & Xf7yx6));
assign Pn7yx6 = (Fo7yx6 & No7yx6);
assign No7yx6 = (~(Iuvmz6[5] & Vg7yx6));
assign Fo7yx6 = (~(Iuvmz6[4] & Dh7yx6));
assign Zm7yx6 = (Vo7yx6 & Dp7yx6);
assign Dp7yx6 = (~(Iuvmz6[8] & Bi7yx6));
assign Vo7yx6 = (~(Iuvmz6[7] & Ji7yx6));
assign Wkq7v6 = (~(Lp7yx6 & Tp7yx6));
assign Tp7yx6 = (~(Be6yx6 & Xovmz6[3]));
assign Lp7yx6 = (Bq7yx6 & Jq7yx6);
assign Jq7yx6 = (~(Mgwmz6[3] & Lt6yx6));
assign Bq7yx6 = (~(Qiwmz6[3] & Tt6yx6));
assign Pkq7v6 = (Lh6yx6 ? Rq7yx6 : J7wmz6[3]);
assign Ikq7v6 = (Fg6yx6 ? N9wmz6[3] : Rq7yx6);
assign Rq7yx6 = (~(Zq7yx6 & Hr7yx6));
assign Hr7yx6 = (Pr7yx6 & Xr7yx6);
assign Xr7yx6 = (~(Iuvmz6[5] & Xf7yx6));
assign Pr7yx6 = (Fs7yx6 & Ns7yx6);
assign Ns7yx6 = (~(Iuvmz6[4] & Vg7yx6));
assign Fs7yx6 = (~(Iuvmz6[8] & Dh7yx6));
assign Zq7yx6 = (Vs7yx6 & Dt7yx6);
assign Dt7yx6 = (~(Iuvmz6[7] & Bi7yx6));
assign Vs7yx6 = (~(Iuvmz6[6] & Ji7yx6));
assign Bkq7v6 = (~(Lt7yx6 & Tt7yx6));
assign Tt7yx6 = (~(Bi6yx6 & Sqvmz6[3]));
assign Lt7yx6 = (Bu7yx6 & Ju7yx6);
assign Ju7yx6 = (~(J7wmz6[3] & Vo6yx6));
assign Bu7yx6 = (~(N9wmz6[3] & Dp6yx6));
assign Ujq7v6 = (Pz5yx6 ? Ru7yx6 : Gyvmz6[3]);
assign Njq7v6 = (Lz4ov6 ? K0wmz6[3] : Ru7yx6);
assign Ru7yx6 = (~(Zu7yx6 & Hv7yx6));
assign Hv7yx6 = (Pv7yx6 & Xv7yx6);
assign Xv7yx6 = (~(Iuvmz6[4] & Xf7yx6));
assign Xf7yx6 = (~(Fw7yx6 & Nw7yx6));
assign Fw7yx6 = (Vw7yx6 & Dx7yx6);
assign Dx7yx6 = (~(Vr5ft6 & P37yx6));
assign Vw7yx6 = (~(X9s7z6[3] & L17yx6));
assign Pv7yx6 = (Lx7yx6 & Tx7yx6);
assign Tx7yx6 = (~(Iuvmz6[8] & Vg7yx6));
assign Vg7yx6 = (~(By7yx6 & Jy7yx6));
assign Jy7yx6 = (Ry7yx6 & Zy7yx6);
assign Zy7yx6 = (Hz7yx6 & Pz7yx6);
assign Pz7yx6 = (~(Tjr7z6[5] & V47yx6));
assign Hz7yx6 = (~(Xz7yx6 & V1s7z6[3]));
assign Ry7yx6 = (F08yx6 & N08yx6);
assign N08yx6 = (~(Gqr7z6[3] & R27yx6));
assign F08yx6 = (~(Cor7z6[3] & N47yx6));
assign By7yx6 = (V08yx6 & D18yx6);
assign D18yx6 = (~(X9s7z6[11] & L17yx6));
assign V08yx6 = (L18yx6 & T18yx6);
assign T18yx6 = (~(P7s7z6[11] & J27yx6));
assign L18yx6 = (~(Wlr7z6[3] & P37yx6));
assign Lx7yx6 = (~(Iuvmz6[7] & Dh7yx6));
assign Dh7yx6 = (~(B28yx6 & J28yx6));
assign J28yx6 = (R28yx6 & Z28yx6);
assign Z28yx6 = (~(Wlr7z6[11] & P37yx6));
assign R28yx6 = (H38yx6 & P38yx6);
assign P38yx6 = (~(Cor7z6[11] & N47yx6));
assign H38yx6 = (~(Gqr7z6[11] & R27yx6));
assign B28yx6 = (X38yx6 & F48yx6);
assign F48yx6 = (~(P7s7z6[19] & J27yx6));
assign X38yx6 = (~(X9s7z6[19] & L17yx6));
assign Zu7yx6 = (N48yx6 & V48yx6);
assign V48yx6 = (~(Iuvmz6[6] & Bi7yx6));
assign Bi7yx6 = (~(D58yx6 & L58yx6));
assign L58yx6 = (T58yx6 & B68yx6);
assign B68yx6 = (~(Wlr7z6[19] & P37yx6));
assign T58yx6 = (J68yx6 & R68yx6);
assign R68yx6 = (~(Cor7z6[19] & N47yx6));
assign J68yx6 = (~(Gqr7z6[19] & R27yx6));
assign D58yx6 = (Z68yx6 & H78yx6);
assign H78yx6 = (~(P7s7z6[27] & J27yx6));
assign Z68yx6 = (~(X9s7z6[27] & L17yx6));
assign N48yx6 = (~(Iuvmz6[5] & Ji7yx6));
assign Ji7yx6 = (~(P78yx6 & X78yx6));
assign X78yx6 = (F88yx6 & N88yx6);
assign N88yx6 = (~(Cor7z6[27] & N47yx6));
assign F88yx6 = (~(Gqr7z6[27] & R27yx6));
assign P78yx6 = (V88yx6 & D98yx6);
assign D98yx6 = (~(Wlr7z6[27] & P37yx6));
assign V88yx6 = (~(X9s7z6[35] & L17yx6));
assign Gjq7v6 = (~(L98yx6 & T98yx6));
assign T98yx6 = (~(Nsvmz6[3] & G05ov6));
assign L98yx6 = (Ba8yx6 & Ja8yx6);
assign Ja8yx6 = (~(Gyvmz6[3] & B15ov6));
assign Ba8yx6 = (~(K0wmz6[3] & I15ov6));
assign Ziq7v6 = (X76yx6 ? Sywmz6[2] : Ra8yx6);
assign Siq7v6 = (R66yx6 ? W0xmz6[2] : Ra8yx6);
assign Ra8yx6 = (~(Za8yx6 & Hb8yx6));
assign Hb8yx6 = (Pb8yx6 & Xb8yx6);
assign Xb8yx6 = (~(Iuvmz6[8] & Fc8yx6));
assign Pb8yx6 = (Nc8yx6 & Vc8yx6);
assign Vc8yx6 = (~(Iuvmz6[7] & Dd8yx6));
assign Nc8yx6 = (~(Iuvmz6[6] & Ld8yx6));
assign Za8yx6 = (Td8yx6 & Be8yx6);
assign Be8yx6 = (~(Iuvmz6[5] & Je8yx6));
assign Td8yx6 = (~(Iuvmz6[4] & Re8yx6));
assign Liq7v6 = (L96yx6 ? Ze8yx6 : Ppwmz6[2]);
assign Eiq7v6 = (F86yx6 ? Trwmz6[2] : Ze8yx6);
assign Ze8yx6 = (~(Hf8yx6 & Pf8yx6));
assign Pf8yx6 = (Xf8yx6 & Fg8yx6);
assign Fg8yx6 = (~(Iuvmz6[7] & Fc8yx6));
assign Xf8yx6 = (Ng8yx6 & Vg8yx6);
assign Vg8yx6 = (~(Iuvmz6[6] & Dd8yx6));
assign Ng8yx6 = (~(Iuvmz6[5] & Ld8yx6));
assign Hf8yx6 = (Dh8yx6 & Lh8yx6);
assign Lh8yx6 = (~(Iuvmz6[4] & Je8yx6));
assign Dh8yx6 = (~(Iuvmz6[8] & Re8yx6));
assign Xhq7v6 = (~(Th8yx6 & Bi8yx6));
assign Bi8yx6 = (~(Ba6yx6 & Cnvmz6[2]));
assign Th8yx6 = (Ji8yx6 & Ri8yx6);
assign Ri8yx6 = (~(Ppwmz6[2] & By6yx6));
assign Ji8yx6 = (~(Trwmz6[2] & Jy6yx6));
assign Qhq7v6 = (Ld6yx6 ? Zi8yx6 : Mgwmz6[2]);
assign Jhq7v6 = (Fc6yx6 ? Qiwmz6[2] : Zi8yx6);
assign Zi8yx6 = (~(Hj8yx6 & Pj8yx6));
assign Pj8yx6 = (Xj8yx6 & Fk8yx6);
assign Fk8yx6 = (~(Iuvmz6[6] & Fc8yx6));
assign Xj8yx6 = (Nk8yx6 & Vk8yx6);
assign Vk8yx6 = (~(Iuvmz6[5] & Dd8yx6));
assign Nk8yx6 = (~(Iuvmz6[4] & Ld8yx6));
assign Hj8yx6 = (Dl8yx6 & Ll8yx6);
assign Ll8yx6 = (~(Iuvmz6[8] & Je8yx6));
assign Dl8yx6 = (~(Iuvmz6[7] & Re8yx6));
assign Chq7v6 = (~(Tl8yx6 & Bm8yx6));
assign Bm8yx6 = (~(Be6yx6 & Xovmz6[2]));
assign Tl8yx6 = (Jm8yx6 & Rm8yx6);
assign Rm8yx6 = (~(Mgwmz6[2] & Lt6yx6));
assign Jm8yx6 = (~(Qiwmz6[2] & Tt6yx6));
assign Vgq7v6 = (Lh6yx6 ? Zm8yx6 : J7wmz6[2]);
assign Ogq7v6 = (Fg6yx6 ? N9wmz6[2] : Zm8yx6);
assign Zm8yx6 = (~(Hn8yx6 & Pn8yx6));
assign Pn8yx6 = (Xn8yx6 & Fo8yx6);
assign Fo8yx6 = (~(Iuvmz6[5] & Fc8yx6));
assign Xn8yx6 = (No8yx6 & Vo8yx6);
assign Vo8yx6 = (~(Iuvmz6[4] & Dd8yx6));
assign No8yx6 = (~(Iuvmz6[8] & Ld8yx6));
assign Hn8yx6 = (Dp8yx6 & Lp8yx6);
assign Lp8yx6 = (~(Iuvmz6[7] & Je8yx6));
assign Dp8yx6 = (~(Iuvmz6[6] & Re8yx6));
assign Hgq7v6 = (~(Tp8yx6 & Bq8yx6));
assign Bq8yx6 = (~(Bi6yx6 & Sqvmz6[2]));
assign Tp8yx6 = (Jq8yx6 & Rq8yx6);
assign Rq8yx6 = (~(J7wmz6[2] & Vo6yx6));
assign Jq8yx6 = (~(N9wmz6[2] & Dp6yx6));
assign Agq7v6 = (Pz5yx6 ? Zq8yx6 : Gyvmz6[2]);
assign Tfq7v6 = (Lz4ov6 ? K0wmz6[2] : Zq8yx6);
assign Zq8yx6 = (~(Hr8yx6 & Pr8yx6));
assign Pr8yx6 = (Xr8yx6 & Fs8yx6);
assign Fs8yx6 = (~(Iuvmz6[4] & Fc8yx6));
assign Fc8yx6 = (~(Ns8yx6 & Vs8yx6));
assign Vs8yx6 = (Dt8yx6 & Dd7yx6);
assign Ns8yx6 = (Lt8yx6 & Tt8yx6);
assign Xr8yx6 = (Bu8yx6 & Ju8yx6);
assign Ju8yx6 = (~(Iuvmz6[8] & Dd8yx6));
assign Dd8yx6 = (~(Ru8yx6 & Zu8yx6));
assign Zu8yx6 = (Hv8yx6 & Pv8yx6);
assign Pv8yx6 = (Xv8yx6 & Fw8yx6);
assign Xv8yx6 = (~(Tjr7z6[4] & V47yx6));
assign Hv8yx6 = (Nw8yx6 & Vw8yx6);
assign Vw8yx6 = (~(Gqr7z6[2] & R27yx6));
assign Nw8yx6 = (~(Cor7z6[2] & N47yx6));
assign Ru8yx6 = (Dx8yx6 & Lx8yx6);
assign Lx8yx6 = (~(Xz7yx6 & V1s7z6[2]));
assign Dx8yx6 = (Tx8yx6 & By8yx6);
assign By8yx6 = (~(X9s7z6[10] & L17yx6));
assign Tx8yx6 = (~(Wlr7z6[2] & P37yx6));
assign Bu8yx6 = (~(Iuvmz6[7] & Ld8yx6));
assign Ld8yx6 = (~(Jy8yx6 & Ry8yx6));
assign Ry8yx6 = (Zy8yx6 & Hz8yx6);
assign Hz8yx6 = (~(Wlr7z6[10] & P37yx6));
assign Zy8yx6 = (Pz8yx6 & Xz8yx6);
assign Xz8yx6 = (~(Cor7z6[10] & N47yx6));
assign Pz8yx6 = (~(Gqr7z6[10] & R27yx6));
assign Jy8yx6 = (F09yx6 & N09yx6);
assign N09yx6 = (~(P7s7z6[18] & J27yx6));
assign F09yx6 = (~(X9s7z6[18] & L17yx6));
assign Hr8yx6 = (V09yx6 & D19yx6);
assign D19yx6 = (~(Iuvmz6[6] & Je8yx6));
assign Je8yx6 = (~(L19yx6 & T19yx6));
assign T19yx6 = (B29yx6 & J29yx6);
assign J29yx6 = (~(Wlr7z6[18] & P37yx6));
assign B29yx6 = (R29yx6 & Z29yx6);
assign Z29yx6 = (~(Cor7z6[18] & N47yx6));
assign R29yx6 = (~(Gqr7z6[18] & R27yx6));
assign L19yx6 = (H39yx6 & P39yx6);
assign P39yx6 = (~(P7s7z6[26] & J27yx6));
assign H39yx6 = (~(X9s7z6[26] & L17yx6));
assign V09yx6 = (~(Iuvmz6[5] & Re8yx6));
assign Re8yx6 = (~(X39yx6 & F49yx6));
assign F49yx6 = (N49yx6 & V49yx6);
assign V49yx6 = (~(Cor7z6[26] & N47yx6));
assign N49yx6 = (~(Gqr7z6[26] & R27yx6));
assign X39yx6 = (D59yx6 & L59yx6);
assign L59yx6 = (~(Wlr7z6[26] & P37yx6));
assign D59yx6 = (~(X9s7z6[34] & L17yx6));
assign Mfq7v6 = (~(T59yx6 & B69yx6));
assign B69yx6 = (~(Nsvmz6[2] & G05ov6));
assign T59yx6 = (J69yx6 & R69yx6);
assign R69yx6 = (~(Gyvmz6[2] & B15ov6));
assign J69yx6 = (~(K0wmz6[2] & I15ov6));
assign Ffq7v6 = (X76yx6 ? Sywmz6[1] : Z69yx6);
assign Yeq7v6 = (R66yx6 ? W0xmz6[1] : Z69yx6);
assign Z69yx6 = (~(H79yx6 & P79yx6));
assign P79yx6 = (X79yx6 & F89yx6);
assign F89yx6 = (~(Iuvmz6[8] & N89yx6));
assign X79yx6 = (V89yx6 & D99yx6);
assign D99yx6 = (~(Iuvmz6[7] & L99yx6));
assign V89yx6 = (~(Iuvmz6[6] & T99yx6));
assign H79yx6 = (Ba9yx6 & Ja9yx6);
assign Ja9yx6 = (~(Iuvmz6[5] & Ra9yx6));
assign Ba9yx6 = (~(Iuvmz6[4] & Za9yx6));
assign Req7v6 = (L96yx6 ? Hb9yx6 : Ppwmz6[1]);
assign Keq7v6 = (F86yx6 ? Trwmz6[1] : Hb9yx6);
assign Hb9yx6 = (~(Pb9yx6 & Xb9yx6));
assign Xb9yx6 = (Fc9yx6 & Nc9yx6);
assign Nc9yx6 = (~(Iuvmz6[7] & N89yx6));
assign Fc9yx6 = (Vc9yx6 & Dd9yx6);
assign Dd9yx6 = (~(Iuvmz6[6] & L99yx6));
assign Vc9yx6 = (~(Iuvmz6[5] & T99yx6));
assign Pb9yx6 = (Ld9yx6 & Td9yx6);
assign Td9yx6 = (~(Iuvmz6[4] & Ra9yx6));
assign Ld9yx6 = (~(Iuvmz6[8] & Za9yx6));
assign Deq7v6 = (~(Be9yx6 & Je9yx6));
assign Je9yx6 = (~(Ba6yx6 & Cnvmz6[1]));
assign Be9yx6 = (Re9yx6 & Ze9yx6);
assign Ze9yx6 = (~(Ppwmz6[1] & By6yx6));
assign Re9yx6 = (~(Trwmz6[1] & Jy6yx6));
assign Wdq7v6 = (Ld6yx6 ? Hf9yx6 : Mgwmz6[1]);
assign Pdq7v6 = (Fc6yx6 ? Qiwmz6[1] : Hf9yx6);
assign Hf9yx6 = (~(Pf9yx6 & Xf9yx6));
assign Xf9yx6 = (Fg9yx6 & Ng9yx6);
assign Ng9yx6 = (~(Iuvmz6[6] & N89yx6));
assign Fg9yx6 = (Vg9yx6 & Dh9yx6);
assign Dh9yx6 = (~(Iuvmz6[5] & L99yx6));
assign Vg9yx6 = (~(Iuvmz6[4] & T99yx6));
assign Pf9yx6 = (Lh9yx6 & Th9yx6);
assign Th9yx6 = (~(Iuvmz6[8] & Ra9yx6));
assign Lh9yx6 = (~(Iuvmz6[7] & Za9yx6));
assign Idq7v6 = (~(Bi9yx6 & Ji9yx6));
assign Ji9yx6 = (~(Be6yx6 & Xovmz6[1]));
assign Bi9yx6 = (Ri9yx6 & Zi9yx6);
assign Zi9yx6 = (~(Mgwmz6[1] & Lt6yx6));
assign Ri9yx6 = (~(Qiwmz6[1] & Tt6yx6));
assign Bdq7v6 = (Lh6yx6 ? Hj9yx6 : J7wmz6[1]);
assign Ucq7v6 = (Fg6yx6 ? N9wmz6[1] : Hj9yx6);
assign Hj9yx6 = (~(Pj9yx6 & Xj9yx6));
assign Xj9yx6 = (Fk9yx6 & Nk9yx6);
assign Nk9yx6 = (~(Iuvmz6[5] & N89yx6));
assign Fk9yx6 = (Vk9yx6 & Dl9yx6);
assign Dl9yx6 = (~(Iuvmz6[4] & L99yx6));
assign Vk9yx6 = (~(Iuvmz6[8] & T99yx6));
assign Pj9yx6 = (Ll9yx6 & Tl9yx6);
assign Tl9yx6 = (~(Iuvmz6[7] & Ra9yx6));
assign Ll9yx6 = (~(Iuvmz6[6] & Za9yx6));
assign Ncq7v6 = (~(Bm9yx6 & Jm9yx6));
assign Jm9yx6 = (~(Bi6yx6 & Sqvmz6[1]));
assign Bm9yx6 = (Rm9yx6 & Zm9yx6);
assign Zm9yx6 = (~(J7wmz6[1] & Vo6yx6));
assign Rm9yx6 = (~(N9wmz6[1] & Dp6yx6));
assign Gcq7v6 = (Pz5yx6 ? Hn9yx6 : Gyvmz6[1]);
assign Zbq7v6 = (Lz4ov6 ? K0wmz6[1] : Hn9yx6);
assign Hn9yx6 = (~(Pn9yx6 & Xn9yx6));
assign Xn9yx6 = (Fo9yx6 & No9yx6);
assign No9yx6 = (~(Iuvmz6[4] & N89yx6));
assign N89yx6 = (~(Vo9yx6 & Dp9yx6));
assign Dp9yx6 = (Lp9yx6 & Dt8yx6);
assign Lp9yx6 = (~(Tp9yx6 | R27yx6));
assign Vo9yx6 = (Bq9yx6 & Tt8yx6);
assign Bq9yx6 = (~(P37yx6 & Jq9yx6));
assign Jq9yx6 = (~(Rq9yx6 ^ Xcr7z6[0]));
assign Fo9yx6 = (Zq9yx6 & Hr9yx6);
assign Hr9yx6 = (~(Iuvmz6[8] & L99yx6));
assign L99yx6 = (~(Pr9yx6 & Xr9yx6));
assign Xr9yx6 = (Fs9yx6 & Ns9yx6);
assign Ns9yx6 = (Vs9yx6 & Dt9yx6);
assign Dt9yx6 = (~(Tjr7z6[3] & V47yx6));
assign Fs9yx6 = (Lt9yx6 & Tt9yx6);
assign Tt9yx6 = (~(Gqr7z6[1] & R27yx6));
assign Lt9yx6 = (~(Xz7yx6 & V1s7z6[1]));
assign Pr9yx6 = (Bu9yx6 & Ju9yx6);
assign Ju9yx6 = (~(X9s7z6[9] & L17yx6));
assign Bu9yx6 = (Ru9yx6 & Zu9yx6);
assign Zu9yx6 = (~(Cor7z6[1] & N47yx6));
assign Ru9yx6 = (~(Wlr7z6[1] & P37yx6));
assign Zq9yx6 = (~(Iuvmz6[7] & T99yx6));
assign T99yx6 = (~(Hv9yx6 & Pv9yx6));
assign Pv9yx6 = (Xv9yx6 & Fw9yx6);
assign Fw9yx6 = (~(Wlr7z6[9] & P37yx6));
assign Xv9yx6 = (Nw9yx6 & Vw9yx6);
assign Vw9yx6 = (~(Cor7z6[9] & N47yx6));
assign Nw9yx6 = (~(Gqr7z6[9] & R27yx6));
assign Hv9yx6 = (Dx9yx6 & Lx9yx6);
assign Lx9yx6 = (~(P7s7z6[17] & J27yx6));
assign Dx9yx6 = (~(X9s7z6[17] & L17yx6));
assign Pn9yx6 = (Tx9yx6 & By9yx6);
assign By9yx6 = (~(Iuvmz6[6] & Ra9yx6));
assign Ra9yx6 = (~(Jy9yx6 & Ry9yx6));
assign Ry9yx6 = (Zy9yx6 & Hz9yx6);
assign Hz9yx6 = (~(Wlr7z6[17] & P37yx6));
assign Zy9yx6 = (Pz9yx6 & Xz9yx6);
assign Xz9yx6 = (~(Cor7z6[17] & N47yx6));
assign Pz9yx6 = (~(Gqr7z6[17] & R27yx6));
assign Jy9yx6 = (F0ayx6 & N0ayx6);
assign N0ayx6 = (~(P7s7z6[25] & J27yx6));
assign F0ayx6 = (~(X9s7z6[25] & L17yx6));
assign Tx9yx6 = (~(Iuvmz6[5] & Za9yx6));
assign Za9yx6 = (~(V0ayx6 & D1ayx6));
assign D1ayx6 = (L1ayx6 & T1ayx6);
assign T1ayx6 = (~(Cor7z6[25] & N47yx6));
assign L1ayx6 = (~(Gqr7z6[25] & R27yx6));
assign V0ayx6 = (B2ayx6 & J2ayx6);
assign J2ayx6 = (~(Wlr7z6[25] & P37yx6));
assign B2ayx6 = (~(X9s7z6[33] & L17yx6));
assign Sbq7v6 = (~(R2ayx6 & Z2ayx6));
assign Z2ayx6 = (~(Nsvmz6[1] & G05ov6));
assign R2ayx6 = (H3ayx6 & P3ayx6);
assign P3ayx6 = (~(Gyvmz6[1] & B15ov6));
assign H3ayx6 = (~(K0wmz6[1] & I15ov6));
assign Lbq7v6 = (X76yx6 ? Sywmz6[0] : X3ayx6);
assign Ebq7v6 = (R66yx6 ? W0xmz6[0] : X3ayx6);
assign X3ayx6 = (~(F4ayx6 & N4ayx6));
assign N4ayx6 = (V4ayx6 & D5ayx6);
assign D5ayx6 = (~(Iuvmz6[8] & L5ayx6));
assign V4ayx6 = (T5ayx6 & B6ayx6);
assign B6ayx6 = (~(Iuvmz6[7] & J6ayx6));
assign T5ayx6 = (~(Iuvmz6[6] & R6ayx6));
assign F4ayx6 = (Z6ayx6 & H7ayx6);
assign H7ayx6 = (~(Iuvmz6[5] & P7ayx6));
assign Z6ayx6 = (~(Iuvmz6[4] & X7ayx6));
assign Xaq7v6 = (L96yx6 ? F8ayx6 : Ppwmz6[0]);
assign Qaq7v6 = (F86yx6 ? Trwmz6[0] : F8ayx6);
assign F8ayx6 = (~(N8ayx6 & V8ayx6));
assign V8ayx6 = (D9ayx6 & L9ayx6);
assign L9ayx6 = (~(Iuvmz6[7] & L5ayx6));
assign D9ayx6 = (T9ayx6 & Baayx6);
assign Baayx6 = (~(Iuvmz6[6] & J6ayx6));
assign T9ayx6 = (~(Iuvmz6[5] & R6ayx6));
assign N8ayx6 = (Jaayx6 & Raayx6);
assign Raayx6 = (~(Iuvmz6[4] & P7ayx6));
assign Jaayx6 = (~(Iuvmz6[8] & X7ayx6));
assign Jaq7v6 = (~(Zaayx6 & Hbayx6));
assign Hbayx6 = (~(Ba6yx6 & Cnvmz6[0]));
assign Zaayx6 = (Pbayx6 & Xbayx6);
assign Xbayx6 = (~(Ppwmz6[0] & By6yx6));
assign Pbayx6 = (~(Trwmz6[0] & Jy6yx6));
assign Caq7v6 = (Ld6yx6 ? Fcayx6 : Mgwmz6[0]);
assign V9q7v6 = (Fc6yx6 ? Qiwmz6[0] : Fcayx6);
assign Fcayx6 = (~(Ncayx6 & Vcayx6));
assign Vcayx6 = (Ddayx6 & Ldayx6);
assign Ldayx6 = (~(Iuvmz6[6] & L5ayx6));
assign Ddayx6 = (Tdayx6 & Beayx6);
assign Beayx6 = (~(Iuvmz6[5] & J6ayx6));
assign Tdayx6 = (~(Iuvmz6[4] & R6ayx6));
assign Ncayx6 = (Jeayx6 & Reayx6);
assign Reayx6 = (~(Iuvmz6[8] & P7ayx6));
assign Jeayx6 = (~(Iuvmz6[7] & X7ayx6));
assign O9q7v6 = (~(Zeayx6 & Hfayx6));
assign Hfayx6 = (~(Be6yx6 & Xovmz6[0]));
assign Zeayx6 = (Pfayx6 & Xfayx6);
assign Xfayx6 = (~(Mgwmz6[0] & Lt6yx6));
assign Pfayx6 = (~(Qiwmz6[0] & Tt6yx6));
assign H9q7v6 = (Lh6yx6 ? Fgayx6 : J7wmz6[0]);
assign A9q7v6 = (Fg6yx6 ? N9wmz6[0] : Fgayx6);
assign Fgayx6 = (~(Ngayx6 & Vgayx6));
assign Vgayx6 = (Dhayx6 & Lhayx6);
assign Lhayx6 = (~(Iuvmz6[5] & L5ayx6));
assign Dhayx6 = (Thayx6 & Biayx6);
assign Biayx6 = (~(Iuvmz6[4] & J6ayx6));
assign Thayx6 = (~(Iuvmz6[8] & R6ayx6));
assign Ngayx6 = (Jiayx6 & Riayx6);
assign Riayx6 = (~(Iuvmz6[7] & P7ayx6));
assign Jiayx6 = (~(Iuvmz6[6] & X7ayx6));
assign T8q7v6 = (~(Ziayx6 & Hjayx6));
assign Hjayx6 = (~(Bi6yx6 & Sqvmz6[0]));
assign Ziayx6 = (Pjayx6 & Xjayx6);
assign Xjayx6 = (~(J7wmz6[0] & Vo6yx6));
assign Pjayx6 = (~(N9wmz6[0] & Dp6yx6));
assign M8q7v6 = (Pz5yx6 ? Fkayx6 : Gyvmz6[0]);
assign F8q7v6 = (Lz4ov6 ? K0wmz6[0] : Fkayx6);
assign Fkayx6 = (~(Nkayx6 & Vkayx6));
assign Vkayx6 = (Dlayx6 & Llayx6);
assign Llayx6 = (~(Iuvmz6[4] & L5ayx6));
assign L5ayx6 = (~(Tlayx6 & Bmayx6));
assign Bmayx6 = (~(Jmayx6 | Rmayx6));
assign Tlayx6 = (Zmayx6 & Lt8yx6);
assign Lt8yx6 = (~(Hnayx6 & Pnayx6));
assign Pnayx6 = (~(Xnayx6 & Ri5yx6));
assign Zmayx6 = (~(X9s7z6[0] & L17yx6));
assign Dlayx6 = (Foayx6 & Noayx6);
assign Noayx6 = (~(Iuvmz6[8] & J6ayx6));
assign J6ayx6 = (~(Voayx6 & Dpayx6));
assign Dpayx6 = (Lpayx6 & Tpayx6);
assign Lpayx6 = (Bqayx6 & Jqayx6);
assign Jqayx6 = (~(Wlr7z6[0] & P37yx6));
assign Bqayx6 = (~(Xz7yx6 & V1s7z6[0]));
assign Voayx6 = (Rqayx6 & Zqayx6);
assign Zqayx6 = (~(Tjr7z6[2] & V47yx6));
assign Rqayx6 = (Hrayx6 & Prayx6);
assign Prayx6 = (~(X9s7z6[8] & L17yx6));
assign Hrayx6 = (~(Cor7z6[0] & N47yx6));
assign Foayx6 = (~(Iuvmz6[7] & R6ayx6));
assign R6ayx6 = (~(Xrayx6 & Fsayx6));
assign Fsayx6 = (Nsayx6 & Vsayx6);
assign Vsayx6 = (~(X9s7z6[16] & L17yx6));
assign Nsayx6 = (Dtayx6 & Ltayx6);
assign Ltayx6 = (~(Wlr7z6[8] & P37yx6));
assign Dtayx6 = (~(Gqr7z6[8] & R27yx6));
assign Xrayx6 = (Ttayx6 & Buayx6);
assign Buayx6 = (~(Tjr7z6[10] & V47yx6));
assign Ttayx6 = (Juayx6 & Ruayx6);
assign Ruayx6 = (~(Cor7z6[8] & N47yx6));
assign Juayx6 = (~(P7s7z6[16] & J27yx6));
assign Nkayx6 = (Zuayx6 & Hvayx6);
assign Hvayx6 = (~(Iuvmz6[6] & P7ayx6));
assign P7ayx6 = (~(Pvayx6 & Xvayx6));
assign Xvayx6 = (Fwayx6 & Nwayx6);
assign Nwayx6 = (~(Wlr7z6[16] & P37yx6));
assign Fwayx6 = (Vwayx6 & Dxayx6);
assign Dxayx6 = (~(Cor7z6[16] & N47yx6));
assign Vwayx6 = (~(Gqr7z6[16] & R27yx6));
assign Pvayx6 = (Lxayx6 & Txayx6);
assign Txayx6 = (~(P7s7z6[24] & J27yx6));
assign Lxayx6 = (~(X9s7z6[24] & L17yx6));
assign Zuayx6 = (~(Iuvmz6[5] & X7ayx6));
assign X7ayx6 = (~(Byayx6 & Jyayx6));
assign Jyayx6 = (Ryayx6 & Zyayx6);
assign Zyayx6 = (~(Cor7z6[24] & N47yx6));
assign Ryayx6 = (~(Gqr7z6[24] & R27yx6));
assign Byayx6 = (Hzayx6 & Pzayx6);
assign Pzayx6 = (~(Wlr7z6[24] & P37yx6));
assign Hzayx6 = (~(X9s7z6[32] & L17yx6));
assign Y7q7v6 = (~(Xzayx6 & F0byx6));
assign F0byx6 = (~(Nsvmz6[0] & G05ov6));
assign Xzayx6 = (N0byx6 & V0byx6);
assign V0byx6 = (~(Gyvmz6[0] & B15ov6));
assign N0byx6 = (~(K0wmz6[0] & I15ov6));
assign R7q7v6 = (D1byx6 & Ixr7z6[1]);
assign D1byx6 = (L1byx6 & Ry5yx6);
assign Ry5yx6 = (~(Zu4yx6 & T1byx6));
assign Zu4yx6 = (!Xv4yx6);
assign L1byx6 = (Alo7x6 | Ixr7z6[0]);
assign Alo7x6 = (~(B2byx6 & U0r7x6));
assign U0r7x6 = (~(Dw4ft6 & Bb9ov6));
assign B2byx6 = (J2byx6 & Z9o7x6);
assign Z9o7x6 = (~(Sk4ft6 & Bb9ov6));
assign J2byx6 = (~(Bb9ov6 & R2byx6));
assign R2byx6 = (M55ft6 | Kg5ft6);
assign Bb9ov6 = (Z2byx6 & O5a7z6);
assign Z2byx6 = (~(A0onv6 | Euget6));
assign K7q7v6 = (~(H3byx6 & P3byx6));
assign P3byx6 = (X3byx6 | Zy3yx6);
assign Zy3yx6 = (!Z24yx6);
assign H3byx6 = (~(Vs27v6 & J24yx6));
assign D7q7v6 = (~(X3byx6 & F4byx6));
assign F4byx6 = (~(Gq37v6 & Fo4yx6));
assign X3byx6 = (N4byx6 & Pr4yx6);
assign Pr4yx6 = (No4yx6 | Dp4yx6);
assign Dp4yx6 = (V4byx6 & L17yx6);
assign N4byx6 = (~(D5byx6 & Xv4yx6));
assign Xv4yx6 = (~(V4byx6 & Hnayx6));
assign W6q7v6 = (!L5byx6);
assign L5byx6 = (Fa5ov6 ? B6byx6 : T5byx6);
assign T5byx6 = (~(J6byx6 & R6byx6));
assign J6byx6 = (~(Ur37v6 | Gq37v6));
assign P6q7v6 = (~(Z6byx6 & H7byx6));
assign H7byx6 = (~(O9xmz6[2] & Ma5ov6));
assign Z6byx6 = (P7byx6 | Fa5ov6);
assign I6q7v6 = (F8byx6 ? X7byx6 : O9xmz6[0]);
assign X7byx6 = (~(N8byx6 & V8byx6));
assign V8byx6 = (~(Vgfnv6 | D9byx6));
assign D9byx6 = (O9xmz6[0] & R6byx6);
assign Vgfnv6 = (~(L9byx6 & T9byx6));
assign T9byx6 = (Babyx6 & Jabyx6);
assign Jabyx6 = (~(TSVALUEB[11] ^ Vcxmz6[11]));
assign Babyx6 = (Rabyx6 & Zabyx6);
assign Zabyx6 = (~(TSVALUEB[12] ^ Vcxmz6[12]));
assign Rabyx6 = (~(TSVALUEB[10] ^ Vcxmz6[10]));
assign L9byx6 = (Hbbyx6 & Pbbyx6);
assign Pbbyx6 = (~(TSVALUEB[8] ^ Vcxmz6[8]));
assign Hbbyx6 = (Xbbyx6 & Fcbyx6);
assign Fcbyx6 = (~(TSVALUEB[9] ^ Vcxmz6[9]));
assign Xbbyx6 = (~(TSVALUEB[7] ^ Vcxmz6[7]));
assign N8byx6 = (Qhfnv6 & Y95ov6);
assign Y95ov6 = (P7byx6 & Xhfnv6);
assign Xhfnv6 = (Ncbyx6 & Vcbyx6);
assign Vcbyx6 = (Ddbyx6 & Ldbyx6);
assign Ldbyx6 = (Tdbyx6 & Bebyx6);
assign Bebyx6 = (~(TSVALUEB[14] ^ Vcxmz6[14]));
assign Tdbyx6 = (~(TSVALUEB[15] ^ Vcxmz6[15]));
assign Ddbyx6 = (Jebyx6 & Rebyx6);
assign Rebyx6 = (~(TSVALUEB[16] ^ Vcxmz6[16]));
assign Jebyx6 = (~(TSVALUEB[17] ^ Vcxmz6[17]));
assign Ncbyx6 = (Zebyx6 & Hfbyx6);
assign Hfbyx6 = (~(TSVALUEB[19] ^ Vcxmz6[19]));
assign Zebyx6 = (Pfbyx6 & Xfbyx6);
assign Xfbyx6 = (~(TSVALUEB[20] ^ Vcxmz6[20]));
assign Pfbyx6 = (~(TSVALUEB[18] ^ Vcxmz6[18]));
assign P7byx6 = (~(Fgbyx6 | X447v6));
assign X447v6 = (~(Sifnv6 & Ngbyx6));
assign Ngbyx6 = (~(P647v6 & Vgbyx6));
assign Vgbyx6 = (~(Ak77z6 & Dhbyx6));
assign Sifnv6 = (Lifnv6 ? Thbyx6 : Lhbyx6);
assign Lifnv6 = (~(R8s7z6[1] | R8s7z6[0]));
assign Thbyx6 = (~(Hr4yx6 & Bibyx6));
assign Bibyx6 = (~(Olfiw6 & Fkfiw6));
assign Lhbyx6 = (Zb1nv6 & Jibyx6);
assign Jibyx6 = (~(Ribyx6 & Fho7v6));
assign Ribyx6 = (Zibyx6 | Fgbyx6);
assign Zb1nv6 = (!Txadt6);
assign Fgbyx6 = (~(Hjbyx6 & Pjbyx6));
assign Pjbyx6 = (Xjbyx6 & Fkbyx6);
assign Fkbyx6 = (~(TSVALUEB[22] ^ Vcxmz6[22]));
assign Xjbyx6 = (Nkbyx6 & Vkbyx6);
assign Vkbyx6 = (~(TSVALUEB[23] ^ Vcxmz6[23]));
assign Nkbyx6 = (~(TSVALUEB[21] ^ Vcxmz6[21]));
assign Hjbyx6 = (Dlbyx6 & Llbyx6);
assign Llbyx6 = (~(TSVALUEB[24] ^ Vcxmz6[24]));
assign Dlbyx6 = (~(TSVALUEB[25] ^ Vcxmz6[25]));
assign Qhfnv6 = (~(TSVALUEB[13] ^ Vcxmz6[13]));
assign B6q7v6 = (~(Tlbyx6 & Bmbyx6));
assign Bmbyx6 = (~(V147v6 & Jmbyx6));
assign Jmbyx6 = (Ma5ov6 | I347v6);
assign Ma5ov6 = (~(Mh5ov6 & F8byx6));
assign Tlbyx6 = (~(Zibyx6 & F8byx6));
assign F8byx6 = (!Fa5ov6);
assign Fa5ov6 = (Rmbyx6 & Zmbyx6);
assign Rmbyx6 = (~(Mh5ov6 & W85ov6));
assign W85ov6 = (~(Hnbyx6 & Pnbyx6));
assign Pnbyx6 = (Xnbyx6 & Fobyx6);
assign Fobyx6 = (~(Sqvmz6[8] & Nk6yx6));
assign Xnbyx6 = (~(Nobyx6 & Vobyx6));
assign Vobyx6 = (~(Dpbyx6 & Lpbyx6));
assign Lpbyx6 = (~(Kms7z6[8] & Kwvmz6[0]));
assign Dpbyx6 = (Tpbyx6 & Bqbyx6);
assign Bqbyx6 = (~(Xovmz6[8] & Kwvmz6[3]));
assign Tpbyx6 = (~(Cnvmz6[8] & Kwvmz6[4]));
assign Hnbyx6 = (Jqbyx6 & Rqbyx6);
assign Rqbyx6 = (Zqbyx6 | Pf5ov6);
assign Jqbyx6 = (~(Nsvmz6[8] & J66yx6));
assign Zibyx6 = (~(Hrbyx6 & Prbyx6));
assign Prbyx6 = (Xrbyx6 & Fsbyx6);
assign Fsbyx6 = (Nsbyx6 & Vsbyx6);
assign Vsbyx6 = (Dtbyx6 & Ltbyx6);
assign Ltbyx6 = (~(TSVALUEB[47] ^ Vcxmz6[47]));
assign Dtbyx6 = (Ttbyx6 & Bubyx6);
assign Bubyx6 = (~(TSVALUEB[43] ^ Vcxmz6[43]));
assign Ttbyx6 = (~(TSVALUEB[45] ^ Vcxmz6[45]));
assign Nsbyx6 = (Jubyx6 & Rubyx6);
assign Rubyx6 = (~(TSVALUEB[40] ^ Vcxmz6[40]));
assign Jubyx6 = (Zubyx6 & Hvbyx6);
assign Hvbyx6 = (~(TSVALUEB[41] ^ Vcxmz6[41]));
assign Zubyx6 = (~(TSVALUEB[44] ^ Vcxmz6[44]));
assign Xrbyx6 = (Pvbyx6 & Xvbyx6);
assign Xvbyx6 = (Fwbyx6 & Nwbyx6);
assign Nwbyx6 = (~(TSVALUEB[34] ^ Vcxmz6[34]));
assign Fwbyx6 = (Vwbyx6 & Dxbyx6);
assign Dxbyx6 = (~(TSVALUEB[36] ^ Vcxmz6[36]));
assign Vwbyx6 = (~(TSVALUEB[38] ^ Vcxmz6[38]));
assign Pvbyx6 = (Lxbyx6 & Txbyx6);
assign Txbyx6 = (~(TSVALUEB[32] ^ Vcxmz6[32]));
assign Lxbyx6 = (~(TSVALUEB[33] ^ Vcxmz6[33]));
assign Hrbyx6 = (Bybyx6 & Jybyx6);
assign Jybyx6 = (Rybyx6 & Zybyx6);
assign Zybyx6 = (Hzbyx6 & Pzbyx6);
assign Pzbyx6 = (~(TSVALUEB[30] ^ Vcxmz6[30]));
assign Hzbyx6 = (Xzbyx6 & F0cyx6);
assign F0cyx6 = (~(TSVALUEB[27] ^ Vcxmz6[27]));
assign Xzbyx6 = (~(TSVALUEB[29] ^ Vcxmz6[29]));
assign Rybyx6 = (N0cyx6 & V0cyx6);
assign V0cyx6 = (~(TSVALUEB[37] ^ Vcxmz6[37]));
assign N0cyx6 = (D1cyx6 & L1cyx6);
assign L1cyx6 = (~(TSVALUEB[39] ^ Vcxmz6[39]));
assign D1cyx6 = (~(TSVALUEB[42] ^ Vcxmz6[42]));
assign Bybyx6 = (T1cyx6 & B2cyx6);
assign B2cyx6 = (J2cyx6 & R2cyx6);
assign R2cyx6 = (~(TSVALUEB[26] ^ Vcxmz6[26]));
assign J2cyx6 = (Z2cyx6 & H3cyx6);
assign H3cyx6 = (~(TSVALUEB[28] ^ Vcxmz6[28]));
assign Z2cyx6 = (~(TSVALUEB[31] ^ Vcxmz6[31]));
assign T1cyx6 = (P3cyx6 & X3cyx6);
assign X3cyx6 = (~(TSVALUEB[35] ^ Vcxmz6[35]));
assign P3cyx6 = (~(TSVALUEB[46] ^ Vcxmz6[46]));
assign U5q7v6 = (Pz5yx6 ? F4cyx6 : Gyvmz6[4]);
assign N5q7v6 = (Lz4ov6 ? K0wmz6[4] : F4cyx6);
assign F4cyx6 = (~(N4cyx6 & V4cyx6));
assign V4cyx6 = (D5cyx6 & L5cyx6);
assign L5cyx6 = (~(Iuvmz6[8] & T5cyx6));
assign D5cyx6 = (B6cyx6 & J6cyx6);
assign J6cyx6 = (~(Iuvmz6[7] & R6cyx6));
assign B6cyx6 = (~(Iuvmz6[6] & Z6cyx6));
assign N4cyx6 = (H7cyx6 & P7cyx6);
assign P7cyx6 = (~(Iuvmz6[5] & X7cyx6));
assign H7cyx6 = (~(Iuvmz6[4] & F8cyx6));
assign G5q7v6 = (~(N8cyx6 & V8cyx6));
assign V8cyx6 = (~(Nsvmz6[4] & G05ov6));
assign N8cyx6 = (D9cyx6 & L9cyx6);
assign L9cyx6 = (~(Gyvmz6[4] & B15ov6));
assign D9cyx6 = (~(K0wmz6[4] & I15ov6));
assign Z4q7v6 = (Lh6yx6 ? T9cyx6 : J7wmz6[4]);
assign S4q7v6 = (Fg6yx6 ? N9wmz6[4] : T9cyx6);
assign T9cyx6 = (~(Bacyx6 & Jacyx6));
assign Jacyx6 = (Racyx6 & Zacyx6);
assign Zacyx6 = (~(Iuvmz6[4] & T5cyx6));
assign Racyx6 = (Hbcyx6 & Pbcyx6);
assign Pbcyx6 = (~(Iuvmz6[8] & R6cyx6));
assign Hbcyx6 = (~(Iuvmz6[7] & Z6cyx6));
assign Bacyx6 = (Xbcyx6 & Fccyx6);
assign Fccyx6 = (~(Iuvmz6[6] & X7cyx6));
assign Xbcyx6 = (~(Iuvmz6[5] & F8cyx6));
assign L4q7v6 = (~(Nccyx6 & Vccyx6));
assign Vccyx6 = (~(Bi6yx6 & Sqvmz6[4]));
assign Nccyx6 = (Ddcyx6 & Ldcyx6);
assign Ldcyx6 = (~(J7wmz6[4] & Vo6yx6));
assign Ddcyx6 = (~(N9wmz6[4] & Dp6yx6));
assign E4q7v6 = (Ld6yx6 ? Tdcyx6 : Mgwmz6[4]);
assign X3q7v6 = (Fc6yx6 ? Qiwmz6[4] : Tdcyx6);
assign Tdcyx6 = (~(Becyx6 & Jecyx6));
assign Jecyx6 = (Recyx6 & Zecyx6);
assign Zecyx6 = (~(Iuvmz6[5] & T5cyx6));
assign Recyx6 = (Hfcyx6 & Pfcyx6);
assign Pfcyx6 = (~(Iuvmz6[4] & R6cyx6));
assign Hfcyx6 = (~(Iuvmz6[8] & Z6cyx6));
assign Becyx6 = (Xfcyx6 & Fgcyx6);
assign Fgcyx6 = (~(Iuvmz6[7] & X7cyx6));
assign Xfcyx6 = (~(Iuvmz6[6] & F8cyx6));
assign Q3q7v6 = (~(Ngcyx6 & Vgcyx6));
assign Vgcyx6 = (~(Be6yx6 & Xovmz6[4]));
assign Ngcyx6 = (Dhcyx6 & Lhcyx6);
assign Lhcyx6 = (~(Mgwmz6[4] & Lt6yx6));
assign Dhcyx6 = (~(Qiwmz6[4] & Tt6yx6));
assign J3q7v6 = (L96yx6 ? Thcyx6 : Ppwmz6[4]);
assign C3q7v6 = (F86yx6 ? Trwmz6[4] : Thcyx6);
assign Thcyx6 = (~(Bicyx6 & Jicyx6));
assign Jicyx6 = (Ricyx6 & Zicyx6);
assign Zicyx6 = (~(Iuvmz6[6] & T5cyx6));
assign Ricyx6 = (Hjcyx6 & Pjcyx6);
assign Pjcyx6 = (~(Iuvmz6[5] & R6cyx6));
assign Hjcyx6 = (~(Iuvmz6[4] & Z6cyx6));
assign Bicyx6 = (Xjcyx6 & Fkcyx6);
assign Fkcyx6 = (~(Iuvmz6[8] & X7cyx6));
assign Xjcyx6 = (~(Iuvmz6[7] & F8cyx6));
assign V2q7v6 = (~(Nkcyx6 & Vkcyx6));
assign Vkcyx6 = (~(Ba6yx6 & Cnvmz6[4]));
assign Nkcyx6 = (Dlcyx6 & Llcyx6);
assign Llcyx6 = (~(Ppwmz6[4] & By6yx6));
assign Dlcyx6 = (~(Trwmz6[4] & Jy6yx6));
assign O2q7v6 = (X76yx6 ? Sywmz6[4] : Tlcyx6);
assign H2q7v6 = (R66yx6 ? W0xmz6[4] : Tlcyx6);
assign Tlcyx6 = (~(Bmcyx6 & Jmcyx6));
assign Jmcyx6 = (Rmcyx6 & Zmcyx6);
assign Zmcyx6 = (~(Iuvmz6[7] & T5cyx6));
assign T5cyx6 = (~(Hncyx6 & Pncyx6));
assign Pncyx6 = (Xncyx6 & Focyx6);
assign Focyx6 = (Nocyx6 & Vocyx6);
assign Vocyx6 = (~(Tjr7z6[6] & V47yx6));
assign Nocyx6 = (~(Xz7yx6 & V1s7z6[4]));
assign Xncyx6 = (Dpcyx6 & Lpcyx6);
assign Lpcyx6 = (~(Gqr7z6[4] & R27yx6));
assign Dpcyx6 = (~(Cor7z6[4] & N47yx6));
assign Hncyx6 = (Tpcyx6 & Bqcyx6);
assign Bqcyx6 = (~(X9s7z6[12] & L17yx6));
assign Tpcyx6 = (Jqcyx6 & Rqcyx6);
assign Rqcyx6 = (~(P7s7z6[12] & J27yx6));
assign Jqcyx6 = (~(Wlr7z6[4] & P37yx6));
assign Rmcyx6 = (Zqcyx6 & Hrcyx6);
assign Hrcyx6 = (~(Iuvmz6[6] & R6cyx6));
assign R6cyx6 = (~(Prcyx6 & Xrcyx6));
assign Xrcyx6 = (Fscyx6 & Nscyx6);
assign Nscyx6 = (~(X9s7z6[20] & L17yx6));
assign Fscyx6 = (Vscyx6 & Dtcyx6);
assign Dtcyx6 = (~(Wlr7z6[12] & P37yx6));
assign Vscyx6 = (~(Gqr7z6[12] & R27yx6));
assign Prcyx6 = (Ltcyx6 & Ttcyx6);
assign Ttcyx6 = (~(Tjr7z6[0] & V47yx6));
assign Ltcyx6 = (Bucyx6 & Jucyx6);
assign Jucyx6 = (~(Cor7z6[12] & N47yx6));
assign Bucyx6 = (~(P7s7z6[20] & J27yx6));
assign Zqcyx6 = (~(Iuvmz6[5] & Z6cyx6));
assign Z6cyx6 = (~(Rucyx6 & Zucyx6));
assign Zucyx6 = (Hvcyx6 & Pvcyx6);
assign Pvcyx6 = (~(Wlr7z6[20] & P37yx6));
assign Hvcyx6 = (Xvcyx6 & Fwcyx6);
assign Fwcyx6 = (~(Cor7z6[20] & N47yx6));
assign Xvcyx6 = (~(Gqr7z6[20] & R27yx6));
assign Rucyx6 = (Nwcyx6 & Vwcyx6);
assign Vwcyx6 = (~(P7s7z6[28] & J27yx6));
assign Nwcyx6 = (~(X9s7z6[28] & L17yx6));
assign Bmcyx6 = (Dxcyx6 & Lxcyx6);
assign Lxcyx6 = (~(Iuvmz6[4] & X7cyx6));
assign X7cyx6 = (~(Txcyx6 & Bycyx6));
assign Bycyx6 = (Jycyx6 & Rycyx6);
assign Rycyx6 = (~(Cor7z6[28] & N47yx6));
assign Jycyx6 = (~(Gqr7z6[28] & R27yx6));
assign Txcyx6 = (Zycyx6 & Hzcyx6);
assign Hzcyx6 = (~(Wlr7z6[28] & P37yx6));
assign Zycyx6 = (~(X9s7z6[36] & L17yx6));
assign Dxcyx6 = (~(Iuvmz6[8] & F8cyx6));
assign F8cyx6 = (~(Pzcyx6 & Xzcyx6));
assign Xzcyx6 = (F0dyx6 & N0dyx6);
assign N0dyx6 = (V0dyx6 | Tpayx6);
assign Tpayx6 = (~(J27yx6 & P7s7z6[8]));
assign F0dyx6 = (D1dyx6 & L1dyx6);
assign D1dyx6 = (~(Dfr7z6[0] & P37yx6));
assign Pzcyx6 = (T1dyx6 & B2dyx6);
assign B2dyx6 = (~(Jhr7z6[0] & N47yx6));
assign T1dyx6 = (J2dyx6 & R2dyx6);
assign R2dyx6 = (~(X9s7z6[4] & L17yx6));
assign J2dyx6 = (~(Nu27v6 & Be7yx6));
assign A2q7v6 = (Pz5yx6 ? Z2dyx6 : Gyvmz6[5]);
assign T1q7v6 = (Lz4ov6 ? K0wmz6[5] : Z2dyx6);
assign Z2dyx6 = (~(H3dyx6 & P3dyx6));
assign P3dyx6 = (X3dyx6 & F4dyx6);
assign F4dyx6 = (~(Iuvmz6[8] & N4dyx6));
assign X3dyx6 = (V4dyx6 & D5dyx6);
assign D5dyx6 = (~(Iuvmz6[7] & L5dyx6));
assign V4dyx6 = (~(Iuvmz6[6] & T5dyx6));
assign H3dyx6 = (B6dyx6 & J6dyx6);
assign J6dyx6 = (~(Iuvmz6[5] & R6dyx6));
assign B6dyx6 = (~(Iuvmz6[4] & Z6dyx6));
assign M1q7v6 = (~(H7dyx6 & P7dyx6));
assign P7dyx6 = (~(Nsvmz6[5] & G05ov6));
assign H7dyx6 = (X7dyx6 & F8dyx6);
assign F8dyx6 = (~(Gyvmz6[5] & B15ov6));
assign X7dyx6 = (~(K0wmz6[5] & I15ov6));
assign F1q7v6 = (Lh6yx6 ? N8dyx6 : J7wmz6[5]);
assign Y0q7v6 = (Fg6yx6 ? N9wmz6[5] : N8dyx6);
assign N8dyx6 = (~(V8dyx6 & D9dyx6));
assign D9dyx6 = (L9dyx6 & T9dyx6);
assign T9dyx6 = (~(Iuvmz6[4] & N4dyx6));
assign L9dyx6 = (Badyx6 & Jadyx6);
assign Jadyx6 = (~(Iuvmz6[8] & L5dyx6));
assign Badyx6 = (~(Iuvmz6[7] & T5dyx6));
assign V8dyx6 = (Radyx6 & Zadyx6);
assign Zadyx6 = (~(Iuvmz6[6] & R6dyx6));
assign Radyx6 = (~(Iuvmz6[5] & Z6dyx6));
assign R0q7v6 = (~(Hbdyx6 & Pbdyx6));
assign Pbdyx6 = (~(Bi6yx6 & Sqvmz6[5]));
assign Hbdyx6 = (Xbdyx6 & Fcdyx6);
assign Fcdyx6 = (~(J7wmz6[5] & Vo6yx6));
assign Xbdyx6 = (~(N9wmz6[5] & Dp6yx6));
assign K0q7v6 = (Ld6yx6 ? Ncdyx6 : Mgwmz6[5]);
assign D0q7v6 = (Fc6yx6 ? Qiwmz6[5] : Ncdyx6);
assign Ncdyx6 = (~(Vcdyx6 & Dddyx6));
assign Dddyx6 = (Lddyx6 & Tddyx6);
assign Tddyx6 = (~(Iuvmz6[5] & N4dyx6));
assign Lddyx6 = (Bedyx6 & Jedyx6);
assign Jedyx6 = (~(Iuvmz6[4] & L5dyx6));
assign Bedyx6 = (~(Iuvmz6[8] & T5dyx6));
assign Vcdyx6 = (Redyx6 & Zedyx6);
assign Zedyx6 = (~(Iuvmz6[7] & R6dyx6));
assign Redyx6 = (~(Iuvmz6[6] & Z6dyx6));
assign Wzp7v6 = (~(Hfdyx6 & Pfdyx6));
assign Pfdyx6 = (~(Be6yx6 & Xovmz6[5]));
assign Hfdyx6 = (Xfdyx6 & Fgdyx6);
assign Fgdyx6 = (~(Mgwmz6[5] & Lt6yx6));
assign Xfdyx6 = (~(Qiwmz6[5] & Tt6yx6));
assign Pzp7v6 = (L96yx6 ? Ngdyx6 : Ppwmz6[5]);
assign Izp7v6 = (F86yx6 ? Trwmz6[5] : Ngdyx6);
assign Ngdyx6 = (~(Vgdyx6 & Dhdyx6));
assign Dhdyx6 = (Lhdyx6 & Thdyx6);
assign Thdyx6 = (~(Iuvmz6[6] & N4dyx6));
assign Lhdyx6 = (Bidyx6 & Jidyx6);
assign Jidyx6 = (~(Iuvmz6[5] & L5dyx6));
assign Bidyx6 = (~(Iuvmz6[4] & T5dyx6));
assign Vgdyx6 = (Ridyx6 & Zidyx6);
assign Zidyx6 = (~(Iuvmz6[8] & R6dyx6));
assign Ridyx6 = (~(Iuvmz6[7] & Z6dyx6));
assign Bzp7v6 = (~(Hjdyx6 & Pjdyx6));
assign Pjdyx6 = (~(Ba6yx6 & Cnvmz6[5]));
assign Hjdyx6 = (Xjdyx6 & Fkdyx6);
assign Fkdyx6 = (~(Ppwmz6[5] & By6yx6));
assign Xjdyx6 = (~(Trwmz6[5] & Jy6yx6));
assign Uyp7v6 = (X76yx6 ? Sywmz6[5] : Nkdyx6);
assign Nyp7v6 = (R66yx6 ? W0xmz6[5] : Nkdyx6);
assign Nkdyx6 = (~(Vkdyx6 & Dldyx6));
assign Dldyx6 = (Lldyx6 & Tldyx6);
assign Tldyx6 = (~(Iuvmz6[7] & N4dyx6));
assign N4dyx6 = (~(Bmdyx6 & Jmdyx6));
assign Jmdyx6 = (Rmdyx6 & Zmdyx6);
assign Zmdyx6 = (Hndyx6 & Pndyx6);
assign Pndyx6 = (~(Tjr7z6[7] & V47yx6));
assign Hndyx6 = (~(Xz7yx6 & V1s7z6[5]));
assign Rmdyx6 = (Xndyx6 & Fodyx6);
assign Fodyx6 = (~(Gqr7z6[5] & R27yx6));
assign Xndyx6 = (~(Cor7z6[5] & N47yx6));
assign Bmdyx6 = (Nodyx6 & Vodyx6);
assign Vodyx6 = (~(X9s7z6[13] & L17yx6));
assign Nodyx6 = (Dpdyx6 & Lpdyx6);
assign Lpdyx6 = (~(P7s7z6[13] & J27yx6));
assign Dpdyx6 = (~(Wlr7z6[5] & P37yx6));
assign Lldyx6 = (Tpdyx6 & Bqdyx6);
assign Bqdyx6 = (~(Iuvmz6[6] & L5dyx6));
assign L5dyx6 = (~(Jqdyx6 & Rqdyx6));
assign Rqdyx6 = (Zqdyx6 & Hrdyx6);
assign Hrdyx6 = (~(X9s7z6[21] & L17yx6));
assign Zqdyx6 = (Prdyx6 & Xrdyx6);
assign Xrdyx6 = (~(Wlr7z6[13] & P37yx6));
assign Prdyx6 = (~(Gqr7z6[13] & R27yx6));
assign Jqdyx6 = (Fsdyx6 & Nsdyx6);
assign Nsdyx6 = (~(Tjr7z6[1] & V47yx6));
assign Fsdyx6 = (Vsdyx6 & Dtdyx6);
assign Dtdyx6 = (~(Cor7z6[13] & N47yx6));
assign Vsdyx6 = (~(P7s7z6[21] & J27yx6));
assign Tpdyx6 = (~(Iuvmz6[5] & T5dyx6));
assign T5dyx6 = (~(Ltdyx6 & Ttdyx6));
assign Ttdyx6 = (Budyx6 & Judyx6);
assign Judyx6 = (~(Wlr7z6[21] & P37yx6));
assign Budyx6 = (Rudyx6 & Zudyx6);
assign Zudyx6 = (~(Cor7z6[21] & N47yx6));
assign Rudyx6 = (~(Gqr7z6[21] & R27yx6));
assign Ltdyx6 = (Hvdyx6 & Pvdyx6);
assign Pvdyx6 = (~(P7s7z6[29] & J27yx6));
assign Hvdyx6 = (~(X9s7z6[29] & L17yx6));
assign Vkdyx6 = (Xvdyx6 & Fwdyx6);
assign Fwdyx6 = (~(Iuvmz6[4] & R6dyx6));
assign R6dyx6 = (~(Nwdyx6 & Vwdyx6));
assign Vwdyx6 = (Dxdyx6 & Lxdyx6);
assign Lxdyx6 = (~(Cor7z6[29] & N47yx6));
assign Dxdyx6 = (~(Gqr7z6[29] & R27yx6));
assign Nwdyx6 = (Txdyx6 & Bydyx6);
assign Bydyx6 = (~(Wlr7z6[29] & P37yx6));
assign Txdyx6 = (~(X9s7z6[37] & L17yx6));
assign Xvdyx6 = (~(Iuvmz6[8] & Z6dyx6));
assign Z6dyx6 = (~(Jydyx6 & Rydyx6));
assign Rydyx6 = (Zydyx6 & Hzdyx6);
assign Hzdyx6 = (~(Jhr7z6[1] & N47yx6));
assign Zydyx6 = (Pzdyx6 & Xzdyx6);
assign Xzdyx6 = (Vs9yx6 | V0dyx6);
assign Vs9yx6 = (~(J27yx6 & P7s7z6[9]));
assign Pzdyx6 = (~(Vs27v6 & Be7yx6));
assign Jydyx6 = (F0eyx6 & N0eyx6);
assign N0eyx6 = (~(X9s7z6[5] & L17yx6));
assign F0eyx6 = (~(Dfr7z6[1] & P37yx6));
assign Gyp7v6 = (Pz5yx6 ? V0eyx6 : Gyvmz6[6]);
assign Zxp7v6 = (Lz4ov6 ? K0wmz6[6] : V0eyx6);
assign V0eyx6 = (~(D1eyx6 & L1eyx6));
assign L1eyx6 = (T1eyx6 & B2eyx6);
assign B2eyx6 = (~(Iuvmz6[8] & J2eyx6));
assign T1eyx6 = (R2eyx6 & Z2eyx6);
assign Z2eyx6 = (~(Iuvmz6[7] & H3eyx6));
assign R2eyx6 = (~(Iuvmz6[6] & P3eyx6));
assign D1eyx6 = (X3eyx6 & F4eyx6);
assign F4eyx6 = (~(Iuvmz6[5] & N4eyx6));
assign X3eyx6 = (~(Iuvmz6[4] & V4eyx6));
assign Sxp7v6 = (~(D5eyx6 & L5eyx6));
assign L5eyx6 = (~(Nsvmz6[6] & G05ov6));
assign D5eyx6 = (T5eyx6 & B6eyx6);
assign B6eyx6 = (~(Gyvmz6[6] & B15ov6));
assign T5eyx6 = (~(K0wmz6[6] & I15ov6));
assign Lxp7v6 = (Lh6yx6 ? J6eyx6 : J7wmz6[6]);
assign Exp7v6 = (Fg6yx6 ? N9wmz6[6] : J6eyx6);
assign J6eyx6 = (~(R6eyx6 & Z6eyx6));
assign Z6eyx6 = (H7eyx6 & P7eyx6);
assign P7eyx6 = (~(Iuvmz6[4] & J2eyx6));
assign H7eyx6 = (X7eyx6 & F8eyx6);
assign F8eyx6 = (~(Iuvmz6[8] & H3eyx6));
assign X7eyx6 = (~(Iuvmz6[7] & P3eyx6));
assign R6eyx6 = (N8eyx6 & V8eyx6);
assign V8eyx6 = (~(Iuvmz6[6] & N4eyx6));
assign N8eyx6 = (~(Iuvmz6[5] & V4eyx6));
assign Xwp7v6 = (~(D9eyx6 & L9eyx6));
assign L9eyx6 = (~(Bi6yx6 & Sqvmz6[6]));
assign D9eyx6 = (T9eyx6 & Baeyx6);
assign Baeyx6 = (~(J7wmz6[6] & Vo6yx6));
assign T9eyx6 = (~(N9wmz6[6] & Dp6yx6));
assign Qwp7v6 = (Ld6yx6 ? Jaeyx6 : Mgwmz6[6]);
assign Jwp7v6 = (Fc6yx6 ? Qiwmz6[6] : Jaeyx6);
assign Jaeyx6 = (~(Raeyx6 & Zaeyx6));
assign Zaeyx6 = (Hbeyx6 & Pbeyx6);
assign Pbeyx6 = (~(Iuvmz6[5] & J2eyx6));
assign Hbeyx6 = (Xbeyx6 & Fceyx6);
assign Fceyx6 = (~(Iuvmz6[4] & H3eyx6));
assign Xbeyx6 = (~(Iuvmz6[8] & P3eyx6));
assign Raeyx6 = (Nceyx6 & Vceyx6);
assign Vceyx6 = (~(Iuvmz6[7] & N4eyx6));
assign Nceyx6 = (~(Iuvmz6[6] & V4eyx6));
assign Cwp7v6 = (~(Ddeyx6 & Ldeyx6));
assign Ldeyx6 = (~(Be6yx6 & Xovmz6[6]));
assign Ddeyx6 = (Tdeyx6 & Beeyx6);
assign Beeyx6 = (~(Mgwmz6[6] & Lt6yx6));
assign Tdeyx6 = (~(Qiwmz6[6] & Tt6yx6));
assign Vvp7v6 = (L96yx6 ? Jeeyx6 : Ppwmz6[6]);
assign Ovp7v6 = (F86yx6 ? Trwmz6[6] : Jeeyx6);
assign Jeeyx6 = (~(Reeyx6 & Zeeyx6));
assign Zeeyx6 = (Hfeyx6 & Pfeyx6);
assign Pfeyx6 = (~(Iuvmz6[6] & J2eyx6));
assign Hfeyx6 = (Xfeyx6 & Fgeyx6);
assign Fgeyx6 = (~(Iuvmz6[5] & H3eyx6));
assign Xfeyx6 = (~(Iuvmz6[4] & P3eyx6));
assign Reeyx6 = (Ngeyx6 & Vgeyx6);
assign Vgeyx6 = (~(Iuvmz6[8] & N4eyx6));
assign Ngeyx6 = (~(Iuvmz6[7] & V4eyx6));
assign Hvp7v6 = (~(Dheyx6 & Lheyx6));
assign Lheyx6 = (~(Ba6yx6 & Cnvmz6[6]));
assign Dheyx6 = (Theyx6 & Bieyx6);
assign Bieyx6 = (~(Ppwmz6[6] & By6yx6));
assign Theyx6 = (~(Trwmz6[6] & Jy6yx6));
assign Avp7v6 = (X76yx6 ? Sywmz6[6] : Jieyx6);
assign Tup7v6 = (R66yx6 ? W0xmz6[6] : Jieyx6);
assign Jieyx6 = (~(Rieyx6 & Zieyx6));
assign Zieyx6 = (Hjeyx6 & Pjeyx6);
assign Pjeyx6 = (~(Iuvmz6[7] & J2eyx6));
assign J2eyx6 = (~(Xjeyx6 & Fkeyx6));
assign Fkeyx6 = (Nkeyx6 & Vkeyx6);
assign Vkeyx6 = (~(X9s7z6[14] & L17yx6));
assign Nkeyx6 = (Dleyx6 & Lleyx6);
assign Lleyx6 = (~(Wlr7z6[6] & P37yx6));
assign Dleyx6 = (~(Gqr7z6[6] & R27yx6));
assign Xjeyx6 = (Tleyx6 & Bmeyx6);
assign Bmeyx6 = (~(Tjr7z6[8] & V47yx6));
assign Tleyx6 = (Jmeyx6 & Rmeyx6);
assign Rmeyx6 = (~(Cor7z6[6] & N47yx6));
assign Jmeyx6 = (~(P7s7z6[14] & J27yx6));
assign Hjeyx6 = (Zmeyx6 & Hneyx6);
assign Hneyx6 = (~(Iuvmz6[6] & H3eyx6));
assign H3eyx6 = (~(Pneyx6 & Xneyx6));
assign Xneyx6 = (Foeyx6 & Noeyx6);
assign Noeyx6 = (~(Wlr7z6[14] & P37yx6));
assign Foeyx6 = (Voeyx6 & Dpeyx6);
assign Dpeyx6 = (~(Cor7z6[14] & N47yx6));
assign Voeyx6 = (~(Gqr7z6[14] & R27yx6));
assign Pneyx6 = (Lpeyx6 & Tpeyx6);
assign Tpeyx6 = (~(P7s7z6[22] & J27yx6));
assign Lpeyx6 = (~(X9s7z6[22] & L17yx6));
assign Zmeyx6 = (~(Iuvmz6[5] & P3eyx6));
assign P3eyx6 = (~(Bqeyx6 & Jqeyx6));
assign Jqeyx6 = (Rqeyx6 & Zqeyx6);
assign Zqeyx6 = (~(Wlr7z6[22] & P37yx6));
assign Rqeyx6 = (Hreyx6 & Preyx6);
assign Preyx6 = (~(Cor7z6[22] & N47yx6));
assign Hreyx6 = (~(Gqr7z6[22] & R27yx6));
assign Bqeyx6 = (Xreyx6 & Fseyx6);
assign Fseyx6 = (~(P7s7z6[30] & J27yx6));
assign Xreyx6 = (~(X9s7z6[30] & L17yx6));
assign Rieyx6 = (Nseyx6 & Vseyx6);
assign Vseyx6 = (~(Iuvmz6[4] & N4eyx6));
assign N4eyx6 = (~(Dteyx6 & Lteyx6));
assign Lteyx6 = (Tteyx6 & Bueyx6);
assign Bueyx6 = (~(Cor7z6[30] & N47yx6));
assign Tteyx6 = (~(Gqr7z6[30] & R27yx6));
assign Dteyx6 = (Jueyx6 & Rueyx6);
assign Rueyx6 = (~(Wlr7z6[30] & P37yx6));
assign Jueyx6 = (~(X9s7z6[38] & L17yx6));
assign Nseyx6 = (~(Iuvmz6[8] & V4eyx6));
assign V4eyx6 = (~(Zueyx6 & Hveyx6));
assign Hveyx6 = (~(Be7yx6 | N47yx6));
assign Zueyx6 = (Pveyx6 & Fw8yx6);
assign Fw8yx6 = (~(J27yx6 & P7s7z6[10]));
assign Pveyx6 = (~(X9s7z6[6] & L17yx6));
assign Mup7v6 = (J24yx6 & Xveyx6);
assign Xveyx6 = (Y26ft6 | Fweyx6);
assign Fweyx6 = (Nweyx6 & Vweyx6);
assign Vweyx6 = (Dxeyx6 & Lxeyx6);
assign Lxeyx6 = (Txeyx6 & P7s7z6[16]);
assign Txeyx6 = (R64yx6 & P7s7z6[8]);
assign R64yx6 = (Byeyx6 & Jyeyx6);
assign Jyeyx6 = (Ryeyx6 & Zyeyx6);
assign Zyeyx6 = (Hzeyx6 & Pzeyx6);
assign Pzeyx6 = (P7s7z6[9] & P7s7z6[10]);
assign Hzeyx6 = (P7s7z6[30] & Bm4yx6);
assign Bm4yx6 = (~(Xz3yx6 | Xzeyx6));
assign Xzeyx6 = (F0fyx6 & N0fyx6);
assign N0fyx6 = (~(V0fyx6 & Zq3yx6));
assign Zq3yx6 = (D1fyx6 ^ Vis7z6[5]);
assign D1fyx6 = (~(Vis7z6[4] & Lt3yx6));
assign V0fyx6 = (Vis7z6[4] & Lt3yx6);
assign Lt3yx6 = (~(Tx3yx6 | Dt3yx6));
assign Dt3yx6 = (!Vis7z6[3]);
assign Tx3yx6 = (~(L1fyx6 & Vis7z6[1]));
assign L1fyx6 = (Vis7z6[0] & Vis7z6[2]);
assign F0fyx6 = (~(Hz3yx6 | Ry3yx6));
assign Ry3yx6 = (T1fyx6 & B2fyx6);
assign B2fyx6 = (J2fyx6 & R2fyx6);
assign R2fyx6 = (~(Zm37v6 & Z2fyx6));
assign Z2fyx6 = (~(Vis7z6[3] & Vis7z6[2]));
assign J2fyx6 = (~(Vis7z6[4] | Vis7z6[5]));
assign T1fyx6 = (~(H3fyx6 | P3fyx6));
assign P3fyx6 = (Zm37v6 ? H56ft6 : X3fyx6);
assign X3fyx6 = (Vis7z6[2] | Vis7z6[3]);
assign H3fyx6 = (~(Vis7z6[1] & Vis7z6[0]));
assign Hz3yx6 = (~(Zm37v6 | H56ft6));
assign Xz3yx6 = (~(We6ft6 ^ Qb6ft6));
assign Ryeyx6 = (F4fyx6 & P7s7z6[13]);
assign F4fyx6 = (P7s7z6[12] & P7s7z6[11]);
assign Byeyx6 = (N4fyx6 & V4fyx6);
assign V4fyx6 = (D5fyx6 & P7s7z6[25]);
assign D5fyx6 = (P7s7z6[19] & P7s7z6[14]);
assign N4fyx6 = (L5fyx6 & P7s7z6[29]);
assign L5fyx6 = (P7s7z6[28] & P7s7z6[27]);
assign Dxeyx6 = (P7s7z6[18] & P7s7z6[17]);
assign Nweyx6 = (T5fyx6 & B6fyx6);
assign B6fyx6 = (J6fyx6 & P7s7z6[22]);
assign J6fyx6 = (P7s7z6[21] & P7s7z6[20]);
assign T5fyx6 = (P7s7z6[26] & P7s7z6[24]);
assign J24yx6 = (Hn4yx6 & Z24yx6);
assign Z24yx6 = (Id6ft6 | Ak6ft6);
assign Hn4yx6 = (~(V4byx6 & J27yx6));
assign Fup7v6 = (Pz5yx6 ? R6fyx6 : Gyvmz6[8]);
assign Pz5yx6 = (~(Hz5yx6 | Z6fyx6));
assign Ytp7v6 = (Lz4ov6 ? K0wmz6[8] : R6fyx6);
assign Lz4ov6 = (~(H7fyx6 & Z6fyx6));
assign H7fyx6 = (!Hz5yx6);
assign Hz5yx6 = (~(P7fyx6 & X7fyx6));
assign R6fyx6 = (Iuvmz6[4] & F8fyx6);
assign Rtp7v6 = (~(N8fyx6 & V8fyx6));
assign V8fyx6 = (~(Nsvmz6[8] & G05ov6));
assign N8fyx6 = (D9fyx6 & L9fyx6);
assign L9fyx6 = (~(Gyvmz6[8] & B15ov6));
assign B15ov6 = (~(V46yx6 | G05ov6));
assign V46yx6 = (!O2wmz6[0]);
assign D9fyx6 = (~(K0wmz6[8] & I15ov6));
assign I15ov6 = (~(G05ov6 | O2wmz6[0]));
assign G05ov6 = (!F46yx6);
assign F46yx6 = (~(T9fyx6 & Xj3yx6));
assign Xj3yx6 = (!J66yx6);
assign J66yx6 = (Kwvmz6[1] & Nobyx6);
assign T9fyx6 = (~(D047v6 & N46yx6));
assign N46yx6 = (~(Bafyx6 & Jafyx6));
assign Bafyx6 = (~(O2wmz6[1] ^ Y4wmz6[1]));
assign Ktp7v6 = (Lh6yx6 ? Rafyx6 : J7wmz6[8]);
assign Lh6yx6 = (Dh6yx6 & Bewmz6[0]);
assign Dtp7v6 = (Fg6yx6 ? N9wmz6[8] : Rafyx6);
assign Fg6yx6 = (~(Dh6yx6 & Vg6yx6));
assign Dh6yx6 = (P7fyx6 & Zafyx6);
assign Rafyx6 = (Iuvmz6[5] & F8fyx6);
assign Wsp7v6 = (~(Hbfyx6 & Pbfyx6));
assign Pbfyx6 = (~(Bi6yx6 & Sqvmz6[8]));
assign Hbfyx6 = (Xbfyx6 & Fcfyx6);
assign Fcfyx6 = (~(J7wmz6[8] & Vo6yx6));
assign Vo6yx6 = (~(Zi6yx6 | Bi6yx6));
assign Zi6yx6 = (!Rbwmz6[0]);
assign Xbfyx6 = (~(N9wmz6[8] & Dp6yx6));
assign Dp6yx6 = (~(Bi6yx6 | Rbwmz6[0]));
assign Bi6yx6 = (Xj6yx6 & Nk3yx6);
assign Nk3yx6 = (!Nk6yx6);
assign Nk6yx6 = (Kwvmz6[2] & Nobyx6);
assign Xj6yx6 = (~(Ly37v6 & Ji6yx6));
assign Ji6yx6 = (~(Ncfyx6 & Vcfyx6));
assign Ncfyx6 = (~(Rbwmz6[1] ^ Bewmz6[1]));
assign Psp7v6 = (Ld6yx6 ? Ddfyx6 : Mgwmz6[8]);
assign Ld6yx6 = (Dd6yx6 & Enwmz6[0]);
assign Isp7v6 = (Fc6yx6 ? Qiwmz6[8] : Ddfyx6);
assign Fc6yx6 = (~(Dd6yx6 & Vc6yx6));
assign Dd6yx6 = (P7fyx6 & Ldfyx6);
assign Ddfyx6 = (Iuvmz6[6] & F8fyx6);
assign Bsp7v6 = (~(Tdfyx6 & Befyx6));
assign Befyx6 = (~(Be6yx6 & Xovmz6[8]));
assign Tdfyx6 = (Jefyx6 & Refyx6);
assign Refyx6 = (~(Mgwmz6[8] & Lt6yx6));
assign Lt6yx6 = (~(Re6yx6 | Be6yx6));
assign Re6yx6 = (!Ukwmz6[0]);
assign Jefyx6 = (~(Qiwmz6[8] & Tt6yx6));
assign Tt6yx6 = (~(Be6yx6 | Ukwmz6[0]));
assign Be6yx6 = (Pf6yx6 & Dl3yx6);
assign Dl3yx6 = (~(Kwvmz6[3] & Nobyx6));
assign Pf6yx6 = (Zefyx6 | Td6yx6);
assign Td6yx6 = (Hffyx6 & Pffyx6);
assign Hffyx6 = (~(Ukwmz6[1] ^ Enwmz6[1]));
assign Zefyx6 = (!Tw37v6);
assign Urp7v6 = (L96yx6 ? Xffyx6 : Ppwmz6[8]);
assign L96yx6 = (D96yx6 & Hwwmz6[0]);
assign Nrp7v6 = (F86yx6 ? Trwmz6[8] : Xffyx6);
assign F86yx6 = (~(D96yx6 & V86yx6));
assign D96yx6 = (P7fyx6 & Fgfyx6);
assign Xffyx6 = (Iuvmz6[7] & F8fyx6);
assign Grp7v6 = (~(Ngfyx6 & Vgfyx6));
assign Vgfyx6 = (~(Ba6yx6 & Cnvmz6[8]));
assign Ngfyx6 = (Dhfyx6 & Lhfyx6);
assign Lhfyx6 = (~(Ppwmz6[8] & By6yx6));
assign By6yx6 = (~(Ra6yx6 | Ba6yx6));
assign Ra6yx6 = (!Xtwmz6[0]);
assign Dhfyx6 = (~(Trwmz6[8] & Jy6yx6));
assign Jy6yx6 = (~(Ba6yx6 | Xtwmz6[0]));
assign Ba6yx6 = (Pb6yx6 & Tl3yx6);
assign Tl3yx6 = (~(Kwvmz6[4] & Nobyx6));
assign Pb6yx6 = (Thfyx6 | T96yx6);
assign T96yx6 = (Bifyx6 & Jifyx6);
assign Bifyx6 = (~(Xtwmz6[1] ^ Hwwmz6[1]));
assign Zqp7v6 = (X76yx6 ? Sywmz6[8] : Rifyx6);
assign X76yx6 = (~(P76yx6 & K5xmz6[0]));
assign Sqp7v6 = (R66yx6 ? W0xmz6[8] : Rifyx6);
assign R66yx6 = (~(P76yx6 & H76yx6));
assign P76yx6 = (P7fyx6 & Zifyx6);
assign Rifyx6 = (Iuvmz6[8] & F8fyx6);
assign F8fyx6 = (~(Hjfyx6 & Pjfyx6));
assign Pjfyx6 = (Xjfyx6 & Fkfyx6);
assign Fkfyx6 = (Nkfyx6 & Ld7yx6);
assign Nkfyx6 = (~(Hsr7z6[0] & Vkfyx6));
assign Xjfyx6 = (Dlfyx6 & Llfyx6);
assign Llfyx6 = (~(Xz7yx6 & C4s7z6[0]));
assign Dlfyx6 = (~(Uur7z6[0] & V47yx6));
assign Hjfyx6 = (Tlfyx6 & Bmfyx6);
assign Bmfyx6 = (Jmfyx6 & Rmfyx6);
assign Rmfyx6 = (~(Y26ft6 & J27yx6));
assign Jmfyx6 = (~(Ixr7z6[0] & P37yx6));
assign Tlfyx6 = (Zmfyx6 & Hnfyx6);
assign Hnfyx6 = (~(Tl6ft6 & L17yx6));
assign Zmfyx6 = (~(Nw5ft6 & N47yx6));
assign Lqp7v6 = (~(Pnfyx6 & Xnfyx6));
assign Xnfyx6 = (~(No3yx6 & Kms7z6[0]));
assign Pnfyx6 = (Fofyx6 & Nofyx6);
assign Nofyx6 = (~(Vofyx6 & Sywmz6[0]));
assign Fofyx6 = (~(Dpfyx6 & W0xmz6[0]));
assign Eqp7v6 = (D25ov6 ? V7xmz6[0] : Lpfyx6);
assign Xpp7v6 = (~(Tpfyx6 & Bqfyx6));
assign Bqfyx6 = (~(No3yx6 & Kms7z6[8]));
assign Tpfyx6 = (Jqfyx6 & Rqfyx6);
assign Rqfyx6 = (~(Vofyx6 & Sywmz6[8]));
assign Jqfyx6 = (~(Dpfyx6 & W0xmz6[8]));
assign Qpp7v6 = (~(Zqfyx6 & Hrfyx6));
assign Hrfyx6 = (~(No3yx6 & Kms7z6[7]));
assign Zqfyx6 = (Prfyx6 & Xrfyx6);
assign Xrfyx6 = (~(Vofyx6 & Sywmz6[7]));
assign Prfyx6 = (~(Dpfyx6 & W0xmz6[7]));
assign Jpp7v6 = (~(Fsfyx6 & Nsfyx6));
assign Nsfyx6 = (~(No3yx6 & Kms7z6[6]));
assign Fsfyx6 = (Vsfyx6 & Dtfyx6);
assign Dtfyx6 = (~(Vofyx6 & Sywmz6[6]));
assign Vsfyx6 = (~(Dpfyx6 & W0xmz6[6]));
assign Cpp7v6 = (D25ov6 ? V7xmz6[6] : Ltfyx6);
assign Vop7v6 = (~(Ttfyx6 & Bufyx6));
assign Bufyx6 = (~(No3yx6 & Kms7z6[5]));
assign Ttfyx6 = (Jufyx6 & Rufyx6);
assign Rufyx6 = (~(Vofyx6 & Sywmz6[5]));
assign Jufyx6 = (~(Dpfyx6 & W0xmz6[5]));
assign Oop7v6 = (D25ov6 ? V7xmz6[5] : Zufyx6);
assign Hop7v6 = (~(Hvfyx6 & Pvfyx6));
assign Pvfyx6 = (~(No3yx6 & Kms7z6[4]));
assign Hvfyx6 = (Xvfyx6 & Fwfyx6);
assign Fwfyx6 = (~(Vofyx6 & Sywmz6[4]));
assign Xvfyx6 = (~(Dpfyx6 & W0xmz6[4]));
assign Aop7v6 = (D25ov6 ? V7xmz6[4] : Nwfyx6);
assign Tnp7v6 = (~(Vwfyx6 & Dxfyx6));
assign Dxfyx6 = (~(No3yx6 & Kms7z6[3]));
assign Vwfyx6 = (Lxfyx6 & Txfyx6);
assign Txfyx6 = (~(Vofyx6 & Sywmz6[3]));
assign Lxfyx6 = (~(Dpfyx6 & W0xmz6[3]));
assign Mnp7v6 = (D25ov6 ? V7xmz6[3] : Byfyx6);
assign Fnp7v6 = (~(Jyfyx6 & Ryfyx6));
assign Ryfyx6 = (~(No3yx6 & Kms7z6[2]));
assign Jyfyx6 = (Zyfyx6 & Hzfyx6);
assign Hzfyx6 = (~(Vofyx6 & Sywmz6[2]));
assign Zyfyx6 = (~(Dpfyx6 & W0xmz6[2]));
assign Ymp7v6 = (D25ov6 ? V7xmz6[2] : Pzfyx6);
assign Rmp7v6 = (~(Xzfyx6 & F0gyx6));
assign F0gyx6 = (~(No3yx6 & Kms7z6[1]));
assign Xzfyx6 = (N0gyx6 & V0gyx6);
assign V0gyx6 = (~(Vofyx6 & Sywmz6[1]));
assign Vofyx6 = (~(Rm3yx6 | No3yx6));
assign Rm3yx6 = (!A3xmz6[0]);
assign N0gyx6 = (~(Dpfyx6 & W0xmz6[1]));
assign Dpfyx6 = (~(No3yx6 | A3xmz6[0]));
assign No3yx6 = (Pn3yx6 & Zi3yx6);
assign Zi3yx6 = (~(Kwvmz6[0] & Nobyx6));
assign Nobyx6 = (!Pj3yx6);
assign Pn3yx6 = (D1gyx6 | Fo3yx6);
assign Fo3yx6 = (L1gyx6 & T1gyx6);
assign L1gyx6 = (~(A3xmz6[1] ^ K5xmz6[1]));
assign Kmp7v6 = (D25ov6 ? V7xmz6[1] : B2gyx6);
assign D25ov6 = (K25ov6 & J2gyx6);
assign J2gyx6 = (~(R2gyx6 & La6ft6));
assign R2gyx6 = (~(Zqbyx6 | Z2gyx6));
assign Z2gyx6 = (H3gyx6 & P3gyx6);
assign P3gyx6 = (R6byx6 & X3gyx6);
assign H3gyx6 = (~(F4gyx6 | N4gyx6));
assign K25ov6 = (V4gyx6 & D5gyx6);
assign D5gyx6 = (~(N4gyx6 & L5gyx6));
assign L5gyx6 = (B6byx6 | O9xmz6[2]);
assign N4gyx6 = (T5gyx6 & F35ov6);
assign F35ov6 = (B6gyx6 & J6gyx6);
assign J6gyx6 = (R6gyx6 & S65ov6);
assign S65ov6 = (~(Fbxmz6[2] & Z6gyx6));
assign R6gyx6 = (~(B85ov6 & H7gyx6));
assign B6gyx6 = (P7gyx6 & X7gyx6);
assign X7gyx6 = (~(F8gyx6 & N8gyx6));
assign N8gyx6 = (~(V8gyx6 | D9gyx6));
assign V8gyx6 = (Byfyx6 | X3gyx6);
assign F8gyx6 = (~(L9gyx6 | Lpfyx6));
assign L9gyx6 = (Pzfyx6 | B2gyx6);
assign T5gyx6 = (~(D95ov6 | I85ov6));
assign I85ov6 = (T9gyx6 & Bagyx6);
assign Bagyx6 = (Jagyx6 & Ragyx6);
assign Jagyx6 = (!B85ov6);
assign T9gyx6 = (Zagyx6 & Hbgyx6);
assign Zagyx6 = (~(Fbxmz6[1] & Fbxmz6[3]));
assign D95ov6 = (~(Pbgyx6 & Xbgyx6));
assign Xbgyx6 = (N75ov6 & Ragyx6);
assign N75ov6 = (~(Fcgyx6 & Fbxmz6[2]));
assign Fcgyx6 = (Ncgyx6 & Vcgyx6);
assign Pbgyx6 = (P7gyx6 & Ddgyx6);
assign Ddgyx6 = (~(Pf5ov6 & Ldgyx6));
assign Ldgyx6 = (~(Tdgyx6 & Begyx6));
assign Begyx6 = (~(Jegyx6 | B2gyx6));
assign Jegyx6 = (D9gyx6 | Byfyx6);
assign Byfyx6 = (~(Regyx6 & Zegyx6));
assign Zegyx6 = (Hfgyx6 & Pfgyx6);
assign Pfgyx6 = (~(Sqvmz6[3] & Kwvmz6[2]));
assign Hfgyx6 = (Xfgyx6 & Fggyx6);
assign Fggyx6 = (~(Nsvmz6[3] & Kwvmz6[1]));
assign Xfgyx6 = (~(Xovmz6[3] & Kwvmz6[3]));
assign Regyx6 = (Nggyx6 & Vggyx6);
assign Vggyx6 = (~(Cnvmz6[3] & Kwvmz6[4]));
assign Nggyx6 = (~(Kms7z6[3] & Kwvmz6[0]));
assign D9gyx6 = (~(Dhgyx6 & Lhgyx6));
assign Lhgyx6 = (Thgyx6 & P15ov6);
assign P15ov6 = (~(Bigyx6 & Jigyx6));
assign Jigyx6 = (Rigyx6 & Zigyx6);
assign Zigyx6 = (~(Xovmz6[7] & Kwvmz6[3]));
assign Rigyx6 = (Hjgyx6 & Pjgyx6);
assign Pjgyx6 = (~(Nsvmz6[7] & Kwvmz6[1]));
assign Hjgyx6 = (~(Sqvmz6[7] & Kwvmz6[2]));
assign Bigyx6 = (Xjgyx6 & Fkgyx6);
assign Fkgyx6 = (~(Cnvmz6[7] & Kwvmz6[4]));
assign Xjgyx6 = (~(Kms7z6[7] & Kwvmz6[0]));
assign Thgyx6 = (!Ltfyx6);
assign Ltfyx6 = (~(Nkgyx6 & Vkgyx6));
assign Vkgyx6 = (Dlgyx6 & Llgyx6);
assign Llgyx6 = (~(Xovmz6[6] & Kwvmz6[3]));
assign Dlgyx6 = (Tlgyx6 & Bmgyx6);
assign Bmgyx6 = (~(Nsvmz6[6] & Kwvmz6[1]));
assign Tlgyx6 = (~(Sqvmz6[6] & Kwvmz6[2]));
assign Nkgyx6 = (Jmgyx6 & Rmgyx6);
assign Rmgyx6 = (~(Cnvmz6[6] & Kwvmz6[4]));
assign Jmgyx6 = (~(Kms7z6[6] & Kwvmz6[0]));
assign Dhgyx6 = (~(Nwfyx6 | Zufyx6));
assign Zufyx6 = (~(Zmgyx6 & Hngyx6));
assign Hngyx6 = (Pngyx6 & Xngyx6);
assign Xngyx6 = (~(Sqvmz6[5] & Kwvmz6[2]));
assign Pngyx6 = (Fogyx6 & Nogyx6);
assign Nogyx6 = (~(Nsvmz6[5] & Kwvmz6[1]));
assign Fogyx6 = (~(Xovmz6[5] & Kwvmz6[3]));
assign Zmgyx6 = (Vogyx6 & Dpgyx6);
assign Dpgyx6 = (~(Cnvmz6[5] & Kwvmz6[4]));
assign Vogyx6 = (~(Kms7z6[5] & Kwvmz6[0]));
assign Nwfyx6 = (~(Lpgyx6 & Tpgyx6));
assign Tpgyx6 = (Bqgyx6 & Jqgyx6);
assign Jqgyx6 = (~(Sqvmz6[4] & Kwvmz6[2]));
assign Bqgyx6 = (Rqgyx6 & Zqgyx6);
assign Zqgyx6 = (~(Nsvmz6[4] & Kwvmz6[1]));
assign Rqgyx6 = (~(Xovmz6[4] & Kwvmz6[3]));
assign Lpgyx6 = (Hrgyx6 & Prgyx6);
assign Prgyx6 = (~(Cnvmz6[4] & Kwvmz6[4]));
assign Hrgyx6 = (~(Kms7z6[4] & Kwvmz6[0]));
assign Tdgyx6 = (~(Lpfyx6 | Pzfyx6));
assign Pzfyx6 = (~(Xrgyx6 & Fsgyx6));
assign Fsgyx6 = (Nsgyx6 & Vsgyx6);
assign Vsgyx6 = (~(Sqvmz6[2] & Kwvmz6[2]));
assign Nsgyx6 = (Dtgyx6 & Ltgyx6);
assign Ltgyx6 = (~(Nsvmz6[2] & Kwvmz6[1]));
assign Dtgyx6 = (~(Xovmz6[2] & Kwvmz6[3]));
assign Xrgyx6 = (Ttgyx6 & Bugyx6);
assign Bugyx6 = (~(Cnvmz6[2] & Kwvmz6[4]));
assign Ttgyx6 = (~(Kms7z6[2] & Kwvmz6[0]));
assign Lpfyx6 = (~(Jugyx6 & Rugyx6));
assign Rugyx6 = (Zugyx6 & Hvgyx6);
assign Hvgyx6 = (~(Kwvmz6[2] & Sqvmz6[0]));
assign Zugyx6 = (Pvgyx6 & Xvgyx6);
assign Xvgyx6 = (~(Nsvmz6[0] & Kwvmz6[1]));
assign Pvgyx6 = (~(Kwvmz6[3] & Xovmz6[0]));
assign Jugyx6 = (Fwgyx6 & Nwgyx6);
assign Nwgyx6 = (~(Kwvmz6[4] & Cnvmz6[0]));
assign Fwgyx6 = (~(Kwvmz6[0] & Kms7z6[0]));
assign P7gyx6 = (Vwgyx6 & Dxgyx6);
assign Dxgyx6 = (~(Lxgyx6 & Txgyx6));
assign Txgyx6 = (~(Fbxmz6[3] & C55ov6));
assign Vwgyx6 = (~(Lxgyx6 & Bygyx6));
assign Bygyx6 = (B6byx6 | O9xmz6[1]);
assign V4gyx6 = (Hbgyx6 & Pj3yx6);
assign Pj3yx6 = (~(Jygyx6 & Pf5ov6));
assign Jygyx6 = (Rygyx6 & Zygyx6);
assign Hbgyx6 = (~(Hzgyx6 & Pzgyx6));
assign Pzgyx6 = (Xzgyx6 & Rygyx6);
assign Rygyx6 = (~(Zqbyx6 & La6ft6));
assign Xzgyx6 = (Eifnv6 & Jch7v6);
assign Hzgyx6 = (F0hyx6 & Pf5ov6);
assign F0hyx6 = (N0hyx6 & V0hyx6);
assign V0hyx6 = (~(D1hyx6 & B6byx6));
assign D1hyx6 = (~(P647v6 & Ak77z6));
assign B2gyx6 = (~(L1hyx6 & T1hyx6));
assign T1hyx6 = (B2hyx6 & J2hyx6);
assign J2hyx6 = (~(Sqvmz6[1] & Kwvmz6[2]));
assign B2hyx6 = (R2hyx6 & Z2hyx6);
assign Z2hyx6 = (~(Nsvmz6[1] & Kwvmz6[1]));
assign R2hyx6 = (~(Xovmz6[1] & Kwvmz6[3]));
assign L1hyx6 = (H3hyx6 & P3hyx6);
assign P3hyx6 = (~(Cnvmz6[1] & Kwvmz6[4]));
assign H3hyx6 = (~(Kms7z6[1] & Kwvmz6[0]));
assign Dmp7v6 = (Ab5ov6 ? X3hyx6 : Kh1nz6[2]);
assign Wlp7v6 = (Ue5ov6 ? X3hyx6 : Mm1nz6[2]);
assign Plp7v6 = (Ne5ov6 ? X3hyx6 : Nn1nz6[2]);
assign Ilp7v6 = (Ge5ov6 ? X3hyx6 : Oo1nz6[2]);
assign X3hyx6 = (~(F4hyx6 & N4hyx6));
assign N4hyx6 = (I347v6 ? D5hyx6 : V4hyx6);
assign D5hyx6 = (L5hyx6 & T5hyx6);
assign T5hyx6 = (B6hyx6 & J6hyx6);
assign J6hyx6 = (~(Mh5ov6 & Vcxmz6[23]));
assign B6hyx6 = (~(Vcxmz6[2] & Gjfnv6));
assign L5hyx6 = (R6hyx6 & Z6hyx6);
assign Z6hyx6 = (~(Hi5ov6 & Vcxmz6[16]));
assign R6hyx6 = (~(Oi5ov6 & Vcxmz6[9]));
assign V4hyx6 = (H7hyx6 & P7hyx6);
assign P7hyx6 = (~(Oi5ov6 & Vcxmz6[35]));
assign H7hyx6 = (X7hyx6 & F8hyx6);
assign F8hyx6 = (~(Gjfnv6 & Vcxmz6[28]));
assign X7hyx6 = (~(Hi5ov6 & Vcxmz6[42]));
assign F4hyx6 = (N8hyx6 & Ragyx6);
assign N8hyx6 = (~(V7xmz6[2] & Pf5ov6));
assign Blp7v6 = (Ab5ov6 ? V8hyx6 : Kh1nz6[3]);
assign Ukp7v6 = (Ue5ov6 ? V8hyx6 : Mm1nz6[3]);
assign Nkp7v6 = (Ne5ov6 ? V8hyx6 : Nn1nz6[3]);
assign Gkp7v6 = (Ge5ov6 ? V8hyx6 : Oo1nz6[3]);
assign V8hyx6 = (~(D9hyx6 & L9hyx6));
assign L9hyx6 = (~(V7xmz6[3] & Pf5ov6));
assign D9hyx6 = (I347v6 ? Bahyx6 : T9hyx6);
assign Bahyx6 = (Jahyx6 & Rahyx6);
assign Rahyx6 = (Zahyx6 & Hbhyx6);
assign Hbhyx6 = (~(Mh5ov6 & Vcxmz6[24]));
assign Zahyx6 = (~(Vcxmz6[3] & Gjfnv6));
assign Jahyx6 = (Pbhyx6 & Xbhyx6);
assign Xbhyx6 = (~(Hi5ov6 & Vcxmz6[17]));
assign Pbhyx6 = (~(Oi5ov6 & Vcxmz6[10]));
assign T9hyx6 = (Fchyx6 & Nchyx6);
assign Nchyx6 = (~(Oi5ov6 & Vcxmz6[36]));
assign Fchyx6 = (Vchyx6 & Ddhyx6);
assign Ddhyx6 = (~(Gjfnv6 & Vcxmz6[29]));
assign Vchyx6 = (~(Hi5ov6 & Vcxmz6[43]));
assign Zjp7v6 = (Ab5ov6 ? Ldhyx6 : Kh1nz6[4]);
assign Sjp7v6 = (Ue5ov6 ? Ldhyx6 : Mm1nz6[4]);
assign Ljp7v6 = (Ne5ov6 ? Ldhyx6 : Nn1nz6[4]);
assign Ejp7v6 = (Ge5ov6 ? Ldhyx6 : Oo1nz6[4]);
assign Ldhyx6 = (~(Tdhyx6 & Behyx6));
assign Behyx6 = (Jehyx6 & Ragyx6);
assign Tdhyx6 = (Rehyx6 & Zehyx6);
assign Zehyx6 = (~(V7xmz6[4] & Pf5ov6));
assign Rehyx6 = (I347v6 ? Pfhyx6 : Hfhyx6);
assign Pfhyx6 = (Xfhyx6 & Fghyx6);
assign Fghyx6 = (Nghyx6 & Vghyx6);
assign Vghyx6 = (~(Mh5ov6 & Vcxmz6[25]));
assign Nghyx6 = (~(Vcxmz6[4] & Gjfnv6));
assign Xfhyx6 = (Dhhyx6 & Lhhyx6);
assign Lhhyx6 = (~(Hi5ov6 & Vcxmz6[18]));
assign Dhhyx6 = (~(Oi5ov6 & Vcxmz6[11]));
assign Hfhyx6 = (Thhyx6 & Bihyx6);
assign Bihyx6 = (~(Oi5ov6 & Vcxmz6[37]));
assign Thhyx6 = (Jihyx6 & Rihyx6);
assign Rihyx6 = (~(Gjfnv6 & Vcxmz6[30]));
assign Jihyx6 = (~(Hi5ov6 & Vcxmz6[44]));
assign Xip7v6 = (Ab5ov6 ? Zihyx6 : Kh1nz6[5]);
assign Qip7v6 = (Ue5ov6 ? Zihyx6 : Mm1nz6[5]);
assign Jip7v6 = (Ne5ov6 ? Zihyx6 : Nn1nz6[5]);
assign Cip7v6 = (Ge5ov6 ? Zihyx6 : Oo1nz6[5]);
assign Zihyx6 = (~(Hjhyx6 & Pjhyx6));
assign Pjhyx6 = (I347v6 ? Fkhyx6 : Xjhyx6);
assign Fkhyx6 = (Nkhyx6 & Vkhyx6);
assign Vkhyx6 = (~(Oi5ov6 & Vcxmz6[12]));
assign Nkhyx6 = (Dlhyx6 & Llhyx6);
assign Llhyx6 = (~(Vcxmz6[5] & Gjfnv6));
assign Dlhyx6 = (~(Hi5ov6 & Vcxmz6[19]));
assign Xjhyx6 = (Tlhyx6 & Bmhyx6);
assign Bmhyx6 = (Jmhyx6 & Ragyx6);
assign Jmhyx6 = (~(Gjfnv6 & Vcxmz6[31]));
assign Tlhyx6 = (Rmhyx6 & Zmhyx6);
assign Zmhyx6 = (~(Hi5ov6 & Vcxmz6[45]));
assign Rmhyx6 = (~(Oi5ov6 & Vcxmz6[38]));
assign Hjhyx6 = (Hnhyx6 & Jehyx6);
assign Hnhyx6 = (~(V7xmz6[5] & Pf5ov6));
assign Vhp7v6 = (Ab5ov6 ? Pnhyx6 : Kh1nz6[6]);
assign Ohp7v6 = (Ue5ov6 ? Pnhyx6 : Mm1nz6[6]);
assign Hhp7v6 = (Ne5ov6 ? Pnhyx6 : Nn1nz6[6]);
assign Ahp7v6 = (Ge5ov6 ? Pnhyx6 : Oo1nz6[6]);
assign Pnhyx6 = (~(Xnhyx6 & Fohyx6));
assign Fohyx6 = (I347v6 ? Vohyx6 : Nohyx6);
assign Vohyx6 = (Dphyx6 & Lphyx6);
assign Lphyx6 = (Tphyx6 & Bqhyx6);
assign Bqhyx6 = (~(V147v6 & Mh5ov6));
assign Mh5ov6 = (!R6byx6);
assign R6byx6 = (~(Jqhyx6 & Rqhyx6));
assign Jqhyx6 = (Fbxmz6[2] & Fbxmz6[3]);
assign Tphyx6 = (~(Vcxmz6[6] & Gjfnv6));
assign Dphyx6 = (Zqhyx6 & Hrhyx6);
assign Hrhyx6 = (~(Hi5ov6 & Vcxmz6[20]));
assign Zqhyx6 = (~(Oi5ov6 & Vcxmz6[13]));
assign Nohyx6 = (Prhyx6 & Xrhyx6);
assign Xrhyx6 = (~(Oi5ov6 & Vcxmz6[39]));
assign Prhyx6 = (Fshyx6 & Nshyx6);
assign Nshyx6 = (~(Gjfnv6 & Vcxmz6[32]));
assign Fshyx6 = (~(Hi5ov6 & Vcxmz6[46]));
assign Xnhyx6 = (Vshyx6 & Jehyx6);
assign Jehyx6 = (~(Dthyx6 & Z6gyx6));
assign Vshyx6 = (~(V7xmz6[6] & Pf5ov6));
assign Tgp7v6 = (Ab5ov6 ? Lthyx6 : Kh1nz6[7]);
assign Ab5ov6 = (Apiiw6 & Tthyx6);
assign Tthyx6 = (~(Cc5ov6 & Buhyx6));
assign Buhyx6 = (~(Juhyx6 & Ruhyx6));
assign Cc5ov6 = (!Hae7v6);
assign Mgp7v6 = (Ue5ov6 ? Lthyx6 : Mm1nz6[7]);
assign Ue5ov6 = (Zuhyx6 & Nl5ov6);
assign Zuhyx6 = (Apiiw6 & Hvhyx6);
assign Fgp7v6 = (Ne5ov6 ? Lthyx6 : Nn1nz6[7]);
assign Ne5ov6 = (Pvhyx6 & Ul5ov6);
assign Pvhyx6 = (Apiiw6 & Xvhyx6);
assign Yfp7v6 = (Ge5ov6 ? Lthyx6 : Oo1nz6[7]);
assign Ge5ov6 = (Fwhyx6 & Apiiw6);
assign Apiiw6 = (Dniiw6 & Nwhyx6);
assign Nwhyx6 = (~(Vwhyx6 & Gl5ov6));
assign Vwhyx6 = (Dxhyx6 | Lxhyx6);
assign Dxhyx6 = (~(Txhyx6 & Byhyx6));
assign Dniiw6 = (~(Jyhyx6 | GATEHCLK));
assign Jyhyx6 = (~(HTMDHBURST[0] | Ue77z6));
assign Fwhyx6 = (Hvhyx6 & Xvhyx6);
assign Xvhyx6 = (!Nl5ov6);
assign Nl5ov6 = (Hae7v6 ? Pp1nz6[1] : Ruhyx6);
assign Hvhyx6 = (!Ul5ov6);
assign Ul5ov6 = (Hae7v6 ? Pp1nz6[0] : Juhyx6);
assign Lthyx6 = (~(Ryhyx6 & Zyhyx6));
assign Zyhyx6 = (Hzhyx6 & Pzhyx6);
assign Pzhyx6 = (~(H7gyx6 & Xzhyx6));
assign Xzhyx6 = (F0iyx6 | Gjfnv6);
assign Gjfnv6 = (B85ov6 & C55ov6);
assign B85ov6 = (Z6gyx6 & Fbxmz6[3]);
assign Z6gyx6 = (~(Ncgyx6 | Fbxmz6[1]));
assign F0iyx6 = (B6byx6 & N0iyx6);
assign N0iyx6 = (Hi5ov6 | Oi5ov6);
assign H7gyx6 = (!U75ov6);
assign U75ov6 = (~(B6byx6 | O9xmz6[0]));
assign B6byx6 = (!I347v6);
assign Hzhyx6 = (~(F4gyx6 | Dhbyx6));
assign Dhbyx6 = (!Ragyx6);
assign Ragyx6 = (~(V0iyx6 & D1iyx6));
assign D1iyx6 = (M35ov6 & C55ov6);
assign V0iyx6 = (Fbxmz6[3] & Ncgyx6);
assign F4gyx6 = (L1iyx6 & T1iyx6);
assign T1iyx6 = (Fbxmz6[0] & Vcgyx6);
assign L1iyx6 = (Fbxmz6[2] & Fbxmz6[1]);
assign Ryhyx6 = (B2iyx6 & J2iyx6);
assign J2iyx6 = (~(V7xmz6[7] & Pf5ov6));
assign B2iyx6 = (R2iyx6 & Z2iyx6);
assign Z2iyx6 = (~(O9xmz6[2] & Hi5ov6));
assign Hi5ov6 = (~(Z65ov6 | Vcgyx6));
assign Z65ov6 = (~(H3iyx6 & Fbxmz6[1]));
assign H3iyx6 = (Fbxmz6[0] & C55ov6);
assign R2iyx6 = (~(Oi5ov6 & O9xmz6[1]));
assign Oi5ov6 = (P3iyx6 & Lxgyx6);
assign Lxgyx6 = (Fbxmz6[1] & Ncgyx6);
assign P3iyx6 = (Fbxmz6[3] & C55ov6);
assign Rfp7v6 = (Dt2yx6 ? N52nz6[6] : X3iyx6);
assign X3iyx6 = (~(F4iyx6 & N4iyx6));
assign N4iyx6 = (~(V4iyx6 & D5iyx6));
assign D5iyx6 = (~(L5iyx6 | T5iyx6));
assign V4iyx6 = (F2f7v6 & B6iyx6);
assign B6iyx6 = (~(J6iyx6 & R6iyx6));
assign R6iyx6 = (~(Z6iyx6 & H7iyx6));
assign Z6iyx6 = (P7iyx6 & X7iyx6);
assign P7iyx6 = (F8iyx6 | R0f7v6);
assign J6iyx6 = (Xv2yx6 | Ik77z6);
assign Xv2yx6 = (!Od77z6);
assign F4iyx6 = (~(J72nz6[0] & Lx2yx6));
assign Kfp7v6 = (~(N8iyx6 & V8iyx6));
assign V8iyx6 = (D9iyx6 & Zu2yx6);
assign Zu2yx6 = (!L9iyx6);
assign D9iyx6 = (~(T9iyx6 & Baiyx6));
assign T9iyx6 = (J72nz6[0] & Ns2yx6);
assign N8iyx6 = (Jaiyx6 & Raiyx6);
assign Raiyx6 = (~(Wye7v6 & Zaiyx6));
assign Jaiyx6 = (~(Z12nz6[0] & Pv2yx6));
assign Dfp7v6 = (~(Hbiyx6 & Pbiyx6));
assign Pbiyx6 = (Xbiyx6 & Fciyx6);
assign Fciyx6 = (~(Nciyx6 & Mqb7z6[0]));
assign Xbiyx6 = (Vciyx6 & Ddiyx6);
assign Vciyx6 = (~(Ldiyx6 & Gh77z6));
assign Hbiyx6 = (Tdiyx6 & Beiyx6);
assign Beiyx6 = (~(Z12nz6[1] & Pv2yx6));
assign Tdiyx6 = (Jeiyx6 & Reiyx6);
assign Reiyx6 = (~(J72nz6[1] & Baiyx6));
assign Jeiyx6 = (~(N52nz6[0] & Zaiyx6));
assign Wep7v6 = (~(Zeiyx6 & Hfiyx6));
assign Hfiyx6 = (Pfiyx6 & Xfiyx6);
assign Xfiyx6 = (~(J72nz6[2] & Baiyx6));
assign Pfiyx6 = (Fgiyx6 & Ngiyx6);
assign Ngiyx6 = (~(Ldiyx6 & Wd77z6));
assign Fgiyx6 = (~(Nciyx6 & Mqb7z6[1]));
assign Zeiyx6 = (Vgiyx6 & Dhiyx6);
assign Dhiyx6 = (~(N52nz6[1] & Zaiyx6));
assign Vgiyx6 = (~(Z12nz6[2] & Pv2yx6));
assign Pep7v6 = (~(Lhiyx6 & Thiyx6));
assign Thiyx6 = (Biiyx6 & Jiiyx6);
assign Jiiyx6 = (~(Nciyx6 & Mqb7z6[2]));
assign Biiyx6 = (Riiyx6 & Ddiyx6);
assign Riiyx6 = (~(Ldiyx6 & Ee77z6));
assign Lhiyx6 = (Ziiyx6 & Hjiyx6);
assign Hjiyx6 = (~(Z12nz6[3] & Pv2yx6));
assign Ziiyx6 = (Pjiyx6 & Xjiyx6);
assign Xjiyx6 = (~(J72nz6[3] & Baiyx6));
assign Pjiyx6 = (~(N52nz6[2] & Zaiyx6));
assign Iep7v6 = (~(Fkiyx6 & Nkiyx6));
assign Nkiyx6 = (Vkiyx6 & Dliyx6);
assign Dliyx6 = (~(Nciyx6 & Mqb7z6[3]));
assign Vkiyx6 = (Lliyx6 & Ddiyx6);
assign Lliyx6 = (~(Ldiyx6 & Cf77z6));
assign Fkiyx6 = (Tliyx6 & Bmiyx6);
assign Bmiyx6 = (~(Z12nz6[4] & Pv2yx6));
assign Tliyx6 = (Jmiyx6 & Rmiyx6);
assign Rmiyx6 = (~(J72nz6[4] & Baiyx6));
assign Jmiyx6 = (~(N52nz6[3] & Zaiyx6));
assign Bep7v6 = (~(Zmiyx6 & Hniyx6));
assign Hniyx6 = (Pniyx6 & Xniyx6);
assign Xniyx6 = (~(Nciyx6 & Mqb7z6[4]));
assign Pniyx6 = (Foiyx6 & Ddiyx6);
assign Foiyx6 = (~(Ldiyx6 & Kf77z6));
assign Zmiyx6 = (Noiyx6 & Voiyx6);
assign Voiyx6 = (~(Z12nz6[5] & Pv2yx6));
assign Noiyx6 = (Dpiyx6 & Lpiyx6);
assign Lpiyx6 = (~(J72nz6[5] & Baiyx6));
assign Dpiyx6 = (~(N52nz6[4] & Zaiyx6));
assign Udp7v6 = (~(Tpiyx6 & Bqiyx6));
assign Bqiyx6 = (Jqiyx6 & Rqiyx6);
assign Rqiyx6 = (~(Nciyx6 & Mqb7z6[5]));
assign Jqiyx6 = (Zqiyx6 & Ddiyx6);
assign Zqiyx6 = (~(Ldiyx6 & Sf77z6));
assign Tpiyx6 = (Hriyx6 & Priyx6);
assign Priyx6 = (~(Z12nz6[6] & Pv2yx6));
assign Hriyx6 = (Xriyx6 & Fsiyx6);
assign Fsiyx6 = (~(J72nz6[6] & Baiyx6));
assign Xriyx6 = (~(N52nz6[5] & Zaiyx6));
assign Ndp7v6 = (~(Nsiyx6 & Vsiyx6));
assign Vsiyx6 = (Dtiyx6 & Ltiyx6);
assign Ltiyx6 = (~(Nciyx6 & Mqb7z6[6]));
assign Nciyx6 = (Ttiyx6 & L9iyx6);
assign Ttiyx6 = (~(Buiyx6 | Juiyx6));
assign Dtiyx6 = (Ruiyx6 & Ddiyx6);
assign Ddiyx6 = (~(Zuiyx6 & L9iyx6));
assign Zuiyx6 = (Juiyx6 & Hviyx6);
assign Hviyx6 = (!Buiyx6);
assign Ruiyx6 = (~(Ldiyx6 & Ag77z6));
assign Ldiyx6 = (Pviyx6 & L9iyx6);
assign L9iyx6 = (Xviyx6 & Fwiyx6);
assign Xviyx6 = (!Lx2yx6);
assign Pviyx6 = (Juiyx6 & Buiyx6);
assign Buiyx6 = (Vwiyx6 ? Nwiyx6 : Hp5ov6);
assign Juiyx6 = (Vwiyx6 ? Qa2nz6[0] : Dxiyx6);
assign Nsiyx6 = (Lxiyx6 & Txiyx6);
assign Txiyx6 = (~(Z12nz6[7] & Pv2yx6));
assign Lxiyx6 = (Byiyx6 & Jyiyx6);
assign Jyiyx6 = (~(J72nz6[7] & Baiyx6));
assign Baiyx6 = (Ryiyx6 & Fwiyx6);
assign Byiyx6 = (~(Zaiyx6 & N52nz6[6]));
assign Zaiyx6 = (~(Pv2yx6 | J23yx6));
assign Pv2yx6 = (!Fwiyx6);
assign Fwiyx6 = (Zyiyx6 & Mo5ov6);
assign Gdp7v6 = (Hziyx6 | Pziyx6);
assign Pziyx6 = (~(Xziyx6 | F0jyx6));
assign F0jyx6 = (D1jyx6 ? V0jyx6 : N0jyx6);
assign N0jyx6 = (Nl1nz6[1] | Ctf7v6);
assign Xziyx6 = (Ld2yx6 | Dl2yx6);
assign Dl2yx6 = (~(L1jyx6 | T1jyx6));
assign L1jyx6 = (B63yx6 ? D53yx6 : J7f7v6);
assign Ld2yx6 = (~(B2jyx6 & Nl1nz6[0]));
assign Hziyx6 = (Nl1nz6[1] ? R2jyx6 : J2jyx6);
assign R2jyx6 = (Mwf7v6 ? Pb2yx6 : Z2jyx6);
assign Z2jyx6 = (D1jyx6 | Qk77z6);
assign J2jyx6 = (H3jyx6 & Fs2yx6);
assign Fs2yx6 = (Qk77z6 & Mwf7v6);
assign H3jyx6 = (Ctf7v6 & Nl1nz6[0]);
assign Zcp7v6 = (P3jyx6 & X3jyx6);
assign Scp7v6 = (~(F4jyx6 & N4jyx6));
assign N4jyx6 = (~(P3jyx6 & V4jyx6));
assign V4jyx6 = (~(D5jyx6 & L5jyx6));
assign L5jyx6 = (~(T5jyx6 & B6jyx6));
assign D5jyx6 = (~(J6jyx6 & R6jyx6));
assign F4jyx6 = (~(Z6jyx6 & H7jyx6));
assign Lcp7v6 = (~(P7jyx6 | X7jyx6));
assign Ecp7v6 = (F8jyx6 & D1jyx6);
assign D1jyx6 = (~(N8jyx6 & V8jyx6));
assign V8jyx6 = (D9jyx6 & L9jyx6);
assign L9jyx6 = (~(P3jyx6 & T9jyx6));
assign T9jyx6 = (~(Bajyx6 & Jajyx6));
assign Jajyx6 = (~(T5jyx6 & Rajyx6));
assign Bajyx6 = (~(J6jyx6 & Zajyx6));
assign D9jyx6 = (~(H7jyx6 & Hbjyx6));
assign Hbjyx6 = (Twhiw6 | Iy1nz6[0]);
assign H7jyx6 = (X3jyx6 | Pbjyx6);
assign Pbjyx6 = (Xbjyx6 & Fcjyx6);
assign Fcjyx6 = (Kf2nz6[2] ? R6jyx6 : B6jyx6);
assign R6jyx6 = (~(Ncjyx6 & Vcjyx6));
assign Vcjyx6 = (Mo5ov6 | Ddjyx6);
assign Ncjyx6 = (Ldjyx6 & Tdjyx6);
assign Ldjyx6 = (~(Z12nz6[5] & Bejyx6));
assign B6jyx6 = (~(Jejyx6 & Rejyx6));
assign Rejyx6 = (~(B63yx6 & Zejyx6));
assign Jejyx6 = (Hfjyx6 & Tdjyx6);
assign Hfjyx6 = (~(Z12nz6[1] & Bejyx6));
assign Xbjyx6 = (Kf2nz6[0] & Pfjyx6);
assign X3jyx6 = (~(Xfjyx6 & Fgjyx6));
assign Fgjyx6 = (~(T5jyx6 & Ngjyx6));
assign Ngjyx6 = (~(Vgjyx6 & Dhjyx6));
assign Dhjyx6 = (Mo5ov6 | Lhjyx6);
assign Vgjyx6 = (Thjyx6 & Tdjyx6);
assign Thjyx6 = (~(Z12nz6[3] & Bejyx6));
assign Xfjyx6 = (~(Bijyx6 & J6jyx6));
assign Bijyx6 = (Bejyx6 ? Z12nz6[7] : Jijyx6);
assign Jijyx6 = (!Rijyx6);
assign Rijyx6 = (Mo5ov6 ? Ca1nv6 : Zijyx6);
assign N8jyx6 = (Hjjyx6 & Pjjyx6);
assign Pjjyx6 = (Xjjyx6 | X7jyx6);
assign X7jyx6 = (Fkjyx6 & Nkjyx6);
assign Nkjyx6 = (~(J6jyx6 & Vkjyx6));
assign Fkjyx6 = (~(T5jyx6 & Dljyx6));
assign Hjjyx6 = (Kf2nz6[1] ? Tljyx6 : Lljyx6);
assign Tljyx6 = (~(Bmjyx6 & Dp2yx6));
assign Bmjyx6 = (Kf2nz6[2] ? Vkjyx6 : Dljyx6);
assign Vkjyx6 = (~(Jmjyx6 & Rmjyx6));
assign Rmjyx6 = (~(B63yx6 & Zmjyx6));
assign Jmjyx6 = (Hnjyx6 & Tdjyx6);
assign Hnjyx6 = (~(Z12nz6[6] & Bejyx6));
assign Dljyx6 = (~(Pnjyx6 & Xnjyx6));
assign Xnjyx6 = (Mo5ov6 | Fojyx6);
assign Pnjyx6 = (Nojyx6 & Tdjyx6);
assign Nojyx6 = (~(Z12nz6[2] & Bejyx6));
assign Lljyx6 = (~(Vojyx6 & Dpjyx6));
assign Dpjyx6 = (~(Kf2nz6[0] & Xjjyx6));
assign Vojyx6 = (Kf2nz6[2] ? Zajyx6 : Rajyx6);
assign Zajyx6 = (~(Lpjyx6 & Tpjyx6));
assign Tpjyx6 = (Mo5ov6 | Bqjyx6);
assign Lpjyx6 = (Jqjyx6 & Tdjyx6);
assign Jqjyx6 = (~(Z12nz6[4] & Bejyx6));
assign Rajyx6 = (~(Rqjyx6 & Zqjyx6));
assign Zqjyx6 = (Mo5ov6 | Hrjyx6);
assign Rqjyx6 = (Prjyx6 & Tdjyx6);
assign Tdjyx6 = (!T1jyx6);
assign T1jyx6 = (Xrjyx6 & Mo5ov6);
assign Prjyx6 = (~(Z12nz6[0] & Bejyx6));
assign F8jyx6 = (~(Fsjyx6 & Nsjyx6));
assign Nsjyx6 = (Vsjyx6 & Hih7v6);
assign Vsjyx6 = (Aih7v6 & Twhiw6);
assign Fsjyx6 = (Vih7v6 & Oih7v6);
assign Xbp7v6 = (~(Dtjyx6 & Ltjyx6));
assign Ltjyx6 = (~(L8wnv6 & Itb7z6[29]));
assign Dtjyx6 = (Ttjyx6 & Bujyx6);
assign Bujyx6 = (~(G9wnv6 & Jujyx6));
assign Jujyx6 = (~(Rujyx6 & Zujyx6));
assign Zujyx6 = (Hvjyx6 & Pvjyx6);
assign Pvjyx6 = (Wawnv6 | Xvjyx6);
assign Wawnv6 = (!Dtm7z6[2]);
assign Hvjyx6 = (~(Dtm7z6[3] & Fwjyx6));
assign Rujyx6 = (Nwjyx6 & Vwjyx6);
assign Vwjyx6 = (~(Dtm7z6[0] & HRDATAD[29]));
assign Nwjyx6 = (~(Dtm7z6[1] & HRDATAS[29]));
assign Ttjyx6 = (~(Fcwnv6 & Ymyhw6));
assign Ymyhw6 = (Dz1nv6 ? Ulxmz6[29] : Aixmz6[29]);
assign Qbp7v6 = (~(Dxjyx6 & Lxjyx6));
assign Lxjyx6 = (~(Txjyx6 & Zec7z6[0]));
assign Dxjyx6 = (Byjyx6 & Jyjyx6);
assign Jyjyx6 = (~(H5xnv6 & Kaxnv6));
assign Kaxnv6 = (~(Ryjyx6 & Zyjyx6));
assign Zyjyx6 = (~(G7piw6 & HRDATAS[0]));
assign Ryjyx6 = (Hzjyx6 & Pzjyx6);
assign Pzjyx6 = (~(K9piw6 & Orwnv6));
assign Hzjyx6 = (~(HRDATAI[0] & Xzjyx6));
assign Byjyx6 = (~(Byc7z6[0] & O5xnv6));
assign Jbp7v6 = (~(F0kyx6 & N0kyx6));
assign N0kyx6 = (~(Txjyx6 & Zec7z6[1]));
assign F0kyx6 = (V0kyx6 & D1kyx6);
assign D1kyx6 = (~(H5xnv6 & B1ynv6));
assign B1ynv6 = (~(L1kyx6 & T1kyx6));
assign T1kyx6 = (~(G7piw6 & HRDATAS[1]));
assign L1kyx6 = (B2kyx6 & J2kyx6);
assign J2kyx6 = (~(K9piw6 & Kud7x6));
assign B2kyx6 = (~(HRDATAI[1] & Xzjyx6));
assign V0kyx6 = (~(Byc7z6[1] & O5xnv6));
assign Cbp7v6 = (~(R2kyx6 & Z2kyx6));
assign Z2kyx6 = (~(Txjyx6 & Zec7z6[2]));
assign R2kyx6 = (H3kyx6 & P3kyx6);
assign P3kyx6 = (~(H5xnv6 & Mwxnv6));
assign Mwxnv6 = (~(X3kyx6 & F4kyx6));
assign F4kyx6 = (~(G7piw6 & HRDATAS[2]));
assign X3kyx6 = (N4kyx6 & V4kyx6);
assign V4kyx6 = (~(K9piw6 & Eyd7x6));
assign N4kyx6 = (~(HRDATAI[2] & Xzjyx6));
assign H3kyx6 = (~(Byc7z6[2] & O5xnv6));
assign Vap7v6 = (~(D5kyx6 & L5kyx6));
assign L5kyx6 = (~(Txjyx6 & Zec7z6[3]));
assign D5kyx6 = (T5kyx6 & B6kyx6);
assign B6kyx6 = (~(H5xnv6 & Xrxnv6));
assign Xrxnv6 = (~(J6kyx6 & R6kyx6));
assign R6kyx6 = (~(G7piw6 & HRDATAS[3]));
assign J6kyx6 = (Z6kyx6 & H7kyx6);
assign H7kyx6 = (~(K9piw6 & R1e7x6));
assign Z6kyx6 = (~(HRDATAI[3] & Xzjyx6));
assign T5kyx6 = (~(Byc7z6[3] & O5xnv6));
assign Oap7v6 = (~(P7kyx6 & X7kyx6));
assign X7kyx6 = (~(Txjyx6 & Zec7z6[4]));
assign P7kyx6 = (F8kyx6 & N8kyx6);
assign N8kyx6 = (~(H5xnv6 & Inxnv6));
assign Inxnv6 = (~(V8kyx6 & D9kyx6));
assign D9kyx6 = (~(G7piw6 & HRDATAS[4]));
assign V8kyx6 = (L9kyx6 & T9kyx6);
assign T9kyx6 = (~(K9piw6 & E5e7x6));
assign L9kyx6 = (~(HRDATAI[4] & Xzjyx6));
assign F8kyx6 = (~(Byc7z6[4] & O5xnv6));
assign Hap7v6 = (~(Bakyx6 & Jakyx6));
assign Jakyx6 = (~(Txjyx6 & Zec7z6[5]));
assign Bakyx6 = (Rakyx6 & Zakyx6);
assign Zakyx6 = (~(H5xnv6 & Tixnv6));
assign Tixnv6 = (~(Hbkyx6 & Pbkyx6));
assign Pbkyx6 = (~(G7piw6 & HRDATAS[5]));
assign Hbkyx6 = (Xbkyx6 & Fckyx6);
assign Fckyx6 = (~(K9piw6 & R8e7x6));
assign Xbkyx6 = (~(HRDATAI[5] & Xzjyx6));
assign Rakyx6 = (~(Byc7z6[5] & O5xnv6));
assign Aap7v6 = (~(Nckyx6 & Vckyx6));
assign Vckyx6 = (~(Txjyx6 & Zec7z6[6]));
assign Nckyx6 = (Ddkyx6 & Ldkyx6);
assign Ldkyx6 = (~(H5xnv6 & Eexnv6));
assign Eexnv6 = (~(Tdkyx6 & Bekyx6));
assign Bekyx6 = (~(G7piw6 & HRDATAS[6]));
assign Tdkyx6 = (Jekyx6 & Rekyx6);
assign Rekyx6 = (~(K9piw6 & Ece7x6));
assign Jekyx6 = (~(HRDATAI[6] & Xzjyx6));
assign Ddkyx6 = (~(Byc7z6[6] & O5xnv6));
assign T9p7v6 = (~(Zekyx6 & Hfkyx6));
assign Hfkyx6 = (~(Txjyx6 & Zec7z6[7]));
assign Zekyx6 = (Pfkyx6 & Xfkyx6);
assign Xfkyx6 = (~(H5xnv6 & N1xnv6));
assign N1xnv6 = (~(Fgkyx6 & Ngkyx6));
assign Ngkyx6 = (~(G7piw6 & HRDATAS[7]));
assign Fgkyx6 = (Vgkyx6 & Dhkyx6);
assign Dhkyx6 = (~(K9piw6 & Rfe7x6));
assign Vgkyx6 = (~(HRDATAI[7] & Xzjyx6));
assign Pfkyx6 = (~(Byc7z6[7] & O5xnv6));
assign M9p7v6 = (~(Lhkyx6 & Thkyx6));
assign Thkyx6 = (~(Txjyx6 & Zec7z6[8]));
assign Lhkyx6 = (Bikyx6 & Jikyx6);
assign Jikyx6 = (~(H5xnv6 & S5znv6));
assign S5znv6 = (~(Rikyx6 & Zikyx6));
assign Zikyx6 = (~(G7piw6 & HRDATAS[8]));
assign Rikyx6 = (Hjkyx6 & Pjkyx6);
assign Pjkyx6 = (~(K9piw6 & Ebf7x6));
assign Hjkyx6 = (~(HRDATAI[8] & Xzjyx6));
assign Bikyx6 = (~(Byc7z6[8] & O5xnv6));
assign F9p7v6 = (~(Xjkyx6 & Fkkyx6));
assign Fkkyx6 = (~(Txjyx6 & Zec7z6[9]));
assign Xjkyx6 = (Nkkyx6 & Vkkyx6);
assign Vkkyx6 = (~(H5xnv6 & D1znv6));
assign D1znv6 = (~(Dlkyx6 & Llkyx6));
assign Llkyx6 = (Tlkyx6 & Bmkyx6);
assign Tlkyx6 = (~(K9piw6 & Rme7x6));
assign Dlkyx6 = (Jmkyx6 & Rmkyx6);
assign Rmkyx6 = (~(HRDATAI[9] & D9piw6));
assign Jmkyx6 = (~(G7piw6 & HRDATAS[9]));
assign Nkkyx6 = (~(Byc7z6[9] & O5xnv6));
assign Y8p7v6 = (~(Zmkyx6 & Hnkyx6));
assign Hnkyx6 = (~(Txjyx6 & Zec7z6[10]));
assign Zmkyx6 = (Pnkyx6 & Xnkyx6);
assign Xnkyx6 = (~(H5xnv6 & Owynv6));
assign Owynv6 = (~(Fokyx6 & Nokyx6));
assign Nokyx6 = (Vokyx6 & Bmkyx6);
assign Vokyx6 = (~(K9piw6 & Eqe7x6));
assign Fokyx6 = (Dpkyx6 & Lpkyx6);
assign Lpkyx6 = (~(HRDATAI[10] & D9piw6));
assign Dpkyx6 = (~(G7piw6 & HRDATAS[10]));
assign Pnkyx6 = (~(Byc7z6[10] & O5xnv6));
assign R8p7v6 = (~(Tpkyx6 & Bqkyx6));
assign Bqkyx6 = (~(Txjyx6 & Zec7z6[11]));
assign Tpkyx6 = (Jqkyx6 & Rqkyx6);
assign Rqkyx6 = (~(H5xnv6 & Zrynv6));
assign Zrynv6 = (~(Zqkyx6 & Hrkyx6));
assign Hrkyx6 = (Prkyx6 & Bmkyx6);
assign Prkyx6 = (~(K9piw6 & Rte7x6));
assign Zqkyx6 = (Xrkyx6 & Fskyx6);
assign Fskyx6 = (~(HRDATAI[11] & D9piw6));
assign Xrkyx6 = (~(G7piw6 & HRDATAS[11]));
assign Jqkyx6 = (~(Byc7z6[11] & O5xnv6));
assign K8p7v6 = (~(Nskyx6 & Vskyx6));
assign Vskyx6 = (~(Txjyx6 & Zec7z6[12]));
assign Nskyx6 = (Dtkyx6 & Ltkyx6);
assign Ltkyx6 = (~(H5xnv6 & Knynv6));
assign Knynv6 = (~(Ttkyx6 & Bukyx6));
assign Bukyx6 = (Jukyx6 & Bmkyx6);
assign Jukyx6 = (~(K9piw6 & Exe7x6));
assign Ttkyx6 = (Rukyx6 & Zukyx6);
assign Zukyx6 = (~(HRDATAI[12] & D9piw6));
assign Rukyx6 = (~(G7piw6 & HRDATAS[12]));
assign Dtkyx6 = (~(Byc7z6[12] & O5xnv6));
assign D8p7v6 = (~(Hvkyx6 & Pvkyx6));
assign Pvkyx6 = (~(Txjyx6 & Zec7z6[13]));
assign Hvkyx6 = (Xvkyx6 & Fwkyx6);
assign Fwkyx6 = (~(H5xnv6 & Viynv6));
assign Viynv6 = (~(Nwkyx6 & Vwkyx6));
assign Vwkyx6 = (Dxkyx6 & Bmkyx6);
assign Dxkyx6 = (~(K9piw6 & R0f7x6));
assign Nwkyx6 = (Lxkyx6 & Txkyx6);
assign Txkyx6 = (~(HRDATAI[13] & D9piw6));
assign Lxkyx6 = (~(G7piw6 & HRDATAS[13]));
assign Xvkyx6 = (~(Byc7z6[13] & O5xnv6));
assign W7p7v6 = (~(Bykyx6 & Jykyx6));
assign Jykyx6 = (~(Byc7z6[14] & O5xnv6));
assign Bykyx6 = (Rykyx6 & Rdtov6);
assign Rykyx6 = (~(H5xnv6 & Geynv6));
assign P7p7v6 = (~(Zykyx6 & Hzkyx6));
assign Hzkyx6 = (~(Txjyx6 & Zec7z6[15]));
assign Zykyx6 = (Pzkyx6 & Xzkyx6);
assign Xzkyx6 = (~(H5xnv6 & R9ynv6));
assign Pzkyx6 = (~(Byc7z6[15] & O5xnv6));
assign I7p7v6 = (~(F0lyx6 & N0lyx6));
assign N0lyx6 = (~(Txjyx6 & Zec7z6[16]));
assign F0lyx6 = (V0lyx6 & D1lyx6);
assign D1lyx6 = (~(H5xnv6 & N6znv6));
assign V0lyx6 = (~(Byc7z6[16] & O5xnv6));
assign B7p7v6 = (~(L1lyx6 & T1lyx6));
assign T1lyx6 = (~(Txjyx6 & Zec7z6[17]));
assign L1lyx6 = (B2lyx6 & J2lyx6);
assign J2lyx6 = (~(H5xnv6 & Y1znv6));
assign Y1znv6 = (~(R2lyx6 & Z2lyx6));
assign Z2lyx6 = (~(G7piw6 & HRDATAS[17]));
assign R2lyx6 = (H3lyx6 & P3lyx6);
assign P3lyx6 = (~(K9piw6 & Agf7x6));
assign H3lyx6 = (~(HRDATAI[17] & X3lyx6));
assign B2lyx6 = (~(Byc7z6[17] & O5xnv6));
assign U6p7v6 = (~(F4lyx6 & N4lyx6));
assign N4lyx6 = (~(Txjyx6 & Zec7z6[18]));
assign F4lyx6 = (V4lyx6 & D5lyx6);
assign D5lyx6 = (~(H5xnv6 & Jxynv6));
assign Jxynv6 = (~(L5lyx6 & T5lyx6));
assign T5lyx6 = (~(G7piw6 & HRDATAS[18]));
assign L5lyx6 = (B6lyx6 & J6lyx6);
assign J6lyx6 = (~(K9piw6 & Njf7x6));
assign B6lyx6 = (~(HRDATAI[18] & X3lyx6));
assign V4lyx6 = (~(Byc7z6[18] & O5xnv6));
assign N6p7v6 = (~(R6lyx6 & Z6lyx6));
assign Z6lyx6 = (~(Txjyx6 & Zec7z6[19]));
assign R6lyx6 = (H7lyx6 & P7lyx6);
assign P7lyx6 = (~(H5xnv6 & Usynv6));
assign Usynv6 = (~(X7lyx6 & F8lyx6));
assign F8lyx6 = (~(G7piw6 & HRDATAS[19]));
assign X7lyx6 = (N8lyx6 & V8lyx6);
assign V8lyx6 = (~(K9piw6 & Anf7x6));
assign N8lyx6 = (~(HRDATAI[19] & X3lyx6));
assign H7lyx6 = (~(Byc7z6[19] & O5xnv6));
assign G6p7v6 = (~(D9lyx6 & L9lyx6));
assign L9lyx6 = (~(Txjyx6 & Zec7z6[20]));
assign D9lyx6 = (T9lyx6 & Balyx6);
assign Balyx6 = (~(H5xnv6 & Foynv6));
assign Foynv6 = (~(Jalyx6 & Ralyx6));
assign Ralyx6 = (~(G7piw6 & HRDATAS[20]));
assign Jalyx6 = (Zalyx6 & Hblyx6);
assign Hblyx6 = (~(K9piw6 & Nqf7x6));
assign Zalyx6 = (~(HRDATAI[20] & X3lyx6));
assign T9lyx6 = (~(Byc7z6[20] & O5xnv6));
assign Z5p7v6 = (~(Pblyx6 & Xblyx6));
assign Xblyx6 = (~(Txjyx6 & Zec7z6[21]));
assign Pblyx6 = (Fclyx6 & Nclyx6);
assign Nclyx6 = (~(H5xnv6 & Qjynv6));
assign Qjynv6 = (~(Vclyx6 & Ddlyx6));
assign Ddlyx6 = (~(G7piw6 & HRDATAS[21]));
assign Vclyx6 = (Ldlyx6 & Tdlyx6);
assign Tdlyx6 = (~(K9piw6 & Auf7x6));
assign Ldlyx6 = (~(HRDATAI[21] & X3lyx6));
assign Fclyx6 = (~(Byc7z6[21] & O5xnv6));
assign S5p7v6 = (~(Belyx6 & Jelyx6));
assign Jelyx6 = (~(Txjyx6 & Zec7z6[22]));
assign Belyx6 = (Relyx6 & Zelyx6);
assign Zelyx6 = (~(H5xnv6 & Bfynv6));
assign Bfynv6 = (~(Hflyx6 & Pflyx6));
assign Pflyx6 = (~(G7piw6 & HRDATAS[22]));
assign Hflyx6 = (Xflyx6 & Fglyx6);
assign Fglyx6 = (~(K9piw6 & Nxf7x6));
assign Xflyx6 = (~(HRDATAI[22] & X3lyx6));
assign Relyx6 = (~(Byc7z6[22] & O5xnv6));
assign L5p7v6 = (~(Nglyx6 & Vglyx6));
assign Vglyx6 = (~(Txjyx6 & Zec7z6[23]));
assign Nglyx6 = (Dhlyx6 & Lhlyx6);
assign Lhlyx6 = (~(H5xnv6 & Maynv6));
assign Maynv6 = (~(Thlyx6 & Bilyx6));
assign Bilyx6 = (~(G7piw6 & HRDATAS[23]));
assign Thlyx6 = (Jilyx6 & Rilyx6);
assign Rilyx6 = (~(K9piw6 & A1g7x6));
assign Jilyx6 = (~(HRDATAI[23] & X3lyx6));
assign Dhlyx6 = (~(Byc7z6[23] & O5xnv6));
assign E5p7v6 = (~(Zilyx6 & Hjlyx6));
assign Hjlyx6 = (~(Txjyx6 & Zec7z6[24]));
assign Zilyx6 = (Pjlyx6 & Xjlyx6);
assign Xjlyx6 = (~(H5xnv6 & P9xnv6));
assign P9xnv6 = (~(Fklyx6 & Nklyx6));
assign Nklyx6 = (~(G7piw6 & HRDATAS[24]));
assign Fklyx6 = (Vklyx6 & Dllyx6);
assign Dllyx6 = (~(K9piw6 & Kdg7x6));
assign Vklyx6 = (~(HRDATAI[24] & X3lyx6));
assign Pjlyx6 = (~(Byc7z6[24] & O5xnv6));
assign X4p7v6 = (~(Lllyx6 & Tllyx6));
assign Tllyx6 = (~(Txjyx6 & Zec7z6[25]));
assign Lllyx6 = (Bmlyx6 & Jmlyx6);
assign Jmlyx6 = (~(H5xnv6 & W1ynv6));
assign W1ynv6 = (~(Rmlyx6 & Zmlyx6));
assign Zmlyx6 = (Hnlyx6 & Pnlyx6);
assign Hnlyx6 = (~(K9piw6 & X9g7x6));
assign Rmlyx6 = (Xnlyx6 & Folyx6);
assign Folyx6 = (~(HRDATAI[25] & D9piw6));
assign Xnlyx6 = (~(G7piw6 & HRDATAS[25]));
assign Bmlyx6 = (~(Byc7z6[25] & O5xnv6));
assign Q4p7v6 = (~(Nolyx6 & Volyx6));
assign Volyx6 = (~(Txjyx6 & Zec7z6[26]));
assign Nolyx6 = (Dplyx6 & Lplyx6);
assign Lplyx6 = (~(H5xnv6 & Hxxnv6));
assign Hxxnv6 = (~(Tplyx6 & Bqlyx6));
assign Bqlyx6 = (Jqlyx6 & Pnlyx6);
assign Jqlyx6 = (~(K9piw6 & Dx98x6));
assign Tplyx6 = (Rqlyx6 & Zqlyx6);
assign Zqlyx6 = (~(HRDATAI[26] & D9piw6));
assign Rqlyx6 = (~(G7piw6 & HRDATAS[26]));
assign Dplyx6 = (~(Byc7z6[26] & O5xnv6));
assign J4p7v6 = (~(Hrlyx6 & Prlyx6));
assign Prlyx6 = (~(Txjyx6 & Zec7z6[27]));
assign Hrlyx6 = (Xrlyx6 & Fslyx6);
assign Fslyx6 = (~(H5xnv6 & Ssxnv6));
assign Ssxnv6 = (~(Nslyx6 & Vslyx6));
assign Vslyx6 = (Dtlyx6 & Pnlyx6);
assign Dtlyx6 = (~(K9piw6 & Dpyxx6));
assign Nslyx6 = (Ltlyx6 & Ttlyx6);
assign Ttlyx6 = (~(HRDATAI[27] & D9piw6));
assign Ltlyx6 = (~(G7piw6 & HRDATAS[27]));
assign Xrlyx6 = (~(Byc7z6[27] & O5xnv6));
assign C4p7v6 = (~(Bulyx6 & Julyx6));
assign Julyx6 = (~(Txjyx6 & Zec7z6[28]));
assign Bulyx6 = (Rulyx6 & Zulyx6);
assign Zulyx6 = (~(H5xnv6 & Doxnv6));
assign Doxnv6 = (~(Hvlyx6 & Pvlyx6));
assign Pvlyx6 = (Xvlyx6 & Pnlyx6);
assign Xvlyx6 = (~(K9piw6 & Dtyxx6));
assign Hvlyx6 = (Fwlyx6 & Nwlyx6);
assign Nwlyx6 = (~(HRDATAI[28] & D9piw6));
assign Fwlyx6 = (~(G7piw6 & HRDATAS[28]));
assign Rulyx6 = (~(Byc7z6[28] & O5xnv6));
assign V3p7v6 = (~(Vwlyx6 & Dxlyx6));
assign Dxlyx6 = (~(Txjyx6 & Zec7z6[29]));
assign Vwlyx6 = (Lxlyx6 & Txlyx6);
assign Txlyx6 = (~(H5xnv6 & Ojxnv6));
assign Ojxnv6 = (~(Bylyx6 & Jylyx6));
assign Jylyx6 = (Rylyx6 & Pnlyx6);
assign Rylyx6 = (~(K9piw6 & Fwjyx6));
assign Bylyx6 = (Zylyx6 & Hzlyx6);
assign Hzlyx6 = (~(HRDATAI[29] & D9piw6));
assign Zylyx6 = (~(G7piw6 & HRDATAS[29]));
assign Lxlyx6 = (~(Byc7z6[29] & O5xnv6));
assign O3p7v6 = (~(Pzlyx6 & Xzlyx6));
assign Xzlyx6 = (~(Txjyx6 & Zec7z6[30]));
assign Pzlyx6 = (F0myx6 & N0myx6);
assign N0myx6 = (~(H5xnv6 & Zexnv6));
assign F0myx6 = (~(Byc7z6[30] & O5xnv6));
assign H3p7v6 = (~(V0myx6 & D1myx6));
assign D1myx6 = (~(Txjyx6 & Zec7z6[31]));
assign V0myx6 = (L1myx6 & T1myx6);
assign T1myx6 = (~(H5xnv6 & P2xnv6));
assign H5xnv6 = (~(O5xnv6 | Txjyx6));
assign Txjyx6 = (!Rdtov6);
assign L1myx6 = (~(Byc7z6[31] & O5xnv6));
assign O5xnv6 = (Opqov6 & Rdtov6);
assign Opqov6 = (!Hpqov6);
assign Hpqov6 = (P6d7z6[2] & Cg1ov6);
assign A3p7v6 = (~(B2myx6 & J2myx6));
assign J2myx6 = (~(R2myx6 & Z2myx6));
assign R2myx6 = (~(Jfonv6 | H3myx6));
assign B2myx6 = (~(P3myx6 & Eqn7z6[0]));
assign T2p7v6 = (~(X3myx6 & F4myx6));
assign F4myx6 = (~(N4myx6 & Z2myx6));
assign N4myx6 = (~(V4myx6 | H3myx6));
assign X3myx6 = (~(Eqn7z6[1] & P3myx6));
assign M2p7v6 = (~(D5myx6 & L5myx6));
assign L5myx6 = (~(Eqn7z6[2] & P3myx6));
assign D5myx6 = (T5myx6 & B6myx6);
assign B6myx6 = (~(Z2myx6 & Jn1ov6));
assign Z2myx6 = (~(P3myx6 | J6myx6));
assign J6myx6 = (!HWRITED);
assign P3myx6 = (R6myx6 & Goonv6);
assign T5myx6 = (~(H3myx6 & HWRITED));
assign HWRITED = (~(Z6myx6 & H7myx6));
assign H7myx6 = (~(Hm1ov6 & Lhmov6));
assign Z6myx6 = (P7myx6 & X7myx6);
assign X7myx6 = (~(I2yet6 & Jn1ov6));
assign P7myx6 = (~(L3bdt6 & Vm1ov6));
assign H3myx6 = (~(R6myx6 | HREADYD));
assign R6myx6 = (~(Eqn7z6[0] & Qtixx6));
assign Qtixx6 = (F8myx6 & I2yet6);
assign F8myx6 = (Qmonv6 & N8myx6);
assign N8myx6 = (~(V8myx6 & Y497z6));
assign V8myx6 = (~(U8oet6 | Qboet6));
assign F2p7v6 = (Wj1ov6 ? X0d7z6[31] : Dvc7z6[31]);
assign Y1p7v6 = (Wj1ov6 ? X0d7z6[30] : Dvc7z6[30]);
assign R1p7v6 = (~(D9myx6 & L9myx6));
assign L9myx6 = (~(Gonov6 & K9d7x6));
assign D9myx6 = (T9myx6 & Bamyx6);
assign Bamyx6 = (~(Jamyx6 & Ramyx6));
assign Ramyx6 = (Zamyx6 & Hbmyx6);
assign Hbmyx6 = (~(D2piw6 & Bpnov6));
assign D2piw6 = (!Qv0ov6);
assign Zamyx6 = (Pbmyx6 & Vs9ov6);
assign Pbmyx6 = (~(Xbmyx6 & Qu1ov6));
assign Qu1ov6 = (Zo1ov6 | Yrc8v6);
assign Yrc8v6 = (~(Ufphw6 | Dwb7z6[4]));
assign Ufphw6 = (~(Ce9iw6 & Fcmyx6));
assign Ce9iw6 = (Ncmyx6 & Vcmyx6);
assign Vcmyx6 = (Ddmyx6 & Ldmyx6);
assign Ddmyx6 = (Tdmyx6 & Bemyx6);
assign Bemyx6 = (!Qij7z6[3]);
assign Ncmyx6 = (X4eet6 & O5a7z6);
assign Zo1ov6 = (Jemyx6 & Remyx6);
assign Jemyx6 = (O5a7z6 & Hulov6);
assign Jamyx6 = (~(Zemyx6 | Hfmyx6));
assign Hfmyx6 = (Jsoov6 ? Pfmyx6 : Kkadt6);
assign Jsoov6 = (~(Kboov6 & A4jhw6));
assign Kboov6 = (!Hu0ov6);
assign Hu0ov6 = (~(Xfmyx6 & Cgc7z6[3]));
assign Xfmyx6 = (Cgc7z6[0] & Cgc7z6[1]);
assign Pfmyx6 = (IFLUSH & Iooov6);
assign Zemyx6 = (~(Vjddt6 & O4piw6));
assign T9myx6 = (~(Fgmyx6 & Ngmyx6));
assign Ngmyx6 = (Vgmyx6 & Jamnv6);
assign Vgmyx6 = (Vs9ov6 & Pj1ov6);
assign Fgmyx6 = (~(A9mnv6 | Ierov6));
assign Ierov6 = (!Rihov6);
assign K1p7v6 = (Wj1ov6 ? X0d7z6[2] : Dvc7z6[2]);
assign D1p7v6 = (Wj1ov6 ? X0d7z6[3] : Dvc7z6[3]);
assign W0p7v6 = (Wj1ov6 ? X0d7z6[4] : Dvc7z6[4]);
assign P0p7v6 = (Wj1ov6 ? X0d7z6[5] : Dvc7z6[5]);
assign I0p7v6 = (Wj1ov6 ? X0d7z6[6] : Dvc7z6[6]);
assign B0p7v6 = (Wj1ov6 ? X0d7z6[7] : Dvc7z6[7]);
assign Uzo7v6 = (Wj1ov6 ? X0d7z6[8] : Dvc7z6[8]);
assign Nzo7v6 = (Wj1ov6 ? X0d7z6[9] : Dvc7z6[9]);
assign Gzo7v6 = (Wj1ov6 ? X0d7z6[10] : Dvc7z6[10]);
assign Zyo7v6 = (Wj1ov6 ? X0d7z6[11] : Dvc7z6[11]);
assign Syo7v6 = (Wj1ov6 ? X0d7z6[12] : Dvc7z6[12]);
assign Lyo7v6 = (Wj1ov6 ? X0d7z6[13] : Dvc7z6[13]);
assign Eyo7v6 = (Wj1ov6 ? X0d7z6[14] : Dvc7z6[14]);
assign Xxo7v6 = (Wj1ov6 ? X0d7z6[15] : Dvc7z6[15]);
assign Qxo7v6 = (Wj1ov6 ? X0d7z6[16] : Dvc7z6[16]);
assign Jxo7v6 = (Wj1ov6 ? X0d7z6[17] : Dvc7z6[17]);
assign Cxo7v6 = (Wj1ov6 ? X0d7z6[18] : Dvc7z6[18]);
assign Vwo7v6 = (Wj1ov6 ? X0d7z6[19] : Dvc7z6[19]);
assign Owo7v6 = (Wj1ov6 ? X0d7z6[20] : Dvc7z6[20]);
assign Hwo7v6 = (Wj1ov6 ? X0d7z6[21] : Dvc7z6[21]);
assign Awo7v6 = (Wj1ov6 ? X0d7z6[22] : Dvc7z6[22]);
assign Tvo7v6 = (Wj1ov6 ? X0d7z6[23] : Dvc7z6[23]);
assign Mvo7v6 = (Wj1ov6 ? X0d7z6[24] : Dvc7z6[24]);
assign Fvo7v6 = (Wj1ov6 ? X0d7z6[25] : Dvc7z6[25]);
assign Yuo7v6 = (Wj1ov6 ? X0d7z6[26] : Dvc7z6[26]);
assign Ruo7v6 = (Wj1ov6 ? X0d7z6[27] : Dvc7z6[27]);
assign Kuo7v6 = (Wj1ov6 ? X0d7z6[28] : Dvc7z6[28]);
assign Duo7v6 = (Wj1ov6 ? X0d7z6[29] : Dvc7z6[29]);
assign Wj1ov6 = (Dhmyx6 & F4xnv6);
assign Dhmyx6 = (Lh1ov6 & Lhmyx6);
assign Wto7v6 = (Thmyx6 | Bimyx6);
assign Bimyx6 = (Jimyx6 ? HPROTI[0] : J5n7z6[0]);
assign Thmyx6 = (R2qhw6 | Fe0iw6);
assign Pto7v6 = (Mr9ov6 ? Fopet6 : HPROTI[0]);
assign Ito7v6 = (~(Rimyx6 & Zimyx6));
assign Zimyx6 = (Hjmyx6 & Pjmyx6);
assign Pjmyx6 = (~(Fe0iw6 & K2bdt6));
assign Fe0iw6 = (Jimyx6 & Uclov6);
assign Hjmyx6 = (~(Xjmyx6 & HPROTI[1]));
assign Rimyx6 = (Fkmyx6 & Nkmyx6);
assign Nkmyx6 = (~(R2qhw6 & Hjqnv6));
assign Fkmyx6 = (~(J5n7z6[1] & Y2qhw6));
assign Bto7v6 = (Mr9ov6 ? Empet6 : HPROTI[1]);
assign Uso7v6 = (~(Vkmyx6 & Dlmyx6));
assign Dlmyx6 = (~(J5n7z6[2] & Y2qhw6));
assign Vkmyx6 = (Llmyx6 & Tlmyx6);
assign Tlmyx6 = (~(Xjmyx6 & Bmmyx6));
assign Llmyx6 = (~(R2qhw6 & Yhqnv6));
assign Nso7v6 = (Mr9ov6 ? Dkpet6 : Bmmyx6);
assign Bmmyx6 = (~(Jmmyx6 & Rmmyx6));
assign Rmmyx6 = (~(Zmmyx6 & Hnmyx6));
assign Zmmyx6 = (Pnmyx6 & Xnmyx6);
assign Pnmyx6 = (~(Fomyx6 & Nomyx6));
assign Nomyx6 = (Vomyx6 & Dpmyx6);
assign Dpmyx6 = (Lpmyx6 & Tpmyx6);
assign Lpmyx6 = (Bqmyx6 & Jqmyx6);
assign Vomyx6 = (Rqmyx6 & Zqmyx6);
assign Fomyx6 = (Hrmyx6 & Prmyx6);
assign Prmyx6 = (Xrmyx6 & Fsmyx6);
assign Xrmyx6 = (Nsmyx6 & Vsmyx6);
assign Hrmyx6 = (Bkkiw6 & Dtmyx6);
assign Jmmyx6 = (~(Ltmyx6 & Ttmyx6));
assign Ttmyx6 = (~(Bumyx6 & Jumyx6));
assign Jumyx6 = (~(Rumyx6 & Zumyx6));
assign Bumyx6 = (Xvmyx6 ? Pvmyx6 : Hvmyx6);
assign Gso7v6 = (~(Fwmyx6 & Nwmyx6));
assign Nwmyx6 = (~(J5n7z6[3] & Y2qhw6));
assign Fwmyx6 = (Vwmyx6 & Dxmyx6);
assign Dxmyx6 = (~(Xjmyx6 & Lxmyx6));
assign Vwmyx6 = (~(R2qhw6 & Pgqnv6));
assign Zro7v6 = (Mr9ov6 ? Cipet6 : Lxmyx6);
assign Lxmyx6 = (~(Txmyx6 & Bymyx6));
assign Bymyx6 = (~(Ltmyx6 & Jymyx6));
assign Jymyx6 = (~(Rymyx6 & Zymyx6));
assign Rymyx6 = (Xvmyx6 & Hzmyx6);
assign Hzmyx6 = (~(Pzmyx6 & Xzmyx6));
assign Pzmyx6 = (Pvmyx6 & F0nyx6);
assign Txmyx6 = (~(Hnmyx6 & N0nyx6));
assign Sro7v6 = (~(V0nyx6 & D1nyx6));
assign D1nyx6 = (~(W2n7z6[0] & Y2qhw6));
assign V0nyx6 = (L1nyx6 & T1nyx6);
assign T1nyx6 = (~(Xjmyx6 & B2nyx6));
assign L1nyx6 = (~(R2qhw6 & Gfqnv6));
assign Lro7v6 = (Mr9ov6 ? Bgpet6 : B2nyx6);
assign B2nyx6 = (~(J2nyx6 & R2nyx6));
assign R2nyx6 = (~(Z2nyx6 & Ltmyx6));
assign Z2nyx6 = (Xvmyx6 ? H3nyx6 : Zumyx6);
assign H3nyx6 = (P3nyx6 & Xzmyx6);
assign P3nyx6 = (~(F0nyx6 | Zymyx6));
assign J2nyx6 = (X3nyx6 | Xnmyx6);
assign Ero7v6 = (~(F4nyx6 & N4nyx6));
assign N4nyx6 = (~(W2n7z6[1] & Y2qhw6));
assign F4nyx6 = (V4nyx6 & D5nyx6);
assign D5nyx6 = (~(Xjmyx6 & L5nyx6));
assign Xjmyx6 = (Jimyx6 & Yq9ov6);
assign V4nyx6 = (~(R2qhw6 & Qdqnv6));
assign R2qhw6 = (Jimyx6 & Fbqnv6);
assign Fbqnv6 = (~(T5nyx6 & B6nyx6));
assign Jimyx6 = (!Y2qhw6);
assign Y2qhw6 = (~(J6nyx6 & X02iw6));
assign X02iw6 = (~(R6nyx6 & Z6nyx6));
assign Z6nyx6 = (~(H7nyx6 | Wwonv6));
assign R6nyx6 = (P7nyx6 & X7nyx6);
assign X7nyx6 = (~(F8nyx6 & Bjhxx6));
assign F8nyx6 = (Ven7z6[2] & Osixx6);
assign P7nyx6 = (~(N8nyx6 & Yjonv6));
assign N8nyx6 = (~(V8nyx6 & D9nyx6));
assign D9nyx6 = (B6nyx6 & L9nyx6);
assign V8nyx6 = (T9nyx6 & Banyx6);
assign J6nyx6 = (~(N0qhw6 & Janyx6));
assign Janyx6 = (~(Ranyx6 & V1eiw6));
assign V1eiw6 = (S12iw6 ^ N22iw6);
assign Ranyx6 = (A4qhw6 & O1eiw6);
assign N0qhw6 = (~(Zanyx6 & Hbnyx6));
assign Hbnyx6 = (S12iw6 & O1eiw6);
assign S12iw6 = (~(Pbnyx6 & Xbnyx6));
assign Xbnyx6 = (~(Fcnyx6 | Wwonv6));
assign Wwonv6 = (Yjonv6 & Yq9ov6);
assign Yq9ov6 = (~(Ncnyx6 & Vcnyx6));
assign Vcnyx6 = (~(Woyet6 & T8gxx6));
assign Fcnyx6 = (~(En9ov6 | Ddnyx6));
assign Pbnyx6 = (Ldnyx6 & Tdnyx6);
assign Tdnyx6 = (Cakiw6 | Benyx6);
assign Zanyx6 = (J2eiw6 & N22iw6);
assign N22iw6 = (~(Jenyx6 & Renyx6));
assign Renyx6 = (Zenyx6 & Ddnyx6);
assign Zenyx6 = (~(Bjhxx6 | Djonv6));
assign Jenyx6 = (Ldnyx6 & Hfnyx6);
assign Hfnyx6 = (~(Enonv6 & Yjonv6));
assign Ldnyx6 = (Pfnyx6 & Xfnyx6);
assign Xfnyx6 = (~(Fgnyx6 & Ngnyx6));
assign Fgnyx6 = (Vgnyx6 & Yjonv6);
assign Pfnyx6 = (Luixx6 & Dhnyx6);
assign J2eiw6 = (!A4qhw6);
assign A4qhw6 = (~(Lhnyx6 & Thnyx6));
assign Thnyx6 = (Binyx6 & Luixx6);
assign Binyx6 = (Dhnyx6 & Jinyx6);
assign Lhnyx6 = (Rinyx6 & Zinyx6);
assign Zinyx6 = (~(Yjonv6 & Hjnyx6));
assign Hjnyx6 = (~(Pjnyx6 & Ncnyx6));
assign Ncnyx6 = (~(Xjnyx6 & T5nyx6));
assign Pjnyx6 = (B6nyx6 & Fknyx6);
assign B6nyx6 = (~(Nknyx6 & Vknyx6));
assign Vknyx6 = (~(Xjnyx6 | Woyet6));
assign Xjnyx6 = (!Wp9ov6);
assign Nknyx6 = (Hryet6 & T8gxx6);
assign T8gxx6 = (Dlnyx6 & T5nyx6);
assign Dlnyx6 = (L9nyx6 & En9ov6);
assign Rinyx6 = (~(Rxonv6 & Vudiw6));
assign Vudiw6 = (!L9nyx6);
assign Rxonv6 = (!Ddnyx6);
assign Ddnyx6 = (~(Uclov6 & Yjonv6));
assign Yjonv6 = (~(Llnyx6 & Tlnyx6));
assign Tlnyx6 = (Bjhxx6 | Znn7z6[0]);
assign Bjhxx6 = (Znn7z6[1] & Ozixx6);
assign Llnyx6 = (~(Qakiw6 & Rxixx6));
assign Uclov6 = (T5nyx6 & Bmnyx6);
assign Bmnyx6 = (~(En9ov6 & L9nyx6));
assign L9nyx6 = (~(Jmnyx6 & Rmnyx6));
assign Rmnyx6 = (~(V4myx6 & Zn9ov6));
assign Jmnyx6 = (~(Zmnyx6 | Go9ov6));
assign T5nyx6 = (Banyx6 & Xm9ov6);
assign Banyx6 = (Vgnyx6 & Fknyx6);
assign Fknyx6 = (!Enonv6);
assign Enonv6 = (Hnnyx6 & Vgnyx6);
assign Hnnyx6 = (Pnnyx6 & Xm9ov6);
assign Xm9ov6 = (!Ngnyx6);
assign Pnnyx6 = (~(Uvixx6 & Qm9ov6));
assign Qm9ov6 = (~(Xnnyx6 & Rj9ov6));
assign Vgnyx6 = (Nvixx6 & No9ov6);
assign No9ov6 = (~(Noonv6 & P6u6x6));
assign Noonv6 = (Dkm7z6[1] & Zuixx6);
assign Nvixx6 = (~(Fonyx6 & Dkm7z6[0]));
assign Fonyx6 = (P6u6x6 & Goonv6);
assign Xqo7v6 = (Mr9ov6 ? Aepet6 : L5nyx6);
assign L5nyx6 = (~(Nonyx6 & Vonyx6));
assign Vonyx6 = (~(Dpnyx6 & Lpnyx6));
assign Lpnyx6 = (Bkfnv6 & Zn3nv6);
assign Dpnyx6 = (Njfnv6 & Hnmyx6);
assign Nonyx6 = (~(Tpnyx6 & Ltmyx6));
assign Tpnyx6 = (Bqnyx6 & Jqnyx6);
assign Jqnyx6 = (~(Rqnyx6 & Zqnyx6));
assign Zqnyx6 = (Hrnyx6 & Prnyx6);
assign Prnyx6 = (Xrnyx6 & Fsnyx6);
assign Fsnyx6 = (~(Nsnyx6 & Hwk7z6[16]));
assign Xrnyx6 = (Vsnyx6 & Dtnyx6);
assign Dtnyx6 = (~(Xzmyx6 & Rumyx6));
assign Vsnyx6 = (~(Ltnyx6 & Zlk7z6[16]));
assign Hrnyx6 = (Ttnyx6 & Bunyx6);
assign Bunyx6 = (~(Junyx6 & P6l7z6[16]));
assign Ttnyx6 = (~(Runyx6 & Xgl7z6[16]));
assign Rqnyx6 = (Zunyx6 & Hvnyx6);
assign Hvnyx6 = (Pvnyx6 & Xvnyx6);
assign Xvnyx6 = (~(Fwnyx6 & Frl7z6[16]));
assign Pvnyx6 = (~(Nwnyx6 & N1m7z6[16]));
assign Zunyx6 = (Vwnyx6 & Dxnyx6);
assign Dxnyx6 = (~(Lxnyx6 & Rbk7z6[16]));
assign Vwnyx6 = (~(Txnyx6 & Vbm7z6[16]));
assign Bqnyx6 = (~(Bynyx6 & Pvmyx6));
assign Pvmyx6 = (Jynyx6 & Rynyx6);
assign Rynyx6 = (Zynyx6 & Hznyx6);
assign Hznyx6 = (Pznyx6 & Xznyx6);
assign Xznyx6 = (~(Nwnyx6 & N1m7z6[14]));
assign Pznyx6 = (~(Lxnyx6 & Rbk7z6[14]));
assign Zynyx6 = (F0oyx6 & N0oyx6);
assign N0oyx6 = (~(Junyx6 & P6l7z6[14]));
assign F0oyx6 = (~(Nsnyx6 & Hwk7z6[14]));
assign Jynyx6 = (V0oyx6 & D1oyx6);
assign D1oyx6 = (L1oyx6 & T1oyx6);
assign T1oyx6 = (~(Fwnyx6 & Frl7z6[14]));
assign L1oyx6 = (~(Ltnyx6 & Zlk7z6[14]));
assign V0oyx6 = (B2oyx6 & J2oyx6);
assign J2oyx6 = (~(Txnyx6 & Vbm7z6[14]));
assign B2oyx6 = (~(Runyx6 & Xgl7z6[14]));
assign Bynyx6 = (Rumyx6 & Zumyx6);
assign Zumyx6 = (!Xzmyx6);
assign Xzmyx6 = (R2oyx6 & Z2oyx6);
assign Z2oyx6 = (H3oyx6 & P3oyx6);
assign P3oyx6 = (X3oyx6 & F4oyx6);
assign F4oyx6 = (~(Runyx6 & Xgl7z6[18]));
assign X3oyx6 = (~(Lxnyx6 & Rbk7z6[18]));
assign H3oyx6 = (N4oyx6 & V4oyx6);
assign V4oyx6 = (~(Junyx6 & P6l7z6[18]));
assign N4oyx6 = (~(Nsnyx6 & Hwk7z6[18]));
assign R2oyx6 = (D5oyx6 & L5oyx6);
assign L5oyx6 = (T5oyx6 & B6oyx6);
assign B6oyx6 = (~(Txnyx6 & Vbm7z6[18]));
assign T5oyx6 = (~(Nwnyx6 & N1m7z6[18]));
assign D5oyx6 = (J6oyx6 & R6oyx6);
assign R6oyx6 = (~(Fwnyx6 & Frl7z6[18]));
assign J6oyx6 = (~(Ltnyx6 & Zlk7z6[18]));
assign Rumyx6 = (Z6oyx6 & Zymyx6);
assign Zymyx6 = (H7oyx6 & P7oyx6);
assign P7oyx6 = (X7oyx6 & F8oyx6);
assign F8oyx6 = (N8oyx6 & V8oyx6);
assign V8oyx6 = (~(Nwnyx6 & N1m7z6[15]));
assign N8oyx6 = (~(Lxnyx6 & Rbk7z6[15]));
assign X7oyx6 = (D9oyx6 & L9oyx6);
assign L9oyx6 = (~(Junyx6 & P6l7z6[15]));
assign D9oyx6 = (~(Nsnyx6 & Hwk7z6[15]));
assign H7oyx6 = (T9oyx6 & Baoyx6);
assign Baoyx6 = (Jaoyx6 & Raoyx6);
assign Raoyx6 = (~(Fwnyx6 & Frl7z6[15]));
assign Jaoyx6 = (~(Ltnyx6 & Zlk7z6[15]));
assign T9oyx6 = (Zaoyx6 & Hboyx6);
assign Hboyx6 = (~(Txnyx6 & Vbm7z6[15]));
assign Zaoyx6 = (~(Runyx6 & Xgl7z6[15]));
assign Z6oyx6 = (Xvmyx6 & Hvmyx6);
assign Hvmyx6 = (!F0nyx6);
assign F0nyx6 = (~(Pboyx6 & Xboyx6));
assign Xboyx6 = (Fcoyx6 & Ncoyx6);
assign Ncoyx6 = (Vcoyx6 & Ddoyx6);
assign Ddoyx6 = (~(Nwnyx6 & N1m7z6[17]));
assign Vcoyx6 = (~(Lxnyx6 & Rbk7z6[17]));
assign Fcoyx6 = (Ldoyx6 & Tdoyx6);
assign Tdoyx6 = (~(Junyx6 & P6l7z6[17]));
assign Ldoyx6 = (~(Nsnyx6 & Hwk7z6[17]));
assign Pboyx6 = (Beoyx6 & Jeoyx6);
assign Jeoyx6 = (Reoyx6 & Zeoyx6);
assign Zeoyx6 = (~(Fwnyx6 & Frl7z6[17]));
assign Reoyx6 = (~(Ltnyx6 & Zlk7z6[17]));
assign Beoyx6 = (Hfoyx6 & Pfoyx6);
assign Pfoyx6 = (~(Txnyx6 & Vbm7z6[17]));
assign Hfoyx6 = (~(Runyx6 & Xgl7z6[17]));
assign Xvmyx6 = (Xfoyx6 & Fgoyx6);
assign Fgoyx6 = (Ngoyx6 & Vgoyx6);
assign Vgoyx6 = (Dhoyx6 & Lhoyx6);
assign Lhoyx6 = (~(Runyx6 & Xgl7z6[19]));
assign Dhoyx6 = (~(Lxnyx6 & Rbk7z6[19]));
assign Ngoyx6 = (Thoyx6 & Bioyx6);
assign Bioyx6 = (~(Junyx6 & P6l7z6[19]));
assign Thoyx6 = (~(Nsnyx6 & Hwk7z6[19]));
assign Xfoyx6 = (Jioyx6 & Rioyx6);
assign Rioyx6 = (Zioyx6 & Hjoyx6);
assign Hjoyx6 = (~(Txnyx6 & Vbm7z6[19]));
assign Zioyx6 = (~(Nwnyx6 & N1m7z6[19]));
assign Jioyx6 = (Pjoyx6 & Xjoyx6);
assign Xjoyx6 = (~(Fwnyx6 & Frl7z6[19]));
assign Pjoyx6 = (~(Ltnyx6 & Zlk7z6[19]));
assign Qqo7v6 = (~(Fkoyx6 & Nkoyx6));
assign Nkoyx6 = (~(Jexmz6[0] & K94iw6));
assign Fkoyx6 = (Vkoyx6 & Dloyx6);
assign Dloyx6 = (~(Lloyx6 & Td9ov6));
assign Td9ov6 = (~(Tloyx6 & Bmoyx6));
assign Bmoyx6 = (Jmoyx6 & Rmoyx6);
assign Rmoyx6 = (~(Zmoyx6 & Orwnv6));
assign Orwnv6 = (~(Hnoyx6 & Pnoyx6));
assign Pnoyx6 = (~(Xnoyx6 & Uea7z6));
assign Uea7z6 = (~(Fooyx6 & Nooyx6));
assign Nooyx6 = (~(HRDATAD[0] & Qln7z6[0]));
assign Fooyx6 = (~(HRDATAS[0] & Qln7z6[1]));
assign Hnoyx6 = (Vooyx6 & Dpoyx6);
assign Dpoyx6 = (~(Lpoyx6 & Tronv6));
assign Tronv6 = (Euonv6 | Zuonv6);
assign Zuonv6 = (~(S7n7z6[1] | S7n7z6[0]));
assign Euonv6 = (!Evadt6);
assign Vooyx6 = (~(Tim7z6[0] & Tpoyx6));
assign Jmoyx6 = (Bqoyx6 | Vrwnv6);
assign Vrwnv6 = (Jqoyx6 & Rqoyx6);
assign Rqoyx6 = (Zqoyx6 & Hroyx6);
assign Hroyx6 = (Proyx6 & Xroyx6);
assign Xroyx6 = (~(Fsoyx6 & Nsoyx6));
assign Fsoyx6 = (Klo7z6[5] & Vsoyx6);
assign Vsoyx6 = (~(Dtoyx6 & Ltoyx6));
assign Ltoyx6 = (Ttoyx6 & Buoyx6);
assign Buoyx6 = (Juoyx6 & Ruoyx6);
assign Ruoyx6 = (~(Hyj7z6[0] & Rbk7z6[0]));
assign Juoyx6 = (~(Hyj7z6[1] & Zlk7z6[0]));
assign Ttoyx6 = (Zuoyx6 & Hvoyx6);
assign Hvoyx6 = (~(Hyj7z6[2] & Hwk7z6[0]));
assign Zuoyx6 = (~(Hyj7z6[3] & P6l7z6[0]));
assign Dtoyx6 = (Pvoyx6 & Xvoyx6);
assign Xvoyx6 = (Fwoyx6 & Nwoyx6);
assign Nwoyx6 = (~(Hyj7z6[4] & Xgl7z6[0]));
assign Fwoyx6 = (~(Hyj7z6[5] & Frl7z6[0]));
assign Pvoyx6 = (Vwoyx6 & Dxoyx6);
assign Dxoyx6 = (~(Hyj7z6[6] & N1m7z6[0]));
assign Vwoyx6 = (~(Hyj7z6[7] & Vbm7z6[0]));
assign Proyx6 = (Lxoyx6 & Txoyx6);
assign Lxoyx6 = (Byoyx6 | Jyoyx6);
assign Jyoyx6 = (Ti2nz6[2] ? Zyoyx6 : Ryoyx6);
assign Ryoyx6 = (~(Hzoyx6 & Ti2nz6[0]));
assign Hzoyx6 = (~(Pzoyx6 | Ti2nz6[3]));
assign Pzoyx6 = (!Xzoyx6);
assign Byoyx6 = (~(Ti2nz6[1] & F0pyx6));
assign Zqoyx6 = (N0pyx6 & V0pyx6);
assign V0pyx6 = (~(D1pyx6 & L1pyx6));
assign L1pyx6 = (~(T1pyx6 & B2pyx6));
assign B2pyx6 = (J2pyx6 & R2pyx6);
assign R2pyx6 = (Z2pyx6 & H3pyx6);
assign H3pyx6 = (P3pyx6 & X3pyx6);
assign X3pyx6 = (F4pyx6 | N4pyx6);
assign F4pyx6 = (~(V4pyx6 & Gthiw6));
assign P3pyx6 = (D5pyx6 & L5pyx6);
assign D5pyx6 = (~(T5pyx6 & B6pyx6));
assign T5pyx6 = (J6pyx6 & R6pyx6);
assign J6pyx6 = (~(Z6pyx6 & H7pyx6));
assign H7pyx6 = (~(P7pyx6 & X7pyx6));
assign X7pyx6 = (F8pyx6 & Xfymz6[9]);
assign F8pyx6 = (~(Xfymz6[10] | Xfymz6[11]));
assign P7pyx6 = (N8pyx6 & Xfymz6[8]);
assign Z6pyx6 = (~(V8pyx6 & At67v6));
assign V8pyx6 = (D9pyx6 & L9pyx6);
assign Z2pyx6 = (T9pyx6 & Bapyx6);
assign Bapyx6 = (~(Jdymz6[0] & Sjd8x6));
assign T9pyx6 = (~(Zt67v6 & Xm4xx6));
assign J2pyx6 = (Japyx6 & Rapyx6);
assign Rapyx6 = (Zapyx6 & Hbpyx6);
assign Hbpyx6 = (~(Zshiw6 & N8pyx6));
assign Zapyx6 = (~(Pbpyx6 & Xbpyx6));
assign Japyx6 = (Fcpyx6 & Ncpyx6);
assign Ncpyx6 = (~(Gh77z6 & Vcpyx6));
assign Fcpyx6 = (~(Biymz6[0] & Ddpyx6));
assign T1pyx6 = (Ldpyx6 & Tdpyx6);
assign Tdpyx6 = (Bepyx6 & Jepyx6);
assign Jepyx6 = (Repyx6 & Zepyx6);
assign Zepyx6 = (~(Ojymz6[0] & Hfpyx6));
assign Repyx6 = (Pfpyx6 & Xfpyx6);
assign Xfpyx6 = (~(Fgpyx6 & Wy67v6));
assign Pfpyx6 = (~(Sgymz6[0] & Ngpyx6));
assign Bepyx6 = (Vgpyx6 & Dhpyx6);
assign Dhpyx6 = (~(Kmymz6[0] & Lhpyx6));
assign Vgpyx6 = (~(Unymz6[0] & Thpyx6));
assign Ldpyx6 = (Bipyx6 & Jipyx6);
assign Jipyx6 = (Ripyx6 & Zipyx6);
assign Zipyx6 = (~(Fjd7v6 & Hjpyx6));
assign Bipyx6 = (Pjpyx6 & Xjpyx6);
assign N0pyx6 = (Fkpyx6 & Nkpyx6);
assign Nkpyx6 = (~(Vkpyx6 & Dlpyx6));
assign Vkpyx6 = (~(Llpyx6 & Tlpyx6));
assign Fkpyx6 = (~(Bmpyx6 & Jmpyx6));
assign Jmpyx6 = (~(Rmpyx6 & Zmpyx6));
assign Zmpyx6 = (Hnpyx6 & Pnpyx6);
assign Pnpyx6 = (Xnpyx6 & Fopyx6);
assign Xnpyx6 = (Nopyx6 & Vopyx6);
assign Hnpyx6 = (Dppyx6 & Lppyx6);
assign Lppyx6 = (~(Tppyx6 & Bqpyx6));
assign Bqpyx6 = (~(Jqpyx6 & Rqpyx6));
assign Rqpyx6 = (~(Yvhiw6 & Zqpyx6));
assign Zqpyx6 = (Txhyx6 | W197z6);
assign Jqpyx6 = (~(Hrpyx6 & Prpyx6));
assign Prpyx6 = (!Y097z6);
assign Dppyx6 = (Xrpyx6 & Fspyx6);
assign Fspyx6 = (~(Nspyx6 & Iy1nz6[0]));
assign Xrpyx6 = (~(Jke7v6 & Vspyx6));
assign Vspyx6 = (~(Dtpyx6 & Ltpyx6));
assign Ltpyx6 = (~(Nl1nz6[0] & Mwhiw6));
assign Dtpyx6 = (~(Eee7v6 & Hiiiw6));
assign Rmpyx6 = (Ttpyx6 & Bupyx6);
assign Bupyx6 = (Jupyx6 & Rupyx6);
assign Rupyx6 = (~(Oo1nz6[0] & Ri3yx6));
assign Jupyx6 = (Zupyx6 & Hvpyx6);
assign Hvpyx6 = (~(Jw1nz6[0] & Pvpyx6));
assign Zupyx6 = (~(Pk1nz6[0] & Xvpyx6));
assign Ttpyx6 = (Fwpyx6 & Nwpyx6);
assign Fwpyx6 = (Vwpyx6 & Dxpyx6);
assign Dxpyx6 = (~(Au1nz6[0] & N82yx6));
assign Jqoyx6 = (Lxpyx6 & Txpyx6);
assign Txpyx6 = (Bypyx6 & Jypyx6);
assign Jypyx6 = (~(Klo7z6[1] & Rypyx6));
assign Rypyx6 = (~(Zypyx6 & Hzpyx6));
assign Hzpyx6 = (Pzpyx6 & Xzpyx6);
assign Xzpyx6 = (F0qyx6 & N0qyx6);
assign N0qyx6 = (V0qyx6 & D1qyx6);
assign D1qyx6 = (~(Kfq7z6[0] & S7hiw6));
assign V0qyx6 = (L1qyx6 & T1qyx6);
assign L1qyx6 = (~(B2qyx6 & J2qyx6));
assign F0qyx6 = (R2qyx6 & Z2qyx6);
assign Z2qyx6 = (~(Hhq7z6[0] & Ydliw6));
assign R2qyx6 = (H3qyx6 & P3qyx6);
assign P3qyx6 = (~(Tbq7z6[0] & Qsgiw6));
assign H3qyx6 = (~(Pdq7z6[0] & Oka8x6));
assign Pzpyx6 = (X3qyx6 & F4qyx6);
assign F4qyx6 = (N4qyx6 & V4qyx6);
assign V4qyx6 = (~(D5qyx6 & Bqp7z6[0]));
assign N4qyx6 = (L5qyx6 & T5qyx6);
assign T5qyx6 = (~(Cjq7z6[0] & Cza8x6));
assign L5qyx6 = (~(Qb4ft6 & B6qyx6));
assign X3qyx6 = (J6qyx6 & R6qyx6);
assign R6qyx6 = (~(Z6qyx6 & Gop7z6[0]));
assign J6qyx6 = (~(H7qyx6 & Rip7z6[0]));
assign Zypyx6 = (P7qyx6 & X7qyx6);
assign X7qyx6 = (F8qyx6 & N8qyx6);
assign N8qyx6 = (V8qyx6 & D9qyx6);
assign D9qyx6 = (~(L9qyx6 & E6p7z6[0]));
assign V8qyx6 = (T9qyx6 & Baqyx6);
assign Baqyx6 = (~(P3a8x6 & Hmp7z6[0]));
assign T9qyx6 = (~(Ua9ov6 & Sgp7z6[0]));
assign F8qyx6 = (Jaqyx6 & Raqyx6);
assign Raqyx6 = (~(Zaqyx6 & G0q7z6[0]));
assign Jaqyx6 = (Hbqyx6 & Pbqyx6);
assign Pbqyx6 = (~(Xbqyx6 & Q8p7z6[0]));
assign Hbqyx6 = (~(Fcqyx6 & B2q7z6[0]));
assign P7qyx6 = (Ncqyx6 & Vcqyx6);
assign Vcqyx6 = (Ddqyx6 & Ldqyx6);
assign Ldqyx6 = (~(Tdqyx6 & Mkp7z6[0]));
assign Ddqyx6 = (Beqyx6 & Jeqyx6);
assign Jeqyx6 = (~(Nao7x6 & I7p7z6[0]));
assign Beqyx6 = (~(Q0a8x6 & Hyp7z6[0]));
assign Ncqyx6 = (Reqyx6 & Zeqyx6);
assign Zeqyx6 = (~(U9p7z6[0] & Hfqyx6));
assign Bypyx6 = (Pfqyx6 & Xfqyx6);
assign Xfqyx6 = (~(Fgqyx6 & Ngqyx6));
assign Fgqyx6 = (~(Vgqyx6 & Dhqyx6));
assign Dhqyx6 = (Lhqyx6 & Thqyx6);
assign Thqyx6 = (Biqyx6 & Jiqyx6);
assign Jiqyx6 = (Riqyx6 & Ziqyx6);
assign Ziqyx6 = (Hjqyx6 & Pjqyx6);
assign Riqyx6 = (Xjqyx6 & Fkqyx6);
assign Xjqyx6 = (~(Nkqyx6 & Vkqyx6));
assign Nkqyx6 = (Dlqyx6 & Llqyx6);
assign Llqyx6 = (~(Tlqyx6 & Bmqyx6));
assign Bmqyx6 = (~(Jmqyx6 & Doadt6));
assign Biqyx6 = (Rmqyx6 & Zmqyx6);
assign Zmqyx6 = (~(Aqadt6 & Hnqyx6));
assign Rmqyx6 = (Pnqyx6 & Xnqyx6);
assign Xnqyx6 = (~(Foqyx6 & A8cet6));
assign Foqyx6 = (Noqyx6 & Voqyx6);
assign Pnqyx6 = (~(Bxi7z6[0] & Dpqyx6));
assign Lhqyx6 = (Lpqyx6 & Tpqyx6);
assign Tpqyx6 = (Bqqyx6 & Jqqyx6);
assign Jqqyx6 = (~(H1j7z6[0] & Rqqyx6));
assign Bqqyx6 = (Zqqyx6 & Hrqyx6);
assign Hrqyx6 = (~(Prqyx6 & Z3j7z6[0]));
assign Zqqyx6 = (~(A0j7z6[0] & Xrqyx6));
assign Lpqyx6 = (Fsqyx6 & Nsqyx6);
assign Nsqyx6 = (~(Bzi7z6[0] & Vsqyx6));
assign Fsqyx6 = (Dtqyx6 & Ltqyx6);
assign Ltqyx6 = (~(Zodet6 & Ttqyx6));
assign Dtqyx6 = (~(Buqyx6 & A0fet6));
assign Vgqyx6 = (Juqyx6 & Ruqyx6);
assign Ruqyx6 = (Zuqyx6 & Hvqyx6);
assign Hvqyx6 = (Pvqyx6 & Xvqyx6);
assign Xvqyx6 = (~(Dri7z6[0] & Fwqyx6));
assign Pvqyx6 = (Nwqyx6 & Vwqyx6);
assign Vwqyx6 = (~(Dxqyx6 & Nob7z6[0]));
assign Nwqyx6 = (~(Wui7z6[0] & Lxqyx6));
assign Zuqyx6 = (Txqyx6 & Byqyx6);
assign Byqyx6 = (~(Jyqyx6 & G5j7z6[0]));
assign Txqyx6 = (Ryqyx6 & Zyqyx6);
assign Zyqyx6 = (~(Bwi7z6[0] & Hzqyx6));
assign Ryqyx6 = (~(Pzqyx6 & G5j7z6[32]));
assign Juqyx6 = (Xzqyx6 & F0ryx6);
assign F0ryx6 = (N0ryx6 & V0ryx6);
assign V0ryx6 = (~(D1ryx6 & Ohj7z6[32]));
assign N0ryx6 = (L1ryx6 & T1ryx6);
assign T1ryx6 = (~(B2ryx6 & M6j7z6[32]));
assign L1ryx6 = (~(J2ryx6 & M6j7z6[0]));
assign Xzqyx6 = (R2ryx6 & Z2ryx6);
assign R2ryx6 = (H3ryx6 & P3ryx6);
assign P3ryx6 = (~(X3ryx6 & Ohj7z6[0]));
assign H3ryx6 = (~(STCALIB[0] & F4ryx6));
assign Pfqyx6 = (~(Klo7z6[2] & N4ryx6));
assign N4ryx6 = (~(V4ryx6 & D5ryx6));
assign D5ryx6 = (L5ryx6 & T5ryx6);
assign T5ryx6 = (B6ryx6 & J6ryx6);
assign J6ryx6 = (~(Q3kiw6 & Zy1ft6));
assign B6ryx6 = (~(R6ryx6 | Z6ryx6));
assign L5ryx6 = (H7ryx6 & P7ryx6);
assign P7ryx6 = (~(Nn1ft6 & K7kiw6));
assign H7ryx6 = (X7ryx6 & F8ryx6);
assign F8ryx6 = (~(Tk1ft6 & M8kiw6));
assign X7ryx6 = (~(Jj1ft6 & H9kiw6));
assign V4ryx6 = (N8ryx6 & V8ryx6);
assign V8ryx6 = (D9ryx6 & L9ryx6);
assign L9ryx6 = (~(Rr1ft6 & U5kiw6));
assign D9ryx6 = (T9ryx6 & Baryx6);
assign Baryx6 = (~(Xo1ft6 & W6kiw6));
assign T9ryx6 = (~(Dm1ft6 & Y7kiw6));
assign N8ryx6 = (Jaryx6 & Raryx6);
assign Raryx6 = (~(Iv1ft6 & G5kiw6));
assign Jaryx6 = (~(Hq1ft6 & I6kiw6));
assign Lxpyx6 = (Zaryx6 & Hbryx6);
assign Zaryx6 = (Pbryx6 & Xbryx6);
assign Xbryx6 = (~(Klo7z6[0] & Fcryx6));
assign Fcryx6 = (~(Ncryx6 & Vcryx6));
assign Vcryx6 = (Ddryx6 & Ldryx6);
assign Ldryx6 = (~(Tdryx6 | Beryx6));
assign Ddryx6 = (Jeryx6 & Reryx6);
assign Reryx6 = (~(Zeryx6 & Hfryx6));
assign Zeryx6 = (Pfryx6 ? Ies7z6[0] : Rj27v6);
assign Jeryx6 = (~(Xfryx6 & Fgryx6));
assign Xfryx6 = (~(Ngryx6 & Vgryx6));
assign Vgryx6 = (~(Dhryx6 & Lhryx6));
assign Lhryx6 = (~(Thryx6 | Zfs7z6[11]));
assign Thryx6 = (Zfs7z6[7] | Zfs7z6[9]);
assign Dhryx6 = (~(I96ft6 | Zfs7z6[10]));
assign Ngryx6 = (~(Biryx6 & Jiryx6));
assign Jiryx6 = (~(Riryx6 | Zqbyx6));
assign Zqbyx6 = (Eee7v6 ? Ziryx6 : Lxhyx6);
assign Lxhyx6 = (Hae7v6 ? Pjryx6 : Hjryx6);
assign Pjryx6 = (~(Xjryx6 & Gl5ov6));
assign Xjryx6 = (~(Pp1nz6[1] & Pp1nz6[0]));
assign Hjryx6 = (Fkryx6 & Nkryx6);
assign Nkryx6 = (~(Juhyx6 ^ Pb3yx6));
assign Pb3yx6 = (~(Xb3yx6 ^ Hi1nz6[0]));
assign Juhyx6 = (Ruhyx6 ^ U81nz6[0]);
assign Fkryx6 = (Vkryx6 & Dlryx6);
assign Dlryx6 = (U81nz6[2] ^ Hi1nz6[2]);
assign Vkryx6 = (Ruhyx6 ^ Xb3yx6);
assign Xb3yx6 = (Y9h7v6 ^ Hi1nz6[2]);
assign Ruhyx6 = (U81nz6[1] ^ U81nz6[2]);
assign Biryx6 = (Llryx6 & Mm27v6);
assign Ncryx6 = (Tlryx6 & Bmryx6);
assign Bmryx6 = (Jmryx6 & Rmryx6);
assign Rmryx6 = (~(Scs7z6[0] & Zmryx6));
assign Jmryx6 = (Hnryx6 | Riryx6);
assign Tlryx6 = (Pnryx6 & Xnryx6);
assign Xnryx6 = (~(Foryx6 & Ig27v6));
assign Pbryx6 = (~(Noryx6 & Phget6));
assign Tloyx6 = (Voryx6 & Dpryx6);
assign Dpryx6 = (~(HRDATAS[0] & Ad47x6));
assign Voryx6 = (~(HRDATAD[0] & Mc47x6));
assign Vkoyx6 = (~(Lpryx6 & I8r7x6));
assign Jqo7v6 = (~(Tpryx6 & Bqryx6));
assign Bqryx6 = (~(Jexmz6[1] & K94iw6));
assign Tpryx6 = (Jqryx6 & Rqryx6);
assign Rqryx6 = (~(Lloyx6 & Ex77x6));
assign Ex77x6 = (~(Zqryx6 & Hrryx6));
assign Hrryx6 = (Prryx6 & Xrryx6);
assign Xrryx6 = (Bqoyx6 | Dud7x6);
assign Dud7x6 = (Fsryx6 & Nsryx6);
assign Nsryx6 = (Vsryx6 & Dtryx6);
assign Dtryx6 = (Ltryx6 & Ttryx6);
assign Ttryx6 = (Buryx6 & Juryx6);
assign Juryx6 = (~(Ruryx6 & Nsoyx6));
assign Ruryx6 = (Klo7z6[5] & Zuryx6);
assign Zuryx6 = (~(Hvryx6 & Pvryx6));
assign Pvryx6 = (Xvryx6 & Fwryx6);
assign Fwryx6 = (Nwryx6 & Vwryx6);
assign Vwryx6 = (~(Hyj7z6[0] & Rbk7z6[1]));
assign Nwryx6 = (~(Hyj7z6[1] & Zlk7z6[1]));
assign Xvryx6 = (Dxryx6 & Lxryx6);
assign Lxryx6 = (~(Hyj7z6[2] & Hwk7z6[1]));
assign Dxryx6 = (~(Hyj7z6[3] & P6l7z6[1]));
assign Hvryx6 = (Txryx6 & Byryx6);
assign Byryx6 = (Jyryx6 & Ryryx6);
assign Ryryx6 = (~(Hyj7z6[4] & Xgl7z6[1]));
assign Jyryx6 = (~(Hyj7z6[5] & Frl7z6[1]));
assign Txryx6 = (Zyryx6 & Hzryx6);
assign Hzryx6 = (~(Hyj7z6[6] & N1m7z6[1]));
assign Zyryx6 = (~(Hyj7z6[7] & Vbm7z6[1]));
assign Buryx6 = (~(Pzryx6 & Tdryx6));
assign Tdryx6 = (Xzryx6 & F0syx6);
assign F0syx6 = (N0syx6 & Zfs7z6[8]);
assign N0syx6 = (V0syx6 & D1syx6);
assign Xzryx6 = (Or27v6 & Llryx6);
assign Pzryx6 = (Klo7z6[0] & L1syx6);
assign Ltryx6 = (T1syx6 & B2syx6);
assign B2syx6 = (~(J2syx6 & R6ryx6));
assign J2syx6 = (Klo7z6[2] & R2syx6);
assign T1syx6 = (~(Bmpyx6 & Z2syx6));
assign Z2syx6 = (~(H3syx6 & P3syx6));
assign P3syx6 = (X3syx6 & F4syx6);
assign F4syx6 = (N4syx6 & V4syx6);
assign N4syx6 = (~(Nspyx6 & Iy1nz6[1]));
assign X3syx6 = (D5syx6 & L5syx6);
assign L5syx6 = (~(Jke7v6 & T5syx6));
assign T5syx6 = (~(B6syx6 & J6syx6));
assign J6syx6 = (~(Nl1nz6[1] & Mwhiw6));
assign Mwhiw6 = (R6syx6 & Z6syx6);
assign Z6syx6 = (~(J02nz6[11] | J02nz6[9]));
assign R6syx6 = (Mhiiw6 & H7syx6);
assign Mhiiw6 = (P7syx6 & X7syx6);
assign X7syx6 = (F8syx6 & J02nz6[6]);
assign F8syx6 = (~(J02nz6[3] | J02nz6[8]));
assign P7syx6 = (N8syx6 & Yvhiw6);
assign B6syx6 = (~(Hae7v6 & Hiiiw6));
assign Hiiiw6 = (V8syx6 & D9syx6);
assign D9syx6 = (L9syx6 & T9syx6);
assign T9syx6 = (!J02nz6[7]);
assign V8syx6 = (Basyx6 & Imiiw6);
assign D5syx6 = (Jasyx6 | B63yx6);
assign H3syx6 = (Rasyx6 & Nwpyx6);
assign Rasyx6 = (Zasyx6 & Hbsyx6);
assign Hbsyx6 = (~(Jw1nz6[1] & Pvpyx6));
assign Zasyx6 = (~(Pk1nz6[1] & Xvpyx6));
assign Vsryx6 = (Pbsyx6 & Xbsyx6);
assign Xbsyx6 = (Fcsyx6 & Ncsyx6);
assign Ncsyx6 = (~(Vcsyx6 & Dlpyx6));
assign Vcsyx6 = (~(Ddsyx6 & Ldsyx6));
assign Fcsyx6 = (~(Tdsyx6 & Ngqyx6));
assign Tdsyx6 = (~(Besyx6 & Jesyx6));
assign Jesyx6 = (Resyx6 & Zesyx6);
assign Zesyx6 = (Hfsyx6 & Pfsyx6);
assign Pfsyx6 = (Xfsyx6 & Fgsyx6);
assign Fgsyx6 = (~(Ngsyx6 & Vgsyx6));
assign Vgsyx6 = (Jmqyx6 & O7adt6);
assign Ngsyx6 = (Vkqyx6 & Dlqyx6);
assign Xfsyx6 = (Dhsyx6 & Pjqyx6);
assign Hfsyx6 = (Lhsyx6 & Thsyx6);
assign Thsyx6 = (~(Bxi7z6[1] & Dpqyx6));
assign Lhsyx6 = (Bisyx6 & Jisyx6);
assign Jisyx6 = (~(Risyx6 & Byi7z6[1]));
assign Risyx6 = (Zisyx6 & Hjsyx6);
assign Bisyx6 = (~(Voqyx6 & Pjsyx6));
assign Pjsyx6 = (~(Xjsyx6 & Fksyx6));
assign Fksyx6 = (~(Nksyx6 & D5cet6));
assign Xjsyx6 = (~(E9cet6 & Noqyx6));
assign Resyx6 = (Vksyx6 & Dlsyx6);
assign Dlsyx6 = (Llsyx6 & Tlsyx6);
assign Tlsyx6 = (~(A0j7z6[1] & Xrqyx6));
assign Llsyx6 = (Bmsyx6 & Jmsyx6);
assign Jmsyx6 = (~(O6cet6 & Hnqyx6));
assign Bmsyx6 = (~(Prqyx6 & Z3j7z6[1]));
assign Vksyx6 = (Rmsyx6 & Zmsyx6);
assign Zmsyx6 = (~(Bzi7z6[1] & Vsqyx6));
assign Rmsyx6 = (Hnsyx6 & Pnsyx6);
assign Pnsyx6 = (~(H1j7z6[1] & Rqqyx6));
assign Hnsyx6 = (~(Buqyx6 & Opeet6));
assign Besyx6 = (Xnsyx6 & Fosyx6);
assign Fosyx6 = (Nosyx6 & Vosyx6);
assign Vosyx6 = (Dpsyx6 & Lpsyx6);
assign Lpsyx6 = (~(Dri7z6[1] & Fwqyx6));
assign Dpsyx6 = (Tpsyx6 & Bqsyx6);
assign Bqsyx6 = (~(Dxqyx6 & Nob7z6[1]));
assign Tpsyx6 = (~(Wui7z6[1] & Lxqyx6));
assign Nosyx6 = (Jqsyx6 & Rqsyx6);
assign Rqsyx6 = (~(Jyqyx6 & G5j7z6[1]));
assign Jqsyx6 = (Zqsyx6 & Hrsyx6);
assign Hrsyx6 = (~(Bwi7z6[1] & Hzqyx6));
assign Zqsyx6 = (~(Pzqyx6 & G5j7z6[33]));
assign Xnsyx6 = (Prsyx6 & Xrsyx6);
assign Xrsyx6 = (Fssyx6 & Nssyx6);
assign Nssyx6 = (~(D1ryx6 & Ohj7z6[33]));
assign Fssyx6 = (Vssyx6 & Dtsyx6);
assign Dtsyx6 = (~(B2ryx6 & M6j7z6[33]));
assign Vssyx6 = (~(J2ryx6 & M6j7z6[1]));
assign Prsyx6 = (Ltsyx6 & Ttsyx6);
assign Ttsyx6 = (~(X3ryx6 & Ohj7z6[1]));
assign Ltsyx6 = (~(STCALIB[1] & F4ryx6));
assign Pbsyx6 = (Busyx6 & Jusyx6);
assign Jusyx6 = (~(D1pyx6 & Rusyx6));
assign Rusyx6 = (~(Zusyx6 & Hvsyx6));
assign Hvsyx6 = (Pvsyx6 & Xvsyx6);
assign Xvsyx6 = (Fwsyx6 & Nwsyx6);
assign Nwsyx6 = (~(Vwsyx6 & Xu67v6));
assign Vwsyx6 = (Zshiw6 & N8pyx6);
assign Fwsyx6 = (Dxsyx6 & Qid8x6);
assign Dxsyx6 = (~(Lxsyx6 & Txsyx6));
assign Txsyx6 = (Xm4xx6 & Bysyx6);
assign Bysyx6 = (!W197z6);
assign Lxsyx6 = (C477v6 & X14xx6);
assign X14xx6 = (!Jysyx6);
assign Pvsyx6 = (Rysyx6 & Zysyx6);
assign Zysyx6 = (~(Biymz6[1] & Ddpyx6));
assign Rysyx6 = (Hzsyx6 & Pzsyx6);
assign Pzsyx6 = (~(Jdymz6[1] & Sjd8x6));
assign Hzsyx6 = (~(Wd77z6 & Vcpyx6));
assign Zusyx6 = (Xzsyx6 & F0tyx6);
assign F0tyx6 = (N0tyx6 & V0tyx6);
assign V0tyx6 = (~(Kmymz6[1] & Lhpyx6));
assign N0tyx6 = (D1tyx6 & L1tyx6);
assign L1tyx6 = (~(Sgymz6[1] & Ngpyx6));
assign D1tyx6 = (~(Ojymz6[1] & Hfpyx6));
assign Xzsyx6 = (T1tyx6 & Xjpyx6);
assign T1tyx6 = (B2tyx6 & J2tyx6);
assign J2tyx6 = (~(Unymz6[1] & Thpyx6));
assign B2tyx6 = (~(Hcymz6[1] & Hjpyx6));
assign Busyx6 = (~(Klo7z6[1] & R2tyx6));
assign R2tyx6 = (~(Z2tyx6 & H3tyx6));
assign H3tyx6 = (P3tyx6 & X3tyx6);
assign X3tyx6 = (F4tyx6 & N4tyx6);
assign N4tyx6 = (V4tyx6 & D5tyx6);
assign D5tyx6 = (~(Pdq7z6[1] & Oka8x6));
assign V4tyx6 = (L5tyx6 & T5tyx6);
assign T5tyx6 = (~(Kfq7z6[1] & S7hiw6));
assign L5tyx6 = (~(Tbq7z6[1] & Qsgiw6));
assign F4tyx6 = (B6tyx6 & J6tyx6);
assign J6tyx6 = (~(R6tyx6 & Z6tyx6));
assign B6tyx6 = (H7tyx6 & P7tyx6);
assign P7tyx6 = (~(Hhq7z6[1] & Ydliw6));
assign H7tyx6 = (~(Cjq7z6[1] & Cza8x6));
assign P3tyx6 = (X7tyx6 & F8tyx6);
assign F8tyx6 = (N8tyx6 & V8tyx6);
assign V8tyx6 = (~(D5qyx6 & Bqp7z6[1]));
assign N8tyx6 = (D9tyx6 & L9tyx6);
assign L9tyx6 = (~(T9tyx6 & Aw77z6));
assign D9tyx6 = (~(Y7q7z6[0] & B6qyx6));
assign X7tyx6 = (Batyx6 & Jatyx6);
assign Jatyx6 = (~(Z6qyx6 & Gop7z6[1]));
assign Batyx6 = (~(H7qyx6 & Rip7z6[1]));
assign Z2tyx6 = (Ratyx6 & Zatyx6);
assign Zatyx6 = (Hbtyx6 & Pbtyx6);
assign Pbtyx6 = (Xbtyx6 & Fctyx6);
assign Fctyx6 = (~(L9qyx6 & E6p7z6[1]));
assign Xbtyx6 = (Nctyx6 & Vctyx6);
assign Vctyx6 = (~(Hmp7z6[1] & P3a8x6));
assign Nctyx6 = (~(Sgp7z6[1] & Ua9ov6));
assign Hbtyx6 = (Ddtyx6 & Ldtyx6);
assign Ldtyx6 = (~(Zaqyx6 & G0q7z6[1]));
assign Ddtyx6 = (Tdtyx6 & Betyx6);
assign Betyx6 = (~(Xbqyx6 & Q8p7z6[1]));
assign Tdtyx6 = (~(Fcqyx6 & B2q7z6[1]));
assign Ratyx6 = (Jetyx6 & Retyx6);
assign Retyx6 = (Zetyx6 & Hftyx6);
assign Hftyx6 = (~(Tdqyx6 & Mkp7z6[1]));
assign Zetyx6 = (Pftyx6 & Xftyx6);
assign Xftyx6 = (~(I7p7z6[1] & Nao7x6));
assign Pftyx6 = (~(Hyp7z6[1] & Q0a8x6));
assign Jetyx6 = (Fgtyx6 & Ngtyx6);
assign Ngtyx6 = (~(U9p7z6[1] & Hfqyx6));
assign Fsryx6 = (Vgtyx6 & Dhtyx6);
assign Dhtyx6 = (Lhtyx6 & Thtyx6);
assign Thtyx6 = (Bityx6 & Jityx6);
assign Jityx6 = (~(Weget6 & Noryx6));
assign Bityx6 = (~(Scs7z6[1] & Rityx6));
assign Lhtyx6 = (Zityx6 & Hjtyx6);
assign Hjtyx6 = (~(Oo1nz6[1] & Pjtyx6));
assign Zityx6 = (~(Au1nz6[1] & Xjtyx6));
assign Vgtyx6 = (Fktyx6 & Nktyx6);
assign Nktyx6 = (Vktyx6 & Dltyx6);
assign Dltyx6 = (~(Ci6ft6 & Lltyx6));
assign Vktyx6 = (~(Ies7z6[1] & Tltyx6));
assign Fktyx6 = (Bmtyx6 & Hbryx6);
assign Hbryx6 = (Jmtyx6 & Rmtyx6);
assign Rmtyx6 = (~(F0pyx6 & Zmtyx6));
assign Zmtyx6 = (~(Hntyx6 & Pntyx6));
assign Hntyx6 = (Xntyx6 & Fotyx6);
assign Jmtyx6 = (Notyx6 & Votyx6);
assign Notyx6 = (~(Hyj7z6[3] & Dlpyx6));
assign Prryx6 = (~(Zmoyx6 & Kud7x6));
assign Kud7x6 = (~(Dptyx6 & Lptyx6));
assign Lptyx6 = (~(Xnoyx6 & Mea7z6));
assign Mea7z6 = (~(Tptyx6 & Bqtyx6));
assign Bqtyx6 = (~(HRDATAD[1] & Qln7z6[0]));
assign Tptyx6 = (~(HRDATAS[1] & Qln7z6[1]));
assign Dptyx6 = (~(Tim7z6[1] & Tpoyx6));
assign Zqryx6 = (Jqtyx6 & Rqtyx6);
assign Rqtyx6 = (~(HRDATAS[1] & Ad47x6));
assign Jqtyx6 = (~(HRDATAD[1] & Mc47x6));
assign Jqryx6 = (~(Lpryx6 & L7q7x6));
assign Cqo7v6 = (~(Zqtyx6 & Hrtyx6));
assign Hrtyx6 = (~(Jexmz6[2] & K94iw6));
assign Zqtyx6 = (Prtyx6 & Xrtyx6);
assign Xrtyx6 = (~(Lloyx6 & Icfov6));
assign Icfov6 = (~(Fstyx6 & Nstyx6));
assign Nstyx6 = (Vstyx6 & Dttyx6);
assign Dttyx6 = (Bqoyx6 | Xxd7x6);
assign Xxd7x6 = (Lttyx6 & Tttyx6);
assign Tttyx6 = (Butyx6 & Jutyx6);
assign Jutyx6 = (Rutyx6 & Zutyx6);
assign Zutyx6 = (Hvtyx6 & Pvtyx6);
assign Pvtyx6 = (~(Xvtyx6 & Nsoyx6));
assign Xvtyx6 = (Klo7z6[5] & Fwtyx6);
assign Fwtyx6 = (~(Nwtyx6 & Vwtyx6));
assign Vwtyx6 = (Dxtyx6 & Lxtyx6);
assign Lxtyx6 = (Txtyx6 & Bytyx6);
assign Bytyx6 = (~(Hyj7z6[0] & Rbk7z6[2]));
assign Txtyx6 = (~(Hyj7z6[1] & Zlk7z6[2]));
assign Dxtyx6 = (Jytyx6 & Rytyx6);
assign Rytyx6 = (~(Hyj7z6[2] & Hwk7z6[2]));
assign Jytyx6 = (~(Hyj7z6[3] & P6l7z6[2]));
assign Nwtyx6 = (Zytyx6 & Hztyx6);
assign Hztyx6 = (Pztyx6 & Xztyx6);
assign Xztyx6 = (~(Hyj7z6[4] & Xgl7z6[2]));
assign Pztyx6 = (~(Hyj7z6[5] & Frl7z6[2]));
assign Zytyx6 = (F0uyx6 & N0uyx6);
assign N0uyx6 = (~(Hyj7z6[6] & N1m7z6[2]));
assign F0uyx6 = (~(Hyj7z6[7] & Vbm7z6[2]));
assign Hvtyx6 = (V0uyx6 & Votyx6);
assign Votyx6 = (~(Hyj7z6[7] & Dlpyx6));
assign V0uyx6 = (D1uyx6 | L1uyx6);
assign L1uyx6 = (Ti2nz6[2] ? T1uyx6 : Zyoyx6);
assign T1uyx6 = (~(Xzoyx6 & B2uyx6));
assign Zyoyx6 = (!J2uyx6);
assign D1uyx6 = (~(F0pyx6 & R2uyx6));
assign Rutyx6 = (Z2uyx6 & H3uyx6);
assign H3uyx6 = (~(P3uyx6 & Pk1nz6[2]));
assign Z2uyx6 = (~(Bmpyx6 & X3uyx6));
assign X3uyx6 = (~(F4uyx6 & N4uyx6));
assign N4uyx6 = (~(Jw1nz6[2] & Pvpyx6));
assign F4uyx6 = (V4uyx6 & D5uyx6);
assign V4uyx6 = (~(L5uyx6 & Imiiw6));
assign L5uyx6 = (~(Fopyx6 & T5uyx6));
assign Butyx6 = (B6uyx6 & J6uyx6);
assign J6uyx6 = (R6uyx6 & Z6uyx6);
assign Z6uyx6 = (~(Noryx6 & Apget6));
assign Noryx6 = (H7uyx6 & P7uyx6);
assign P7uyx6 = (Dtj7z6[4] & M59iw6);
assign M59iw6 = (!Dtj7z6[3]);
assign H7uyx6 = (Dtj7z6[2] & X7uyx6);
assign R6uyx6 = (F8uyx6 & N8uyx6);
assign N8uyx6 = (~(V8uyx6 & Dlpyx6));
assign Dlpyx6 = (~(D9uyx6 & L9uyx6));
assign L9uyx6 = (~(Q9eiw6 & X7uyx6));
assign D9uyx6 = (~(T9uyx6 & Klo7z6[5]));
assign V8uyx6 = (~(Bauyx6 & Jauyx6));
assign Jauyx6 = (!Hyj7z6[4]);
assign Bauyx6 = (Llpyx6 & Ddsyx6);
assign F8uyx6 = (Rauyx6 | Zauyx6);
assign B6uyx6 = (Hbuyx6 & Pbuyx6);
assign Pbuyx6 = (~(Klo7z6[2] & Xbuyx6));
assign Xbuyx6 = (~(Fcuyx6 & Ncuyx6));
assign Ncuyx6 = (Vcuyx6 & Dduyx6);
assign Dduyx6 = (Lduyx6 & Tduyx6);
assign Tduyx6 = (~(Nqo7z6[0] & M8kiw6));
assign Lduyx6 = (Beuyx6 & Jeuyx6);
assign Jeuyx6 = (~(Reuyx6 & Zeuyx6));
assign Zeuyx6 = (Hfuyx6 & Upeiw6);
assign Reuyx6 = (Pfuyx6 & Z4p7z6[5]);
assign Beuyx6 = (~(R6ryx6 & Z4p7z6[2]));
assign Vcuyx6 = (Xfuyx6 & Fguyx6);
assign Fguyx6 = (~(Fpo7z6[0] & H9kiw6));
assign Xfuyx6 = (~(Ouo7z6[0] & K7kiw6));
assign Fcuyx6 = (Nguyx6 & Vguyx6);
assign Vguyx6 = (Dhuyx6 & Lhuyx6);
assign Lhuyx6 = (~(T2p7z6[2] & U5kiw6));
assign Dhuyx6 = (Thuyx6 & Biuyx6);
assign Biuyx6 = (~(Hxo7z6[0] & W6kiw6));
assign Thuyx6 = (~(Vro7z6[0] & Y7kiw6));
assign Nguyx6 = (Jiuyx6 & Riuyx6);
assign Riuyx6 = (~(W3p7z6[2] & G5kiw6));
assign Jiuyx6 = (~(A0p7z6[0] & I6kiw6));
assign Hbuyx6 = (~(D1pyx6 & Ziuyx6));
assign Ziuyx6 = (~(Hjuyx6 & Pjuyx6));
assign Pjuyx6 = (Xjuyx6 & Fkuyx6);
assign Fkuyx6 = (Nkuyx6 & Vkuyx6);
assign Vkuyx6 = (~(Jdymz6[2] & Sjd8x6));
assign Nkuyx6 = (Dluyx6 & Lluyx6);
assign Lluyx6 = (~(Tluyx6 & Bmuyx6));
assign Tluyx6 = (Gthiw6 & L9pyx6);
assign Dluyx6 = (~(Xbpyx6 & Jmuyx6));
assign Jmuyx6 = (D9pyx6 | Pbpyx6);
assign Xjuyx6 = (Rmuyx6 & Zmuyx6);
assign Zmuyx6 = (~(Tn77v6 & Xm4xx6));
assign Rmuyx6 = (~(Ee77z6 & Vcpyx6));
assign Hjuyx6 = (Hnuyx6 & Pnuyx6);
assign Pnuyx6 = (Xnuyx6 & Fouyx6);
assign Fouyx6 = (~(Biymz6[2] & Ddpyx6));
assign Xnuyx6 = (~(Kmymz6[2] & Lhpyx6));
assign Hnuyx6 = (Nouyx6 & Vouyx6);
assign Vouyx6 = (~(Hcymz6[2] & Hjpyx6));
assign Lttyx6 = (Dpuyx6 & Lpuyx6);
assign Lpuyx6 = (Tpuyx6 & Bquyx6);
assign Bquyx6 = (Jquyx6 & Rquyx6);
assign Rquyx6 = (~(Beryx6 & Klo7z6[0]));
assign Beryx6 = (Zquyx6 & Hruyx6);
assign Hruyx6 = (~(Pruyx6 | Or27v6));
assign Zquyx6 = (~(Xruyx6 | Hnryx6));
assign Jquyx6 = (Fsuyx6 & Nsuyx6);
assign Nsuyx6 = (~(Vsuyx6 & Ngqyx6));
assign Vsuyx6 = (~(Dtuyx6 & Ltuyx6));
assign Ltuyx6 = (Ttuyx6 & Buuyx6);
assign Buuyx6 = (Juuyx6 & Ruuyx6);
assign Ruuyx6 = (Zuuyx6 & Hvuyx6);
assign Hvuyx6 = (~(Voqyx6 & Pvuyx6));
assign Pvuyx6 = (~(Xvuyx6 & Fwuyx6));
assign Fwuyx6 = (~(U3cet6 & Nksyx6));
assign Xvuyx6 = (Nwuyx6 & Vwuyx6);
assign Vwuyx6 = (~(Koaiw6 & Dxuyx6));
assign Nwuyx6 = (Lxuyx6 | Axaiw6);
assign Zuuyx6 = (Txuyx6 & Fkqyx6);
assign Fkqyx6 = (~(Byuyx6 & Koaiw6));
assign Byuyx6 = (Jyuyx6 & Ryuyx6);
assign Ryuyx6 = (~(Zyuyx6 & Hzuyx6));
assign Txuyx6 = (~(Pzuyx6 & Xzuyx6));
assign Pzuyx6 = (Dpadt6 & Vkqyx6);
assign Juuyx6 = (F0vyx6 & N0vyx6);
assign N0vyx6 = (~(Bxi7z6[2] & Dpqyx6));
assign F0vyx6 = (~(A0j7z6[2] & Xrqyx6));
assign Ttuyx6 = (V0vyx6 & D1vyx6);
assign D1vyx6 = (L1vyx6 & T1vyx6);
assign T1vyx6 = (~(H1j7z6[2] & Rqqyx6));
assign L1vyx6 = (~(Ayeet6 & Buqyx6));
assign V0vyx6 = (B2vyx6 & J2vyx6);
assign J2vyx6 = (~(Dxqyx6 & Nob7z6[2]));
assign B2vyx6 = (~(Wui7z6[2] & Lxqyx6));
assign Dtuyx6 = (R2vyx6 & Z2vyx6);
assign Z2vyx6 = (H3vyx6 & P3vyx6);
assign P3vyx6 = (X3vyx6 & F4vyx6);
assign F4vyx6 = (~(Pzqyx6 & G5j7z6[34]));
assign X3vyx6 = (N4vyx6 & V4vyx6);
assign V4vyx6 = (~(Dri7z6[2] & Fwqyx6));
assign N4vyx6 = (~(Bwi7z6[2] & Hzqyx6));
assign H3vyx6 = (D5vyx6 & L5vyx6);
assign L5vyx6 = (~(Jyqyx6 & G5j7z6[2]));
assign D5vyx6 = (~(B2ryx6 & M6j7z6[34]));
assign R2vyx6 = (T5vyx6 & B6vyx6);
assign B6vyx6 = (J6vyx6 & R6vyx6);
assign R6vyx6 = (~(J2ryx6 & M6j7z6[2]));
assign J6vyx6 = (~(D1ryx6 & Ohj7z6[34]));
assign T5vyx6 = (Z6vyx6 & H7vyx6);
assign H7vyx6 = (~(X3ryx6 & Ohj7z6[2]));
assign Z6vyx6 = (~(STCALIB[2] & F4ryx6));
assign Fsuyx6 = (~(Klo7z6[1] & P7vyx6));
assign P7vyx6 = (~(X7vyx6 & F8vyx6));
assign F8vyx6 = (N8vyx6 & V8vyx6);
assign V8vyx6 = (D9vyx6 & L9vyx6);
assign L9vyx6 = (T9vyx6 & Bavyx6);
assign Bavyx6 = (~(Kfq7z6[2] & S7hiw6));
assign T9vyx6 = (Javyx6 & Ravyx6);
assign Javyx6 = (~(Zavyx6 & B2qyx6));
assign Zavyx6 = (~(Zveiw6 | Hbvyx6));
assign D9vyx6 = (Pbvyx6 & Xbvyx6);
assign Xbvyx6 = (~(Hhq7z6[2] & Ydliw6));
assign Pbvyx6 = (Fcvyx6 & Ncvyx6);
assign Ncvyx6 = (~(Tbq7z6[2] & Qsgiw6));
assign Fcvyx6 = (~(Pdq7z6[2] & Oka8x6));
assign N8vyx6 = (Vcvyx6 & Ddvyx6);
assign Ddvyx6 = (Ldvyx6 & Tdvyx6);
assign Tdvyx6 = (~(Y7q7z6[1] & B6qyx6));
assign Ldvyx6 = (Bevyx6 & Jevyx6);
assign Jevyx6 = (~(Cjq7z6[2] & Cza8x6));
assign Bevyx6 = (~(T9tyx6 & Sv77z6));
assign Vcvyx6 = (Revyx6 & Zevyx6);
assign Zevyx6 = (~(D5qyx6 & Bqp7z6[2]));
assign Revyx6 = (~(Z6qyx6 & Gop7z6[2]));
assign X7vyx6 = (Hfvyx6 & Pfvyx6);
assign Pfvyx6 = (Xfvyx6 & Fgvyx6);
assign Fgvyx6 = (Ngvyx6 & Vgvyx6);
assign Vgvyx6 = (~(Ua9ov6 & Sgp7z6[2]));
assign Ngvyx6 = (Dhvyx6 & Lhvyx6);
assign Lhvyx6 = (~(H7qyx6 & Rip7z6[2]));
assign Dhvyx6 = (~(P3a8x6 & Hmp7z6[2]));
assign Xfvyx6 = (Thvyx6 & Bivyx6);
assign Bivyx6 = (~(Fcqyx6 & B2q7z6[2]));
assign Thvyx6 = (Jivyx6 & Rivyx6);
assign Rivyx6 = (~(L9qyx6 & E6p7z6[2]));
assign Jivyx6 = (~(Xbqyx6 & Q8p7z6[2]));
assign Hfvyx6 = (Zivyx6 & Hjvyx6);
assign Hjvyx6 = (Pjvyx6 & Xjvyx6);
assign Xjvyx6 = (~(Q0a8x6 & Hyp7z6[2]));
assign Pjvyx6 = (Fkvyx6 & Nkvyx6);
assign Nkvyx6 = (~(Zaqyx6 & G0q7z6[2]));
assign Fkvyx6 = (~(Nao7x6 & I7p7z6[2]));
assign Zivyx6 = (Vkvyx6 & Dlvyx6);
assign Dlvyx6 = (~(Tdqyx6 & Mkp7z6[2]));
assign Vkvyx6 = (~(U9p7z6[2] & Hfqyx6));
assign Tpuyx6 = (Llvyx6 & Tlvyx6);
assign Tlvyx6 = (~(Scs7z6[2] & Rityx6));
assign Llvyx6 = (Txoyx6 | Bmvyx6);
assign Dpuyx6 = (Jmvyx6 & Rmvyx6);
assign Rmvyx6 = (Zmvyx6 & Hnvyx6);
assign Hnvyx6 = (~(Oo1nz6[2] & Pjtyx6));
assign Zmvyx6 = (~(Au1nz6[2] & Xjtyx6));
assign Jmvyx6 = (Pnvyx6 & Xnvyx6);
assign Xnvyx6 = (~(X66ft6 & Lltyx6));
assign Pnvyx6 = (~(Ies7z6[2] & Tltyx6));
assign Vstyx6 = (~(HRDATAS[2] & Ad47x6));
assign Fstyx6 = (Fovyx6 & Novyx6);
assign Novyx6 = (~(HRDATAD[2] & Mc47x6));
assign Fovyx6 = (~(Zmoyx6 & Eyd7x6));
assign Eyd7x6 = (~(Vovyx6 & Dpvyx6));
assign Dpvyx6 = (~(Xnoyx6 & Eea7z6));
assign Eea7z6 = (~(Lpvyx6 & Tpvyx6));
assign Tpvyx6 = (~(HRDATAD[2] & Qln7z6[0]));
assign Lpvyx6 = (~(HRDATAS[2] & Qln7z6[1]));
assign Vovyx6 = (~(Tim7z6[2] & Tpoyx6));
assign Prtyx6 = (~(Lpryx6 & Vcq7x6));
assign Vpo7v6 = (~(Bqvyx6 & Jqvyx6));
assign Jqvyx6 = (~(Jexmz6[3] & K94iw6));
assign Bqvyx6 = (Rqvyx6 & Zqvyx6);
assign Zqvyx6 = (~(Lloyx6 & Mmlov6));
assign Mmlov6 = (~(Hrvyx6 & Prvyx6));
assign Prvyx6 = (Xrvyx6 & Fsvyx6);
assign Fsvyx6 = (Bqoyx6 | K1e7x6);
assign K1e7x6 = (Nsvyx6 & Vsvyx6);
assign Vsvyx6 = (Dtvyx6 & Ltvyx6);
assign Ltvyx6 = (Ttvyx6 & Buvyx6);
assign Buvyx6 = (Juvyx6 & Ruvyx6);
assign Ruvyx6 = (~(Zuvyx6 & Nsoyx6));
assign Zuvyx6 = (Klo7z6[5] & Hvvyx6);
assign Hvvyx6 = (~(Pvvyx6 & Xvvyx6));
assign Xvvyx6 = (Fwvyx6 & Nwvyx6);
assign Nwvyx6 = (Vwvyx6 & Dxvyx6);
assign Dxvyx6 = (~(Hyj7z6[0] & Rbk7z6[3]));
assign Vwvyx6 = (~(Hyj7z6[1] & Zlk7z6[3]));
assign Fwvyx6 = (Lxvyx6 & Txvyx6);
assign Txvyx6 = (~(Hyj7z6[2] & Hwk7z6[3]));
assign Lxvyx6 = (~(Hyj7z6[3] & P6l7z6[3]));
assign Pvvyx6 = (Byvyx6 & Jyvyx6);
assign Jyvyx6 = (Ryvyx6 & Zyvyx6);
assign Zyvyx6 = (~(Hyj7z6[4] & Xgl7z6[3]));
assign Ryvyx6 = (~(Hyj7z6[5] & Frl7z6[3]));
assign Byvyx6 = (Hzvyx6 & Pzvyx6);
assign Pzvyx6 = (~(Hyj7z6[6] & N1m7z6[3]));
assign Hzvyx6 = (~(Hyj7z6[7] & Vbm7z6[3]));
assign Juvyx6 = (~(Bmpyx6 & Xzvyx6));
assign Xzvyx6 = (~(F0wyx6 & N0wyx6));
assign N0wyx6 = (V0wyx6 & D1wyx6);
assign D1wyx6 = (L1wyx6 & Nopyx6);
assign Nopyx6 = (~(T1wyx6 & J02nz6[5]));
assign T1wyx6 = (B2wyx6 & Imiiw6);
assign V0wyx6 = (J2wyx6 & R2wyx6);
assign R2wyx6 = (~(Nspyx6 & Gie7v6));
assign Nspyx6 = (Z2wyx6 & Puhiw6);
assign J2wyx6 = (~(H3wyx6 & Rgiiw6));
assign H3wyx6 = (Jke7v6 & Imiiw6);
assign F0wyx6 = (P3wyx6 & Nwpyx6);
assign Nwpyx6 = (X3wyx6 & F4wyx6);
assign F4wyx6 = (~(Z2wyx6 & Hrpyx6));
assign X3wyx6 = (D5uyx6 & N4wyx6);
assign D5uyx6 = (~(Pvpyx6 & Imiiw6));
assign Imiiw6 = (!J02nz6[2]);
assign P3wyx6 = (V4wyx6 & D5wyx6);
assign D5wyx6 = (~(Jw1nz6[3] & Pvpyx6));
assign Pvpyx6 = (Pmiiw6 & Jke7v6);
assign Pmiiw6 = (N8syx6 & Basyx6);
assign Basyx6 = (L5wyx6 & T5wyx6);
assign T5wyx6 = (~(J02nz6[3] | J02nz6[6]));
assign L5wyx6 = (B6wyx6 & Thiiw6);
assign N8syx6 = (J02nz6[5] & J02nz6[7]);
assign V4wyx6 = (~(Pk1nz6[3] & Xvpyx6));
assign Ttvyx6 = (J6wyx6 & R6wyx6);
assign R6wyx6 = (Txoyx6 | Z6wyx6);
assign J6wyx6 = (Rauyx6 | Hnryx6);
assign Rauyx6 = (~(H7wyx6 & Klo7z6[0]));
assign H7wyx6 = (~(Xruyx6 | Riryx6));
assign Riryx6 = (!P7wyx6);
assign Dtvyx6 = (X7wyx6 & F8wyx6);
assign F8wyx6 = (~(Klo7z6[1] & N8wyx6));
assign N8wyx6 = (~(V8wyx6 & D9wyx6));
assign D9wyx6 = (L9wyx6 & T9wyx6);
assign T9wyx6 = (Bawyx6 & Jawyx6);
assign Jawyx6 = (Rawyx6 & Zawyx6);
assign Zawyx6 = (~(Pdq7z6[3] & Oka8x6));
assign Rawyx6 = (Hbwyx6 & Pbwyx6);
assign Pbwyx6 = (~(Kfq7z6[3] & S7hiw6));
assign Hbwyx6 = (~(Tbq7z6[3] & Qsgiw6));
assign Bawyx6 = (Xbwyx6 & Fcwyx6);
assign Fcwyx6 = (~(T9tyx6 & Kv77z6));
assign Xbwyx6 = (Ncwyx6 & Vcwyx6);
assign Vcwyx6 = (~(Hhq7z6[3] & Ydliw6));
assign Ncwyx6 = (~(Cjq7z6[3] & Cza8x6));
assign L9wyx6 = (Ddwyx6 & Ldwyx6);
assign Ldwyx6 = (Tdwyx6 & Bewyx6);
assign Bewyx6 = (~(Z6qyx6 & Gop7z6[3]));
assign Tdwyx6 = (Jewyx6 & Rewyx6);
assign Rewyx6 = (~(Y7q7z6[2] & B6qyx6));
assign Jewyx6 = (~(D5qyx6 & Bqp7z6[3]));
assign Ddwyx6 = (Zewyx6 & Hfwyx6);
assign Hfwyx6 = (~(H7qyx6 & Rip7z6[3]));
assign Zewyx6 = (~(P3a8x6 & Hmp7z6[3]));
assign V8wyx6 = (Pfwyx6 & Xfwyx6);
assign Xfwyx6 = (Fgwyx6 & Ngwyx6);
assign Ngwyx6 = (Vgwyx6 & Dhwyx6);
assign Dhwyx6 = (~(Xbqyx6 & Q8p7z6[3]));
assign Vgwyx6 = (Lhwyx6 & Thwyx6);
assign Thwyx6 = (~(Ua9ov6 & Sgp7z6[3]));
assign Lhwyx6 = (~(L9qyx6 & E6p7z6[3]));
assign Fgwyx6 = (Biwyx6 & Jiwyx6);
assign Jiwyx6 = (~(Fcqyx6 & B2q7z6[3]));
assign Biwyx6 = (~(Zaqyx6 & G0q7z6[3]));
assign Pfwyx6 = (Riwyx6 & Ziwyx6);
assign Ziwyx6 = (Hjwyx6 & Pjwyx6);
assign Pjwyx6 = (~(Tdqyx6 & Mkp7z6[3]));
assign Hjwyx6 = (Xjwyx6 & Fkwyx6);
assign Fkwyx6 = (~(Nao7x6 & I7p7z6[3]));
assign Xjwyx6 = (~(Q0a8x6 & Hyp7z6[3]));
assign Riwyx6 = (Reqyx6 & Nkwyx6);
assign Nkwyx6 = (~(U9p7z6[3] & Hfqyx6));
assign Reqyx6 = (Fgtyx6 & Vkwyx6);
assign Vkwyx6 = (~(B2qyx6 & R6tyx6));
assign X7wyx6 = (Dlwyx6 & Llwyx6);
assign Llwyx6 = (~(Scs7z6[3] & Rityx6));
assign Rityx6 = (Klo7z6[0] & Zmryx6);
assign Dlwyx6 = (~(Tlwyx6 & Ngqyx6));
assign Tlwyx6 = (~(Bmwyx6 & Jmwyx6));
assign Jmwyx6 = (Rmwyx6 & Zmwyx6);
assign Zmwyx6 = (Hnwyx6 & Pnwyx6);
assign Pnwyx6 = (Xnwyx6 & Fowyx6);
assign Fowyx6 = (~(Nowyx6 & Vveet6));
assign Nowyx6 = (Buqyx6 & Cwadt6);
assign Xnwyx6 = (Vowyx6 & Pjqyx6);
assign Pjqyx6 = (~(Dpwyx6 & Jyuyx6));
assign Vowyx6 = (~(Lpwyx6 & Koaiw6));
assign Lpwyx6 = (Voqyx6 & Jyuyx6);
assign Hnwyx6 = (Tpwyx6 & Bqwyx6);
assign Bqwyx6 = (~(Bxi7z6[3] & Dpqyx6));
assign Tpwyx6 = (~(Dradt6 & Hnqyx6));
assign Rmwyx6 = (Jqwyx6 & Rqwyx6);
assign Rqwyx6 = (Zqwyx6 & Hrwyx6);
assign Hrwyx6 = (~(H1j7z6[3] & Rqqyx6));
assign Zqwyx6 = (Prwyx6 & Xrwyx6);
assign Xrwyx6 = (~(Prqyx6 & Z3j7z6[3]));
assign Prwyx6 = (~(A0j7z6[3] & Xrqyx6));
assign Jqwyx6 = (Fswyx6 & Nswyx6);
assign Nswyx6 = (~(Bzi7z6[3] & Vsqyx6));
assign Fswyx6 = (~(Dxqyx6 & Nob7z6[3]));
assign Bmwyx6 = (Vswyx6 & Dtwyx6);
assign Dtwyx6 = (Ltwyx6 & Ttwyx6);
assign Ttwyx6 = (Buwyx6 & Juwyx6);
assign Juwyx6 = (~(Bwi7z6[3] & Hzqyx6));
assign Buwyx6 = (Ruwyx6 & Zuwyx6);
assign Zuwyx6 = (~(Wui7z6[3] & Lxqyx6));
assign Ruwyx6 = (~(Dri7z6[3] & Fwqyx6));
assign Ltwyx6 = (Hvwyx6 & Pvwyx6);
assign Pvwyx6 = (~(Pzqyx6 & G5j7z6[35]));
assign Hvwyx6 = (~(Jyqyx6 & G5j7z6[3]));
assign Vswyx6 = (Xvwyx6 & Fwwyx6);
assign Fwwyx6 = (Nwwyx6 & Vwwyx6);
assign Vwwyx6 = (~(D1ryx6 & Ohj7z6[35]));
assign Nwwyx6 = (Dxwyx6 & Lxwyx6);
assign Lxwyx6 = (~(B2ryx6 & M6j7z6[35]));
assign Dxwyx6 = (~(J2ryx6 & M6j7z6[3]));
assign Xvwyx6 = (Txwyx6 & Bywyx6);
assign Bywyx6 = (~(X3ryx6 & Ohj7z6[3]));
assign Txwyx6 = (~(STCALIB[3] & F4ryx6));
assign Nsvyx6 = (Jywyx6 & Rywyx6);
assign Rywyx6 = (Zywyx6 & Hzwyx6);
assign Hzwyx6 = (Pzwyx6 & Xzwyx6);
assign Xzwyx6 = (~(D1pyx6 & F0xyx6));
assign F0xyx6 = (~(N0xyx6 & V0xyx6));
assign V0xyx6 = (D1xyx6 & L1xyx6);
assign L1xyx6 = (T1xyx6 & B2xyx6);
assign B2xyx6 = (~(Jdymz6[3] & Sjd8x6));
assign Sjd8x6 = (Zshiw6 & J2xyx6);
assign T1xyx6 = (R2xyx6 & L5pyx6);
assign D1xyx6 = (Z2xyx6 & H3xyx6);
assign H3xyx6 = (~(Gm77v6 & Xm4xx6));
assign Xm4xx6 = (Gthiw6 & P3xyx6);
assign N0xyx6 = (X3xyx6 & F4xyx6);
assign F4xyx6 = (N4xyx6 & V4xyx6);
assign V4xyx6 = (~(Kmymz6[3] & Lhpyx6));
assign N4xyx6 = (D5xyx6 & L5xyx6);
assign L5xyx6 = (~(Cf77z6 & Vcpyx6));
assign D5xyx6 = (~(Biymz6[3] & Ddpyx6));
assign X3xyx6 = (Nouyx6 & T5xyx6);
assign T5xyx6 = (~(Hcymz6[3] & Hjpyx6));
assign Nouyx6 = (B6xyx6 & J6xyx6);
assign J6xyx6 = (R6xyx6 & Z6xyx6);
assign Z6xyx6 = (~(Lzqnv6 & Thpyx6));
assign R6xyx6 = (~(Zcsnv6 & Ngpyx6));
assign B6xyx6 = (Ripyx6 & H7xyx6);
assign H7xyx6 = (~(Eg4xx6 & Hfpyx6));
assign Ripyx6 = (Qid8x6 & P7xyx6);
assign P7xyx6 = (~(Gthiw6 & Xbpyx6));
assign Qid8x6 = (!Ljd8x6);
assign Ljd8x6 = (D9pyx6 & Zshiw6);
assign Pzwyx6 = (~(Klo7z6[2] & X7xyx6));
assign X7xyx6 = (~(F8xyx6 & N8xyx6));
assign N8xyx6 = (V8xyx6 & D9xyx6);
assign D9xyx6 = (L9xyx6 & T9xyx6);
assign T9xyx6 = (~(Nqo7z6[1] & M8kiw6));
assign L9xyx6 = (Baxyx6 & Jaxyx6);
assign Baxyx6 = (~(R6ryx6 & Pfuyx6));
assign V8xyx6 = (Raxyx6 & Zaxyx6);
assign Zaxyx6 = (~(Fpo7z6[1] & H9kiw6));
assign Raxyx6 = (~(Ouo7z6[1] & K7kiw6));
assign F8xyx6 = (Hbxyx6 & Pbxyx6);
assign Pbxyx6 = (Xbxyx6 & Fcxyx6);
assign Fcxyx6 = (~(T2p7z6[3] & U5kiw6));
assign Xbxyx6 = (Ncxyx6 & Vcxyx6);
assign Vcxyx6 = (~(Hxo7z6[1] & W6kiw6));
assign Ncxyx6 = (~(Vro7z6[1] & Y7kiw6));
assign Hbxyx6 = (Ddxyx6 & Ldxyx6);
assign Ldxyx6 = (~(W3p7z6[3] & G5kiw6));
assign Ddxyx6 = (~(A0p7z6[1] & I6kiw6));
assign Zywyx6 = (Tdxyx6 & Bexyx6);
assign Bexyx6 = (~(Oo1nz6[3] & Pjtyx6));
assign Tdxyx6 = (~(Au1nz6[3] & Xjtyx6));
assign Jywyx6 = (Jexyx6 & Bmtyx6);
assign Bmtyx6 = (Rexyx6 & Zexyx6);
assign Zexyx6 = (Hfxyx6 | Txoyx6);
assign Txoyx6 = (~(Pfxyx6 & F0pyx6));
assign Hfxyx6 = (R2uyx6 | Ti2nz6[2]);
assign Rexyx6 = (~(Xfxyx6 & Klo7z6[0]));
assign Jexyx6 = (Fgxyx6 & Ngxyx6);
assign Ngxyx6 = (~(Lltyx6 & D86ft6));
assign Fgxyx6 = (~(Ies7z6[3] & Tltyx6));
assign Xrvyx6 = (~(Zmoyx6 & R1e7x6));
assign R1e7x6 = (~(Vgxyx6 & Dhxyx6));
assign Dhxyx6 = (~(Xnoyx6 & Wda7z6));
assign Wda7z6 = (~(Lhxyx6 & Thxyx6));
assign Thxyx6 = (~(HRDATAD[3] & Qln7z6[0]));
assign Lhxyx6 = (~(HRDATAS[3] & Qln7z6[1]));
assign Vgxyx6 = (~(Tim7z6[3] & Tpoyx6));
assign Hrvyx6 = (Bixyx6 & Jixyx6);
assign Jixyx6 = (~(HRDATAS[3] & Ad47x6));
assign Bixyx6 = (~(HRDATAD[3] & Mc47x6));
assign Rqvyx6 = (~(Lpryx6 & Fiq7x6));
assign Opo7v6 = (~(Rixyx6 & Zixyx6));
assign Zixyx6 = (~(Jexmz6[4] & K94iw6));
assign Rixyx6 = (Hjxyx6 & Pjxyx6);
assign Pjxyx6 = (~(Lloyx6 & Cb77x6));
assign Cb77x6 = (~(Xjxyx6 & Fkxyx6));
assign Fkxyx6 = (Nkxyx6 & Vkxyx6);
assign Vkxyx6 = (Bqoyx6 | X4e7x6);
assign X4e7x6 = (Dlxyx6 & Llxyx6);
assign Llxyx6 = (Tlxyx6 & Bmxyx6);
assign Bmxyx6 = (Jmxyx6 & Rmxyx6);
assign Rmxyx6 = (Zmxyx6 & Hnxyx6);
assign Hnxyx6 = (~(Pnxyx6 & Nsoyx6));
assign Pnxyx6 = (Klo7z6[5] & Xnxyx6);
assign Xnxyx6 = (~(Foxyx6 & Noxyx6));
assign Noxyx6 = (Voxyx6 & Dpxyx6);
assign Dpxyx6 = (Lpxyx6 & Tpxyx6);
assign Tpxyx6 = (~(Hyj7z6[0] & Rbk7z6[4]));
assign Lpxyx6 = (~(Hyj7z6[1] & Zlk7z6[4]));
assign Voxyx6 = (Bqxyx6 & Jqxyx6);
assign Jqxyx6 = (~(Hyj7z6[2] & Hwk7z6[4]));
assign Bqxyx6 = (~(Hyj7z6[3] & P6l7z6[4]));
assign Foxyx6 = (Rqxyx6 & Zqxyx6);
assign Zqxyx6 = (Hrxyx6 & Prxyx6);
assign Prxyx6 = (~(Hyj7z6[4] & Xgl7z6[4]));
assign Hrxyx6 = (~(Hyj7z6[5] & Frl7z6[4]));
assign Rqxyx6 = (Xrxyx6 & Fsxyx6);
assign Fsxyx6 = (~(Hyj7z6[6] & N1m7z6[4]));
assign Xrxyx6 = (~(Hyj7z6[7] & Vbm7z6[4]));
assign Zmxyx6 = (~(Nsxyx6 & J2uyx6));
assign Nsxyx6 = (F0pyx6 & R2uyx6);
assign Jmxyx6 = (Vsxyx6 & Dtxyx6);
assign Dtxyx6 = (~(Bmpyx6 & Ltxyx6));
assign Ltxyx6 = (~(Ttxyx6 & Buxyx6));
assign Buxyx6 = (Juxyx6 & N4wyx6);
assign Juxyx6 = (Ruxyx6 & Vopyx6);
assign Vopyx6 = (~(Zuxyx6 & Hvxyx6));
assign Hvxyx6 = (Pvxyx6 & B6wyx6);
assign Pvxyx6 = (Xvxyx6 & L9syx6);
assign Zuxyx6 = (J02nz6[3] & J02nz6[2]);
assign Ttxyx6 = (Fwxyx6 & Nwxyx6);
assign Nwxyx6 = (~(Pk1nz6[4] & Xvpyx6));
assign Fwxyx6 = (Vwxyx6 & L1wyx6);
assign Vsxyx6 = (~(D1pyx6 & Dxxyx6));
assign Dxxyx6 = (~(Lxxyx6 & Txxyx6));
assign Txxyx6 = (Byxyx6 & Jyxyx6);
assign Jyxyx6 = (Ryxyx6 & Zyxyx6);
assign Zyxyx6 = (~(Hzxyx6 & Eg4xx6));
assign Eg4xx6 = (Pzxyx6 & Ojymz6[3]);
assign Pzxyx6 = (Ojymz6[1] & Ojymz6[0]);
assign Hzxyx6 = (Hfpyx6 & Jf4xx6);
assign Jf4xx6 = (!Ojymz6[2]);
assign Ryxyx6 = (Xzxyx6 & F0yyx6);
assign F0yyx6 = (~(N0yyx6 & Lzqnv6));
assign Lzqnv6 = (V0yyx6 & Unymz6[3]);
assign V0yyx6 = (Unymz6[1] & Unymz6[0]);
assign N0yyx6 = (Thpyx6 & Qyqnv6);
assign Qyqnv6 = (!Unymz6[2]);
assign Xzxyx6 = (~(D1yyx6 & Zcsnv6));
assign Zcsnv6 = (L1yyx6 & Sgymz6[3]);
assign L1yyx6 = (Sgymz6[1] & Sgymz6[0]);
assign D1yyx6 = (Ngpyx6 & Xbsnv6);
assign Xbsnv6 = (!Sgymz6[2]);
assign Byxyx6 = (T1yyx6 & B2yyx6);
assign B2yyx6 = (~(J2yyx6 & V4pyx6));
assign J2yyx6 = (D9pyx6 & F02nv6);
assign T1yyx6 = (~(Kf77z6 & Vcpyx6));
assign Lxxyx6 = (R2yyx6 & Z2yyx6);
assign Z2yyx6 = (H3yyx6 & P3yyx6);
assign P3yyx6 = (~(Hcymz6[4] & Hjpyx6));
assign H3yyx6 = (X3yyx6 & F4yyx6);
assign F4yyx6 = (~(Biymz6[4] & Ddpyx6));
assign X3yyx6 = (~(Feymz6[0] & Fgpyx6));
assign R2yyx6 = (N4yyx6 & Xjpyx6);
assign Xjpyx6 = (V4yyx6 & D5yyx6);
assign D5yyx6 = (~(L5yyx6 & T5yyx6));
assign T5yyx6 = (Bmuyx6 & B6yyx6);
assign B6yyx6 = (J6yyx6 & R6pyx6);
assign Bmuyx6 = (Xfymz6[7] & Xfymz6[6]);
assign L5yyx6 = (R6yyx6 & Xfymz6[3]);
assign R6yyx6 = (Xfymz6[2] & L9pyx6);
assign V4yyx6 = (R2xyx6 & Z6yyx6);
assign Tlxyx6 = (H7yyx6 & P7yyx6);
assign P7yyx6 = (~(Klo7z6[1] & X7yyx6));
assign X7yyx6 = (~(F8yyx6 & N8yyx6));
assign N8yyx6 = (V8yyx6 & D9yyx6);
assign D9yyx6 = (L9yyx6 & T9yyx6);
assign T9yyx6 = (Bayyx6 & T1qyx6);
assign Bayyx6 = (~(Kfq7z6[4] & S7hiw6));
assign L9yyx6 = (Jayyx6 & Rayyx6);
assign Rayyx6 = (~(Tbq7z6[4] & Qsgiw6));
assign Jayyx6 = (~(Pdq7z6[4] & Oka8x6));
assign V8yyx6 = (Zayyx6 & Hbyyx6);
assign Hbyyx6 = (Pbyyx6 & Xbyyx6);
assign Xbyyx6 = (~(Hhq7z6[4] & Ydliw6));
assign Pbyyx6 = (~(Cjq7z6[4] & Cza8x6));
assign Zayyx6 = (Fcyyx6 & Ncyyx6);
assign Ncyyx6 = (~(Vcyyx6 & R6tyx6));
assign Fcyyx6 = (~(T9tyx6 & Cv77z6));
assign F8yyx6 = (Ddyyx6 & Ldyyx6);
assign Ldyyx6 = (Tdyyx6 & Beyyx6);
assign Beyyx6 = (Jeyyx6 & Reyyx6);
assign Reyyx6 = (~(Y7q7z6[3] & B6qyx6));
assign Jeyyx6 = (~(D5qyx6 & Bqp7z6[4]));
assign Tdyyx6 = (Zeyyx6 & Hfyyx6);
assign Hfyyx6 = (~(L9qyx6 & E6p7z6[4]));
assign Zeyyx6 = (~(Fcqyx6 & B2q7z6[4]));
assign Ddyyx6 = (Pfyyx6 & Fgtyx6);
assign Pfyyx6 = (Xfyyx6 & Fgyyx6);
assign Fgyyx6 = (~(Tdqyx6 & Mkp7z6[4]));
assign Xfyyx6 = (~(U9p7z6[4] & Hfqyx6));
assign H7yyx6 = (Ngyyx6 & Vgyyx6);
assign Vgyyx6 = (~(Klo7z6[2] & Dhyyx6));
assign Dhyyx6 = (~(Lhyyx6 & Thyyx6));
assign Thyyx6 = (Biyyx6 & Jiyyx6);
assign Jiyyx6 = (Riyyx6 & Ziyyx6);
assign Ziyyx6 = (~(Ouo7z6[2] & K7kiw6));
assign Riyyx6 = (Hjyyx6 & Pjyyx6);
assign Pjyyx6 = (~(Nqo7z6[2] & M8kiw6));
assign Hjyyx6 = (~(Fpo7z6[2] & H9kiw6));
assign Biyyx6 = (Xjyyx6 & Fkyyx6);
assign Fkyyx6 = (~(Hxo7z6[2] & W6kiw6));
assign Xjyyx6 = (~(Vro7z6[2] & Y7kiw6));
assign Lhyyx6 = (Nkyyx6 & Vkyyx6);
assign Vkyyx6 = (Dlyyx6 & Llyyx6);
assign Llyyx6 = (~(T2p7z6[4] & U5kiw6));
assign Dlyyx6 = (~(W3p7z6[4] & G5kiw6));
assign Nkyyx6 = (Tlyyx6 & Bmyyx6);
assign Bmyyx6 = (~(A0p7z6[2] & I6kiw6));
assign Ngyyx6 = (~(Jmyyx6 & Ngqyx6));
assign Jmyyx6 = (~(Rmyyx6 & Zmyyx6));
assign Zmyyx6 = (Hnyyx6 & Pnyyx6);
assign Pnyyx6 = (Xnyyx6 & Foyyx6);
assign Foyyx6 = (Noyyx6 & Voyyx6);
assign Voyyx6 = (~(Dpyyx6 & Lpyyx6));
assign Dpyyx6 = (Jyuyx6 & Tpyyx6);
assign Noyyx6 = (Hjqyx6 & Bqyyx6);
assign Xnyyx6 = (Jqyyx6 & Rqyyx6);
assign Rqyyx6 = (~(Esadt6 & Hnqyx6));
assign Jqyyx6 = (Zqyyx6 & Hryyx6);
assign Hryyx6 = (~(Pryyx6 & L2cet6));
assign Pryyx6 = (Nksyx6 & Voqyx6);
assign Zqyyx6 = (~(Bxi7z6[4] & Dpqyx6));
assign Dpqyx6 = (Xryyx6 & Voqyx6);
assign Hnyyx6 = (Fsyyx6 & Nsyyx6);
assign Nsyyx6 = (Vsyyx6 & Dtyyx6);
assign Dtyyx6 = (~(Brdet6 & Ttqyx6));
assign Vsyyx6 = (Ltyyx6 & Ttyyx6);
assign Ttyyx6 = (~(A0j7z6[4] & Xrqyx6));
assign Ltyyx6 = (~(H1j7z6[4] & Rqqyx6));
assign Fsyyx6 = (Buyyx6 & Juyyx6);
assign Juyyx6 = (~(Bzi7z6[4] & Vsqyx6));
assign Buyyx6 = (~(Dxqyx6 & Nob7z6[4]));
assign Rmyyx6 = (Ruyyx6 & Zuyyx6);
assign Zuyyx6 = (Hvyyx6 & Pvyyx6);
assign Pvyyx6 = (Xvyyx6 & Fwyyx6);
assign Fwyyx6 = (~(Bwi7z6[4] & Hzqyx6));
assign Xvyyx6 = (Nwyyx6 & Vwyyx6);
assign Vwyyx6 = (~(Wui7z6[4] & Lxqyx6));
assign Nwyyx6 = (~(Dri7z6[4] & Fwqyx6));
assign Hvyyx6 = (Dxyyx6 & Lxyyx6);
assign Lxyyx6 = (~(B2ryx6 & M6j7z6[36]));
assign Dxyyx6 = (Txyyx6 & Byyyx6);
assign Byyyx6 = (~(Pzqyx6 & G5j7z6[36]));
assign Txyyx6 = (~(Jyqyx6 & G5j7z6[4]));
assign Ruyyx6 = (Jyyyx6 & Ryyyx6);
assign Ryyyx6 = (Zyyyx6 & Hzyyx6);
assign Hzyyx6 = (~(X3ryx6 & Ohj7z6[4]));
assign Zyyyx6 = (Pzyyx6 & Xzyyx6);
assign Xzyyx6 = (~(J2ryx6 & M6j7z6[4]));
assign Pzyyx6 = (~(D1ryx6 & Ohj7z6[36]));
assign Jyyyx6 = (F0zyx6 & N0zyx6);
assign N0zyx6 = (~(STCALIB[4] & F4ryx6));
assign Dlxyx6 = (V0zyx6 & D1zyx6);
assign D1zyx6 = (L1zyx6 & T1zyx6);
assign T1zyx6 = (~(Au1nz6[4] & Xjtyx6));
assign L1zyx6 = (B2zyx6 & J2zyx6);
assign J2zyx6 = (R2zyx6 | Ap27v6);
assign B2zyx6 = (~(Oo1nz6[4] & Pjtyx6));
assign V0zyx6 = (Z2zyx6 & H3zyx6);
assign Z2zyx6 = (P3zyx6 & X3zyx6);
assign X3zyx6 = (~(Og6ft6 & Lltyx6));
assign P3zyx6 = (~(Ies7z6[4] & Tltyx6));
assign Nkxyx6 = (~(Zmoyx6 & E5e7x6));
assign E5e7x6 = (~(F4zyx6 & N4zyx6));
assign N4zyx6 = (~(Qco7v6 & Xnoyx6));
assign F4zyx6 = (~(Tim7z6[4] & Tpoyx6));
assign Xjxyx6 = (V4zyx6 & D5zyx6);
assign D5zyx6 = (~(HRDATAS[4] & Ad47x6));
assign V4zyx6 = (~(HRDATAD[4] & Mc47x6));
assign Hjxyx6 = (~(Lpryx6 & Pnq7x6));
assign Hpo7v6 = (~(L5zyx6 & T5zyx6));
assign T5zyx6 = (~(Jexmz6[5] & K94iw6));
assign L5zyx6 = (B6zyx6 & J6zyx6);
assign J6zyx6 = (~(Lloyx6 & C477x6));
assign C477x6 = (~(R6zyx6 & Z6zyx6));
assign Z6zyx6 = (H7zyx6 & P7zyx6);
assign P7zyx6 = (Bqoyx6 | K8e7x6);
assign K8e7x6 = (X7zyx6 & F8zyx6);
assign F8zyx6 = (N8zyx6 & V8zyx6);
assign V8zyx6 = (D9zyx6 & L9zyx6);
assign L9zyx6 = (T9zyx6 & R2zyx6);
assign T9zyx6 = (~(P3uyx6 & Pk1nz6[5]));
assign D9zyx6 = (Bazyx6 & Jazyx6);
assign Jazyx6 = (~(Bmpyx6 & Razyx6));
assign Razyx6 = (~(Vwpyx6 & N4wyx6));
assign N4wyx6 = (~(Zazyx6 & Hrpyx6));
assign Zazyx6 = (Tppyx6 & J02nz6[8]);
assign Vwpyx6 = (Hbzyx6 & V4syx6);
assign V4syx6 = (~(Pbzyx6 & Hrpyx6));
assign Bmpyx6 = (Kniiw6 & Klo7z6[3]);
assign Bazyx6 = (~(Xbzyx6 & Fczyx6));
assign Fczyx6 = (~(Nczyx6 & Vczyx6));
assign Vczyx6 = (Ddzyx6 & Ldzyx6);
assign Ldzyx6 = (Tdzyx6 & Bezyx6);
assign Bezyx6 = (~(Hyj7z6[0] & Rbk7z6[5]));
assign Tdzyx6 = (~(Hyj7z6[1] & Zlk7z6[5]));
assign Ddzyx6 = (Jezyx6 & Rezyx6);
assign Rezyx6 = (~(Hyj7z6[2] & Hwk7z6[5]));
assign Jezyx6 = (~(Hyj7z6[3] & P6l7z6[5]));
assign Nczyx6 = (Zezyx6 & Hfzyx6);
assign Hfzyx6 = (Pfzyx6 & Xfzyx6);
assign Xfzyx6 = (~(Hyj7z6[4] & Xgl7z6[5]));
assign Pfzyx6 = (~(Hyj7z6[5] & Frl7z6[5]));
assign Zezyx6 = (Fgzyx6 & Ngzyx6);
assign Ngzyx6 = (~(Hyj7z6[6] & N1m7z6[5]));
assign Fgzyx6 = (~(Hyj7z6[7] & Vbm7z6[5]));
assign N8zyx6 = (Vgzyx6 & Dhzyx6);
assign Dhzyx6 = (~(D1pyx6 & Lhzyx6));
assign Lhzyx6 = (~(Thzyx6 & Bizyx6));
assign Bizyx6 = (Jizyx6 & Rizyx6);
assign Rizyx6 = (Zizyx6 & Hjzyx6);
assign Hjzyx6 = (~(Sf77z6 & Vcpyx6));
assign Zizyx6 = (Pjzyx6 & R2xyx6);
assign R2xyx6 = (~(Ied8x6 & Xbpyx6));
assign Pjzyx6 = (~(D9pyx6 & Xbpyx6));
assign Jizyx6 = (Xjzyx6 & Fkzyx6);
assign Fkzyx6 = (~(Biymz6[5] & Ddpyx6));
assign Xjzyx6 = (~(Feymz6[1] & Fgpyx6));
assign Thzyx6 = (Nkzyx6 & Vkzyx6);
assign Vkzyx6 = (Dlzyx6 & Llzyx6);
assign Llzyx6 = (~(Sgymz6[2] & Ngpyx6));
assign Dlzyx6 = (~(Ojymz6[2] & Hfpyx6));
assign Nkzyx6 = (Pjpyx6 & Tlzyx6);
assign Tlzyx6 = (~(Unymz6[2] & Thpyx6));
assign Vgzyx6 = (Bmzyx6 & Jmzyx6);
assign Jmzyx6 = (~(Rmzyx6 & Zmzyx6));
assign Zmzyx6 = (~(Hnzyx6 & Pnzyx6));
assign Pnzyx6 = (Xnzyx6 & Fozyx6);
assign Fozyx6 = (Nozyx6 & Vozyx6);
assign Vozyx6 = (~(Hyj7z6[0] & Dfk7z6[5]));
assign Nozyx6 = (~(Hyj7z6[1] & Lpk7z6[5]));
assign Xnzyx6 = (Dpzyx6 & Lpzyx6);
assign Lpzyx6 = (~(Hyj7z6[2] & Tzk7z6[5]));
assign Dpzyx6 = (~(Hyj7z6[3] & Bal7z6[5]));
assign Hnzyx6 = (Tpzyx6 & Bqzyx6);
assign Bqzyx6 = (Jqzyx6 & Rqzyx6);
assign Rqzyx6 = (~(Hyj7z6[4] & Jkl7z6[5]));
assign Jqzyx6 = (~(Hyj7z6[5] & Rul7z6[5]));
assign Tpzyx6 = (Zqzyx6 & Hrzyx6);
assign Hrzyx6 = (~(Hyj7z6[6] & Z4m7z6[5]));
assign Zqzyx6 = (~(Hyj7z6[7] & Hfm7z6[5]));
assign Bmzyx6 = (~(Klo7z6[2] & Przyx6));
assign Przyx6 = (~(Xrzyx6 & Fszyx6));
assign Fszyx6 = (Nszyx6 & Vszyx6);
assign Vszyx6 = (Dtzyx6 & Ltzyx6);
assign Ltzyx6 = (~(Fpo7z6[3] & H9kiw6));
assign Dtzyx6 = (Ttzyx6 & Jaxyx6);
assign Jaxyx6 = (~(Buzyx6 & R6ryx6));
assign R6ryx6 = (Juzyx6 & Hfuyx6);
assign Juzyx6 = (!Ruzyx6);
assign Buzyx6 = (Z4p7z6[1] & R2syx6);
assign Ttzyx6 = (~(Nqo7z6[3] & M8kiw6));
assign Nszyx6 = (Zuzyx6 & Hvzyx6);
assign Hvzyx6 = (~(Hxo7z6[3] & W6kiw6));
assign Zuzyx6 = (Pvzyx6 & Xvzyx6);
assign Xvzyx6 = (~(Vitet6 & S4kiw6));
assign Pvzyx6 = (~(Ouo7z6[3] & K7kiw6));
assign Xrzyx6 = (Fwzyx6 & Nwzyx6);
assign Nwzyx6 = (Vwzyx6 & Dxzyx6);
assign Dxzyx6 = (~(W3p7z6[5] & G5kiw6));
assign Vwzyx6 = (Lxzyx6 & Txzyx6);
assign Txzyx6 = (~(Vro7z6[3] & Y7kiw6));
assign Lxzyx6 = (~(T2p7z6[5] & U5kiw6));
assign Fwzyx6 = (Byzyx6 & Jyzyx6);
assign Byzyx6 = (Tlyyx6 & Ryzyx6);
assign Ryzyx6 = (~(A0p7z6[3] & I6kiw6));
assign X7zyx6 = (Zyzyx6 & Hzzyx6);
assign Hzzyx6 = (Pzzyx6 & Xzzyx6);
assign Xzzyx6 = (~(Oo1nz6[5] & Pjtyx6));
assign Pzzyx6 = (F00zx6 & N00zx6);
assign N00zx6 = (~(V00zx6 & Ngqyx6));
assign V00zx6 = (~(D10zx6 & L10zx6));
assign L10zx6 = (T10zx6 & B20zx6);
assign B20zx6 = (J20zx6 & R20zx6);
assign R20zx6 = (Z20zx6 & H30zx6);
assign H30zx6 = (P30zx6 & X30zx6);
assign X30zx6 = (~(H1j7z6[5] & Rqqyx6));
assign P30zx6 = (F40zx6 & N40zx6);
assign N40zx6 = (~(V40zx6 & Ffj7z6[0]));
assign F40zx6 = (~(A0j7z6[5] & Xrqyx6));
assign Z20zx6 = (D50zx6 & L50zx6);
assign L50zx6 = (~(Zsdet6 & Ttqyx6));
assign D50zx6 = (~(Qteet6 & Buqyx6));
assign J20zx6 = (T50zx6 & B60zx6);
assign B60zx6 = (J60zx6 & 1'b1);
assign J60zx6 = (~(Dxqyx6 & Nob7z6[5]));
assign T50zx6 = (R60zx6 & Z60zx6);
assign Z60zx6 = (~(Wui7z6[5] & Lxqyx6));
assign R60zx6 = (~(Dri7z6[5] & Fwqyx6));
assign T10zx6 = (H70zx6 & P70zx6);
assign P70zx6 = (X70zx6 & F80zx6);
assign F80zx6 = (N80zx6 & V80zx6);
assign V80zx6 = (~(D90zx6 & Lgj7z6[180]));
assign N80zx6 = (L90zx6 & T90zx6);
assign T90zx6 = (~(Bwi7z6[5] & Hzqyx6));
assign L90zx6 = (~(Ba0zx6 & Nbj7z6[0]));
assign X70zx6 = (Ja0zx6 & Ra0zx6);
assign Ra0zx6 = (~(Za0zx6 & Lgj7z6[168]));
assign Ja0zx6 = (~(Hb0zx6 & Lgj7z6[156]));
assign H70zx6 = (Pb0zx6 & Xb0zx6);
assign Xb0zx6 = (Fc0zx6 & Nc0zx6);
assign Nc0zx6 = (~(Vc0zx6 & Lgj7z6[144]));
assign Fc0zx6 = (~(Dd0zx6 & Lgj7z6[132]));
assign Pb0zx6 = (Ld0zx6 & Td0zx6);
assign Td0zx6 = (~(Be0zx6 & Lgj7z6[120]));
assign Ld0zx6 = (~(Je0zx6 & Lgj7z6[108]));
assign D10zx6 = (Re0zx6 & Ze0zx6);
assign Ze0zx6 = (Hf0zx6 & Pf0zx6);
assign Pf0zx6 = (Xf0zx6 & Fg0zx6);
assign Fg0zx6 = (Ng0zx6 & Vg0zx6);
assign Vg0zx6 = (~(Dh0zx6 & Lgj7z6[72]));
assign Ng0zx6 = (Lh0zx6 & Th0zx6);
assign Th0zx6 = (~(Bi0zx6 & Lgj7z6[96]));
assign Lh0zx6 = (~(Ji0zx6 & Lgj7z6[84]));
assign Xf0zx6 = (Ri0zx6 & Zi0zx6);
assign Zi0zx6 = (~(Hj0zx6 & Lgj7z6[60]));
assign Ri0zx6 = (~(Pj0zx6 & Lgj7z6[48]));
assign Hf0zx6 = (Xj0zx6 & Fk0zx6);
assign Fk0zx6 = (Nk0zx6 & Vk0zx6);
assign Vk0zx6 = (~(Dl0zx6 & Lgj7z6[36]));
assign Nk0zx6 = (~(Ll0zx6 & Lgj7z6[24]));
assign Xj0zx6 = (Tl0zx6 & Bm0zx6);
assign Bm0zx6 = (~(Jm0zx6 & Lgj7z6[12]));
assign Tl0zx6 = (~(Rm0zx6 & Lgj7z6[0]));
assign Re0zx6 = (Zm0zx6 & Hn0zx6);
assign Hn0zx6 = (Pn0zx6 & Xn0zx6);
assign Xn0zx6 = (Fo0zx6 & No0zx6);
assign No0zx6 = (~(B2ryx6 & M6j7z6[37]));
assign Fo0zx6 = (Vo0zx6 & Dp0zx6);
assign Dp0zx6 = (~(Pzqyx6 & G5j7z6[37]));
assign Vo0zx6 = (~(Jyqyx6 & G5j7z6[5]));
assign Pn0zx6 = (Lp0zx6 & Tp0zx6);
assign Tp0zx6 = (~(J2ryx6 & M6j7z6[5]));
assign Lp0zx6 = (~(D1ryx6 & Ohj7z6[37]));
assign Zm0zx6 = (Bq0zx6 & Jq0zx6);
assign Jq0zx6 = (Rq0zx6 & Zq0zx6);
assign Zq0zx6 = (~(X3ryx6 & Ohj7z6[5]));
assign Rq0zx6 = (~(STCALIB[5] & F4ryx6));
assign Bq0zx6 = (F0zyx6 & Hr0zx6);
assign F0zyx6 = (Pr0zx6 & Xr0zx6);
assign Xr0zx6 = (~(Fs0zx6 & Voqyx6));
assign F00zx6 = (~(Klo7z6[1] & Ns0zx6));
assign Ns0zx6 = (~(Vs0zx6 & Dt0zx6));
assign Dt0zx6 = (Lt0zx6 & Tt0zx6);
assign Tt0zx6 = (Bu0zx6 & Ju0zx6);
assign Ju0zx6 = (Ru0zx6 & Zu0zx6);
assign Zu0zx6 = (~(Pdq7z6[5] & Oka8x6));
assign Ru0zx6 = (Hv0zx6 & Pv0zx6);
assign Pv0zx6 = (~(Kfq7z6[5] & S7hiw6));
assign Hv0zx6 = (~(Tbq7z6[5] & Qsgiw6));
assign Bu0zx6 = (Xv0zx6 & Fw0zx6);
assign Fw0zx6 = (~(Hhq7z6[5] & Ydliw6));
assign Xv0zx6 = (~(Cjq7z6[5] & Cza8x6));
assign Lt0zx6 = (Nw0zx6 & Vw0zx6);
assign Vw0zx6 = (Dx0zx6 & Lx0zx6);
assign Lx0zx6 = (~(T9tyx6 & Uu77z6));
assign Dx0zx6 = (~(X9q7z6[0] & B6qyx6));
assign Nw0zx6 = (Tx0zx6 & By0zx6);
assign By0zx6 = (~(D5qyx6 & Bqp7z6[5]));
assign Tx0zx6 = (~(Dm2ft6 & P3a8x6));
assign Vs0zx6 = (Jy0zx6 & Ry0zx6);
assign Ry0zx6 = (Zy0zx6 & Hz0zx6);
assign Hz0zx6 = (Pz0zx6 & Xz0zx6);
assign Xz0zx6 = (~(Fcqyx6 & B2q7z6[5]));
assign Pz0zx6 = (F01zx6 & N01zx6);
assign N01zx6 = (~(Ei2ft6 & Ua9ov6));
assign F01zx6 = (~(L9qyx6 & E6p7z6[5]));
assign Zy0zx6 = (V01zx6 & D11zx6);
assign D11zx6 = (~(M12ft6 & Nao7x6));
assign V01zx6 = (~(Gs2ft6 & Q0a8x6));
assign Jy0zx6 = (L11zx6 & T11zx6);
assign T11zx6 = (B21zx6 & J21zx6);
assign J21zx6 = (~(Tdqyx6 & Mkp7z6[5]));
assign B21zx6 = (~(U9p7z6[5] & Hfqyx6));
assign L11zx6 = (R21zx6 & Fgtyx6);
assign Fgtyx6 = (Ravyx6 & Z21zx6);
assign Z21zx6 = (~(Z6tyx6 & J2qyx6));
assign Zyzyx6 = (H31zx6 & H3zyx6);
assign H3zyx6 = (P31zx6 & X31zx6);
assign X31zx6 = (F41zx6 | Pnryx6);
assign Pnryx6 = (~(N41zx6 | Xfxyx6));
assign Xfxyx6 = (V41zx6 & D51zx6);
assign D51zx6 = (L51zx6 & Xruyx6);
assign P31zx6 = (~(T51zx6 & B61zx6));
assign B61zx6 = (J61zx6 & Z6wyx6);
assign J61zx6 = (~(Ti2nz6[1] & Bmvyx6));
assign T51zx6 = (J2uyx6 & F0pyx6);
assign H31zx6 = (R61zx6 & Z61zx6);
assign Z61zx6 = (~(Au1nz6[5] & Xjtyx6));
assign R61zx6 = (~(Ies7z6[5] & Tltyx6));
assign H7zyx6 = (~(Zmoyx6 & R8e7x6));
assign R8e7x6 = (~(H71zx6 & P71zx6));
assign P71zx6 = (~(Xnoyx6 & Oda7z6));
assign Oda7z6 = (~(X71zx6 & F81zx6));
assign F81zx6 = (~(HRDATAD[5] & Qln7z6[0]));
assign X71zx6 = (~(HRDATAS[5] & Qln7z6[1]));
assign H71zx6 = (~(Tim7z6[5] & Tpoyx6));
assign R6zyx6 = (N81zx6 & V81zx6);
assign V81zx6 = (~(HRDATAS[5] & Ad47x6));
assign N81zx6 = (~(HRDATAD[5] & Mc47x6));
assign B6zyx6 = (~(Lpryx6 & Zsq7x6));
assign Apo7v6 = (~(D91zx6 & L91zx6));
assign L91zx6 = (~(Jexmz6[6] & K94iw6));
assign D91zx6 = (T91zx6 & Ba1zx6);
assign Ba1zx6 = (~(Lloyx6 & Cx67x6));
assign Cx67x6 = (~(Ja1zx6 & Ra1zx6));
assign Ra1zx6 = (Za1zx6 & Hb1zx6);
assign Hb1zx6 = (Bqoyx6 | Xbe7x6);
assign Xbe7x6 = (Pb1zx6 & Xb1zx6);
assign Xb1zx6 = (Fc1zx6 & Nc1zx6);
assign Nc1zx6 = (Vc1zx6 & Dd1zx6);
assign Dd1zx6 = (~(D1pyx6 & Ld1zx6));
assign Ld1zx6 = (~(Td1zx6 & Be1zx6));
assign Be1zx6 = (Je1zx6 & Re1zx6);
assign Re1zx6 = (Ze1zx6 & Z6yyx6);
assign Ze1zx6 = (~(Hf1zx6 & Fy67v6));
assign Hf1zx6 = (Pbpyx6 & Zshiw6);
assign Je1zx6 = (Pf1zx6 & Xf1zx6);
assign Xf1zx6 = (~(Ag77z6 & Vcpyx6));
assign Pf1zx6 = (~(Biymz6[6] & Ddpyx6));
assign Td1zx6 = (Fg1zx6 & Ng1zx6);
assign Ng1zx6 = (Vg1zx6 & Y0jhy6);
assign Y0jhy6 = (~(Feymz6[2] & Fgpyx6));
assign Vg1zx6 = (~(Sgymz6[3] & Ngpyx6));
assign Fg1zx6 = (G1jhy6 & O1jhy6);
assign O1jhy6 = (~(Ojymz6[3] & Hfpyx6));
assign G1jhy6 = (~(Unymz6[3] & Thpyx6));
assign Vc1zx6 = (W1jhy6 & E2jhy6);
assign E2jhy6 = (~(M2jhy6 & U2jhy6));
assign M2jhy6 = (C3jhy6 & K3jhy6);
assign C3jhy6 = (~(S3jhy6 & A4jhy6));
assign A4jhy6 = (I4jhy6 & Q4jhy6);
assign Q4jhy6 = (Y4jhy6 & G5jhy6);
assign G5jhy6 = (~(Hyj7z6[3] & Tobiw6));
assign Y4jhy6 = (~(Hyj7z6[2] & Mobiw6));
assign I4jhy6 = (O5jhy6 & W5jhy6);
assign W5jhy6 = (~(Hyj7z6[1] & Fobiw6));
assign O5jhy6 = (~(Hyj7z6[5] & Apbiw6));
assign S3jhy6 = (E6jhy6 & M6jhy6);
assign M6jhy6 = (U6jhy6 & C7jhy6);
assign C7jhy6 = (~(Hyj7z6[6] & Hpbiw6));
assign U6jhy6 = (~(Hyj7z6[7] & Opbiw6));
assign E6jhy6 = (K7jhy6 & S7jhy6);
assign S7jhy6 = (~(Hyj7z6[0] & Dfk7z6[6]));
assign K7jhy6 = (~(Hyj7z6[4] & Jkl7z6[6]));
assign W1jhy6 = (~(P3uyx6 & Pk1nz6[6]));
assign P3uyx6 = (A8jhy6 & Klo7z6[3]);
assign Fc1zx6 = (I8jhy6 & Q8jhy6);
assign Q8jhy6 = (~(Klo7z6[1] & Y8jhy6));
assign Y8jhy6 = (~(G9jhy6 & O9jhy6));
assign O9jhy6 = (W9jhy6 & Eajhy6);
assign Eajhy6 = (Majhy6 & Uajhy6);
assign Uajhy6 = (Cbjhy6 & Ravyx6);
assign Cbjhy6 = (~(Kfq7z6[6] & S7hiw6));
assign Majhy6 = (Kbjhy6 & Sbjhy6);
assign Sbjhy6 = (~(Tbq7z6[6] & Qsgiw6));
assign Kbjhy6 = (~(Pdq7z6[6] & Oka8x6));
assign W9jhy6 = (Acjhy6 & Icjhy6);
assign Icjhy6 = (~(R6tyx6 & Qcjhy6));
assign Acjhy6 = (Ycjhy6 & Gdjhy6);
assign Gdjhy6 = (~(Hhq7z6[6] & Ydliw6));
assign Ycjhy6 = (~(Cjq7z6[6] & Cza8x6));
assign G9jhy6 = (Odjhy6 & Wdjhy6);
assign Wdjhy6 = (Eejhy6 & Mejhy6);
assign Mejhy6 = (Uejhy6 & Cfjhy6);
assign Cfjhy6 = (~(T9tyx6 & Mu77z6));
assign Uejhy6 = (~(X9q7z6[1] & B6qyx6));
assign Eejhy6 = (Kfjhy6 & Sfjhy6);
assign Sfjhy6 = (~(D5qyx6 & Bqp7z6[6]));
assign Kfjhy6 = (~(L9qyx6 & E6p7z6[6]));
assign Odjhy6 = (Agjhy6 & Igjhy6);
assign Igjhy6 = (~(U9p7z6[6] & Hfqyx6));
assign Agjhy6 = (Qgjhy6 & Ygjhy6);
assign Ygjhy6 = (~(Fcqyx6 & B2q7z6[6]));
assign Qgjhy6 = (~(Tdqyx6 & Mkp7z6[6]));
assign I8jhy6 = (Ghjhy6 & Ohjhy6);
assign Ohjhy6 = (~(Whjhy6 & Ngqyx6));
assign Whjhy6 = (~(Eijhy6 & Mijhy6));
assign Mijhy6 = (Uijhy6 & Cjjhy6);
assign Cjjhy6 = (Kjjhy6 & Sjjhy6);
assign Sjjhy6 = (Akjhy6 & Ikjhy6);
assign Ikjhy6 = (Qkjhy6 & Ykjhy6);
assign Ykjhy6 = (~(A0j7z6[6] & Xrqyx6));
assign Qkjhy6 = (Gljhy6 & Oljhy6);
assign Oljhy6 = (~(Wljhy6 & Lpyyx6));
assign Wljhy6 = (Koaiw6 & Jyuyx6);
assign Gljhy6 = (~(V40zx6 & Ffj7z6[1]));
assign Akjhy6 = (Emjhy6 & Mmjhy6);
assign Mmjhy6 = (~(H1j7z6[6] & Rqqyx6));
assign Emjhy6 = (~(Zudet6 & Ttqyx6));
assign Kjjhy6 = (Umjhy6 & Cnjhy6);
assign Cnjhy6 = (Knjhy6 & Snjhy6);
assign Snjhy6 = (~(Dxqyx6 & Nob7z6[6]));
assign Knjhy6 = (~(Wui7z6[6] & Lxqyx6));
assign Umjhy6 = (Aojhy6 & Iojhy6);
assign Iojhy6 = (~(Dri7z6[6] & Fwqyx6));
assign Aojhy6 = (~(Bwi7z6[6] & Hzqyx6));
assign Uijhy6 = (Qojhy6 & Yojhy6);
assign Yojhy6 = (Gpjhy6 & Opjhy6);
assign Opjhy6 = (Wpjhy6 & Eqjhy6);
assign Eqjhy6 = (~(Ba0zx6 & Nbj7z6[1]));
assign Wpjhy6 = (~(D90zx6 & Lgj7z6[181]));
assign Gpjhy6 = (Mqjhy6 & Uqjhy6);
assign Uqjhy6 = (~(Za0zx6 & Lgj7z6[169]));
assign Mqjhy6 = (~(Hb0zx6 & Lgj7z6[157]));
assign Qojhy6 = (Crjhy6 & Krjhy6);
assign Krjhy6 = (Srjhy6 & Asjhy6);
assign Asjhy6 = (~(Vc0zx6 & Lgj7z6[145]));
assign Srjhy6 = (~(Dd0zx6 & Lgj7z6[133]));
assign Crjhy6 = (Isjhy6 & Qsjhy6);
assign Qsjhy6 = (~(Be0zx6 & Lgj7z6[121]));
assign Isjhy6 = (~(Je0zx6 & Lgj7z6[109]));
assign Eijhy6 = (Ysjhy6 & Gtjhy6);
assign Gtjhy6 = (Otjhy6 & Wtjhy6);
assign Wtjhy6 = (Eujhy6 & Mujhy6);
assign Mujhy6 = (Uujhy6 & Cvjhy6);
assign Cvjhy6 = (~(Bi0zx6 & Lgj7z6[97]));
assign Uujhy6 = (~(Ji0zx6 & Lgj7z6[85]));
assign Eujhy6 = (Kvjhy6 & Svjhy6);
assign Svjhy6 = (~(Dh0zx6 & Lgj7z6[73]));
assign Kvjhy6 = (~(Hj0zx6 & Lgj7z6[61]));
assign Otjhy6 = (Awjhy6 & Iwjhy6);
assign Iwjhy6 = (Qwjhy6 & Ywjhy6);
assign Ywjhy6 = (~(Pj0zx6 & Lgj7z6[49]));
assign Qwjhy6 = (~(Dl0zx6 & Lgj7z6[37]));
assign Awjhy6 = (Gxjhy6 & Oxjhy6);
assign Oxjhy6 = (~(Ll0zx6 & Lgj7z6[25]));
assign Gxjhy6 = (~(Jm0zx6 & Lgj7z6[13]));
assign Ysjhy6 = (Wxjhy6 & Eyjhy6);
assign Eyjhy6 = (Myjhy6 & Uyjhy6);
assign Uyjhy6 = (Czjhy6 & Kzjhy6);
assign Kzjhy6 = (~(Rm0zx6 & Lgj7z6[1]));
assign Czjhy6 = (~(Pzqyx6 & G5j7z6[38]));
assign Myjhy6 = (Szjhy6 & A0khy6);
assign A0khy6 = (~(Jyqyx6 & G5j7z6[6]));
assign Szjhy6 = (~(B2ryx6 & M6j7z6[38]));
assign Wxjhy6 = (I0khy6 & Q0khy6);
assign Q0khy6 = (Y0khy6 & G1khy6);
assign G1khy6 = (~(J2ryx6 & M6j7z6[6]));
assign Y0khy6 = (~(D1ryx6 & Ohj7z6[38]));
assign I0khy6 = (O1khy6 & W1khy6);
assign W1khy6 = (~(X3ryx6 & Ohj7z6[6]));
assign O1khy6 = (~(STCALIB[6] & F4ryx6));
assign Ghjhy6 = (~(Klo7z6[2] & E2khy6));
assign E2khy6 = (~(M2khy6 & U2khy6));
assign U2khy6 = (C3khy6 & K3khy6);
assign K3khy6 = (S3khy6 & A4khy6);
assign A4khy6 = (~(Ugtet6 & S4kiw6));
assign S3khy6 = (I4khy6 & Q4khy6);
assign Q4khy6 = (~(Nqo7z6[4] & M8kiw6));
assign I4khy6 = (~(Fpo7z6[4] & H9kiw6));
assign C3khy6 = (Y4khy6 & G5khy6);
assign G5khy6 = (~(Ouo7z6[4] & K7kiw6));
assign Y4khy6 = (~(Hxo7z6[4] & W6kiw6));
assign M2khy6 = (O5khy6 & W5khy6);
assign W5khy6 = (E6khy6 & M6khy6);
assign M6khy6 = (~(W3p7z6[6] & G5kiw6));
assign E6khy6 = (U6khy6 & C7khy6);
assign C7khy6 = (~(Vro7z6[4] & Y7kiw6));
assign U6khy6 = (~(T2p7z6[6] & U5kiw6));
assign O5khy6 = (Jyzyx6 & K7khy6);
assign K7khy6 = (~(A0p7z6[4] & I6kiw6));
assign Jyzyx6 = (S7khy6 & A8khy6);
assign Pb1zx6 = (I8khy6 & Q8khy6);
assign Q8khy6 = (Y8khy6 & G9khy6);
assign G9khy6 = (~(Oo1nz6[6] & Pjtyx6));
assign Y8khy6 = (O9khy6 & W9khy6);
assign W9khy6 = (Fotyx6 | Eakhy6);
assign Eakhy6 = (!F0pyx6);
assign O9khy6 = (R2zyx6 | Xruyx6);
assign I8khy6 = (Makhy6 & Uakhy6);
assign Uakhy6 = (~(Au1nz6[6] & Xjtyx6));
assign Makhy6 = (~(Ies7z6[6] & Tltyx6));
assign Za1zx6 = (~(Zmoyx6 & Ece7x6));
assign Ece7x6 = (~(Cbkhy6 & Kbkhy6));
assign Kbkhy6 = (~(Xnoyx6 & Gda7z6));
assign Gda7z6 = (~(Sbkhy6 & Ackhy6));
assign Ackhy6 = (~(HRDATAD[6] & Qln7z6[0]));
assign Sbkhy6 = (~(HRDATAS[6] & Qln7z6[1]));
assign Cbkhy6 = (~(Tim7z6[6] & Tpoyx6));
assign Ja1zx6 = (Ickhy6 & Qckhy6);
assign Qckhy6 = (~(HRDATAS[6] & Ad47x6));
assign Ickhy6 = (~(HRDATAD[6] & Mc47x6));
assign T91zx6 = (~(Lpryx6 & Lzq7x6));
assign Too7v6 = (~(Yckhy6 & Gdkhy6));
assign Gdkhy6 = (~(Jexmz6[7] & K94iw6));
assign Yckhy6 = (Odkhy6 & Wdkhy6);
assign Wdkhy6 = (~(Lloyx6 & Hp67x6));
assign Hp67x6 = (~(Eekhy6 & Mekhy6));
assign Mekhy6 = (Uekhy6 & Cfkhy6);
assign Cfkhy6 = (Bqoyx6 | Kfe7x6);
assign Kfe7x6 = (Kfkhy6 & Sfkhy6);
assign Sfkhy6 = (Agkhy6 & Igkhy6);
assign Igkhy6 = (Qgkhy6 & R2zyx6);
assign R2zyx6 = (~(Ygkhy6 & Ghkhy6));
assign Ghkhy6 = (~(Hnryx6 | Ohkhy6));
assign Ygkhy6 = (Klo7z6[0] & Or27v6);
assign Qgkhy6 = (~(Whkhy6 & U2jhy6));
assign Whkhy6 = (Eikhy6 & K3jhy6);
assign Eikhy6 = (~(Mikhy6 & Uikhy6));
assign Uikhy6 = (Cjkhy6 & Kjkhy6);
assign Kjkhy6 = (Sjkhy6 & Akkhy6);
assign Akkhy6 = (~(Hyj7z6[3] & Lrbiw6));
assign Sjkhy6 = (~(Hyj7z6[2] & Xqbiw6));
assign Cjkhy6 = (Ikkhy6 & Qkkhy6);
assign Qkkhy6 = (~(Hyj7z6[1] & Jqbiw6));
assign Ikkhy6 = (~(Hyj7z6[5] & Gsbiw6));
assign Mikhy6 = (Ykkhy6 & Glkhy6);
assign Glkhy6 = (Olkhy6 & Wlkhy6);
assign Wlkhy6 = (~(Hyj7z6[6] & Usbiw6));
assign Olkhy6 = (~(Hyj7z6[7] & Btbiw6));
assign Ykkhy6 = (Emkhy6 & Mmkhy6);
assign Mmkhy6 = (~(Hyj7z6[0] & Dfk7z6[7]));
assign Emkhy6 = (~(Hyj7z6[4] & Jkl7z6[7]));
assign Agkhy6 = (Umkhy6 & Cnkhy6);
assign Cnkhy6 = (~(Knkhy6 & Ngqyx6));
assign Knkhy6 = (~(Snkhy6 & Aokhy6));
assign Aokhy6 = (Iokhy6 & Qokhy6);
assign Qokhy6 = (Yokhy6 & Gpkhy6);
assign Gpkhy6 = (Opkhy6 & Wpkhy6);
assign Wpkhy6 = (Eqkhy6 & Mqkhy6);
assign Mqkhy6 = (~(A0j7z6[7] & Xrqyx6));
assign Eqkhy6 = (Uqkhy6 & Crkhy6);
assign Crkhy6 = (~(Prqyx6 & Z3j7z6[7]));
assign Uqkhy6 = (~(V40zx6 & Ffj7z6[2]));
assign Opkhy6 = (Krkhy6 & Srkhy6);
assign Srkhy6 = (~(H1j7z6[7] & Rqqyx6));
assign Krkhy6 = (~(Ywdet6 & Ttqyx6));
assign Yokhy6 = (Askhy6 & Iskhy6);
assign Iskhy6 = (Qskhy6 & Yskhy6);
assign Yskhy6 = (~(Bzi7z6[7] & Vsqyx6));
assign Qskhy6 = (~(Dxqyx6 & Nob7z6[7]));
assign Askhy6 = (Gtkhy6 & Otkhy6);
assign Otkhy6 = (~(Wui7z6[7] & Lxqyx6));
assign Gtkhy6 = (~(Dri7z6[7] & Fwqyx6));
assign Iokhy6 = (Wtkhy6 & Eukhy6);
assign Eukhy6 = (Mukhy6 & Uukhy6);
assign Uukhy6 = (Cvkhy6 & Kvkhy6);
assign Kvkhy6 = (~(Qti7z6[7] & Svkhy6));
assign Cvkhy6 = (Awkhy6 & Iwkhy6);
assign Iwkhy6 = (~(Bwi7z6[7] & Hzqyx6));
assign Awkhy6 = (~(Ba0zx6 & Nbj7z6[2]));
assign Mukhy6 = (Qwkhy6 & Ywkhy6);
assign Ywkhy6 = (~(D90zx6 & Lgj7z6[182]));
assign Qwkhy6 = (~(Za0zx6 & Lgj7z6[170]));
assign Wtkhy6 = (Gxkhy6 & Oxkhy6);
assign Oxkhy6 = (Wxkhy6 & Eykhy6);
assign Eykhy6 = (~(Hb0zx6 & Lgj7z6[158]));
assign Wxkhy6 = (~(Vc0zx6 & Lgj7z6[146]));
assign Gxkhy6 = (Mykhy6 & Uykhy6);
assign Uykhy6 = (~(Dd0zx6 & Lgj7z6[134]));
assign Mykhy6 = (~(Be0zx6 & Lgj7z6[122]));
assign Snkhy6 = (Czkhy6 & Kzkhy6);
assign Kzkhy6 = (Szkhy6 & A0lhy6);
assign A0lhy6 = (I0lhy6 & Q0lhy6);
assign Q0lhy6 = (Y0lhy6 & G1lhy6);
assign G1lhy6 = (~(Ji0zx6 & Lgj7z6[86]));
assign Y0lhy6 = (O1lhy6 & W1lhy6);
assign W1lhy6 = (~(Je0zx6 & Lgj7z6[110]));
assign O1lhy6 = (~(Bi0zx6 & Lgj7z6[98]));
assign I0lhy6 = (E2lhy6 & M2lhy6);
assign M2lhy6 = (~(Dh0zx6 & Lgj7z6[74]));
assign E2lhy6 = (~(Hj0zx6 & Lgj7z6[62]));
assign Szkhy6 = (U2lhy6 & C3lhy6);
assign C3lhy6 = (K3lhy6 & S3lhy6);
assign S3lhy6 = (~(Pj0zx6 & Lgj7z6[50]));
assign K3lhy6 = (~(Dl0zx6 & Lgj7z6[38]));
assign U2lhy6 = (A4lhy6 & I4lhy6);
assign I4lhy6 = (~(Ll0zx6 & Lgj7z6[26]));
assign A4lhy6 = (~(Jm0zx6 & Lgj7z6[14]));
assign Czkhy6 = (Q4lhy6 & Y4lhy6);
assign Y4lhy6 = (G5lhy6 & O5lhy6);
assign O5lhy6 = (W5lhy6 & E6lhy6);
assign E6lhy6 = (~(Jyqyx6 & G5j7z6[7]));
assign W5lhy6 = (M6lhy6 & U6lhy6);
assign U6lhy6 = (~(Rm0zx6 & Lgj7z6[2]));
assign M6lhy6 = (~(Pzqyx6 & G5j7z6[39]));
assign G5lhy6 = (C7lhy6 & K7lhy6);
assign K7lhy6 = (~(B2ryx6 & M6j7z6[39]));
assign C7lhy6 = (~(J2ryx6 & M6j7z6[7]));
assign Q4lhy6 = (S7lhy6 & A8lhy6);
assign A8lhy6 = (I8lhy6 & Q8lhy6);
assign Q8lhy6 = (~(D1ryx6 & Ohj7z6[39]));
assign I8lhy6 = (~(X3ryx6 & Ohj7z6[7]));
assign S7lhy6 = (Hr0zx6 & Y8lhy6);
assign Y8lhy6 = (~(STCALIB[7] & F4ryx6));
assign Hr0zx6 = (Hjqyx6 & G9lhy6);
assign G9lhy6 = (~(Lpyyx6 & Jyuyx6));
assign Hjqyx6 = (~(O9lhy6 & Koaiw6));
assign O9lhy6 = (Hjsyx6 & Jyuyx6);
assign Jyuyx6 = (Dxuyx6 & Toi7z6[5]);
assign Dxuyx6 = (W9lhy6 & Ealhy6);
assign W9lhy6 = (~(Malhy6 | Ualhy6));
assign Umkhy6 = (~(Klo7z6[1] & Cblhy6));
assign Cblhy6 = (~(Kblhy6 & Sblhy6));
assign Sblhy6 = (Aclhy6 & Iclhy6);
assign Iclhy6 = (Qclhy6 & Yclhy6);
assign Yclhy6 = (Gdlhy6 & Ravyx6);
assign Gdlhy6 = (~(Kfq7z6[7] & S7hiw6));
assign S7hiw6 = (~(Odlhy6 | Wdlhy6));
assign Qclhy6 = (Eelhy6 & Melhy6);
assign Melhy6 = (~(Tbq7z6[7] & Qsgiw6));
assign Qsgiw6 = (B2qyx6 & Uelhy6);
assign Uelhy6 = (!Cflhy6);
assign Eelhy6 = (~(Pdq7z6[7] & Oka8x6));
assign Oka8x6 = (~(Odlhy6 | Kflhy6));
assign Aclhy6 = (Sflhy6 & Aglhy6);
assign Aglhy6 = (Iglhy6 & Qglhy6);
assign Qglhy6 = (~(Hhq7z6[7] & Ydliw6));
assign Ydliw6 = (~(Yglhy6 | Cflhy6));
assign Iglhy6 = (~(Cjq7z6[7] & Cza8x6));
assign Cza8x6 = (~(Cflhy6 | Ghlhy6));
assign Sflhy6 = (Ohlhy6 & Whlhy6);
assign Whlhy6 = (~(T9tyx6 & Eu77z6));
assign Ohlhy6 = (~(X9q7z6[2] & B6qyx6));
assign Kblhy6 = (Eilhy6 & Milhy6);
assign Milhy6 = (Uilhy6 & Cjlhy6);
assign Cjlhy6 = (Kjlhy6 & Sjlhy6);
assign Sjlhy6 = (~(D5qyx6 & Bqp7z6[7]));
assign Kjlhy6 = (~(L9qyx6 & E6p7z6[7]));
assign Uilhy6 = (Aklhy6 & Iklhy6);
assign Iklhy6 = (~(Fcqyx6 & B2q7z6[7]));
assign Aklhy6 = (~(Nao7x6 & W22ft6));
assign Eilhy6 = (Qklhy6 & R21zx6);
assign R21zx6 = (T1qyx6 & Yklhy6);
assign Yklhy6 = (~(R6tyx6 & Bxeiw6));
assign R6tyx6 = (Gllhy6 & Af4ft6);
assign T1qyx6 = (~(Qcjhy6 & J2qyx6));
assign J2qyx6 = (~(Ollhy6 | Zveiw6));
assign Zveiw6 = (!Af4ft6);
assign Ollhy6 = (~(Nmq7z6[5] & Nmq7z6[3]));
assign Qklhy6 = (Wllhy6 & Emlhy6);
assign Emlhy6 = (~(Tdqyx6 & Mkp7z6[7]));
assign Wllhy6 = (~(U9p7z6[7] & Hfqyx6));
assign Kfkhy6 = (Mmlhy6 & Umlhy6);
assign Umlhy6 = (Cnlhy6 & Knlhy6);
assign Knlhy6 = (~(Klo7z6[3] & Snlhy6));
assign Snlhy6 = (~(Aolhy6 & Iolhy6));
assign Iolhy6 = (Qolhy6 & Yolhy6);
assign Yolhy6 = (~(Mphiw6 & Gplhy6));
assign Gplhy6 = (~(Oplhy6 & Wplhy6));
assign Wplhy6 = (Eqlhy6 & Mqlhy6);
assign Mqlhy6 = (Uqlhy6 & Crlhy6);
assign Crlhy6 = (~(Pbpyx6 & Zshiw6));
assign Zshiw6 = (Krlhy6 & Srlhy6);
assign Srlhy6 = (Xfymz6[5] & Aslhy6);
assign Krlhy6 = (L9pyx6 & Xfymz6[7]);
assign Uqlhy6 = (~(Biymz6[7] & Ddpyx6));
assign Eqlhy6 = (Islhy6 & Qslhy6);
assign Qslhy6 = (~(Vv67v6 & Fgpyx6));
assign Islhy6 = (~(Sgymz6[4] & Ngpyx6));
assign Oplhy6 = (Yslhy6 & N4yyx6);
assign N4yyx6 = (Pjpyx6 & Gtlhy6);
assign Gtlhy6 = (~(N8pyx6 & Xbpyx6));
assign Pjpyx6 = (Z2xyx6 & Otlhy6);
assign Otlhy6 = (~(Wtlhy6 & Eulhy6));
assign Eulhy6 = (Xfymz6[2] & Xbpyx6);
assign Wtlhy6 = (Xfymz6[4] & Xfymz6[3]);
assign Z2xyx6 = (~(J2xyx6 & Xbpyx6));
assign Xbpyx6 = (L9pyx6 & Mulhy6);
assign Yslhy6 = (Uulhy6 & Cvlhy6);
assign Cvlhy6 = (~(Ojymz6[4] & Hfpyx6));
assign Uulhy6 = (~(Unymz6[4] & Thpyx6));
assign Qolhy6 = (Kvlhy6 & Svlhy6);
assign Svlhy6 = (~(Kniiw6 & Awlhy6));
assign Awlhy6 = (~(Hbzyx6 & Ruxyx6));
assign Ruxyx6 = (~(Iwlhy6 & J02nz6[5]));
assign Iwlhy6 = (B2wyx6 & J02nz6[2]);
assign B2wyx6 = (!T5uyx6);
assign T5uyx6 = (~(Qwlhy6 & Ywlhy6));
assign Qwlhy6 = (J02nz6[4] & Xvxyx6);
assign Hbzyx6 = (Gxlhy6 & Vwxyx6);
assign Vwxyx6 = (~(Oxlhy6 & J02nz6[2]));
assign Oxlhy6 = (!Fopyx6);
assign Fopyx6 = (~(Wxlhy6 & Tppyx6));
assign Wxlhy6 = (J02nz6[4] & J02nz6[8]);
assign Gxlhy6 = (L1wyx6 & Eylhy6);
assign L1wyx6 = (~(Mylhy6 & Pbzyx6));
assign Pbzyx6 = (Uylhy6 & Ywlhy6);
assign Ywlhy6 = (~(Czlhy6 | J02nz6[3]));
assign Uylhy6 = (J02nz6[5] & Xvxyx6);
assign Mylhy6 = (J02nz6[2] & Puhiw6);
assign Kvlhy6 = (~(Kzlhy6 & Szlhy6));
assign Szlhy6 = (~(Fotyx6 & A0mhy6));
assign A0mhy6 = (~(J2uyx6 & I0mhy6));
assign I0mhy6 = (~(Q0mhy6 & Y0mhy6));
assign Y0mhy6 = (~(Ti2nz6[1] & Ti2nz6[2]));
assign J2uyx6 = (~(B2uyx6 | G1mhy6));
assign Fotyx6 = (~(Pfxyx6 & O1mhy6));
assign Pfxyx6 = (~(G1mhy6 | Ti2nz6[0]));
assign G1mhy6 = (~(Ti2nz6[3] & Xzoyx6));
assign Xzoyx6 = (~(W1mhy6 | Ti2nz6[4]));
assign Aolhy6 = (E2mhy6 & M2mhy6);
assign M2mhy6 = (~(Oo1nz6[7] & U2mhy6));
assign E2mhy6 = (C3mhy6 & K3mhy6);
assign K3mhy6 = (~(Pk1nz6[7] & A8jhy6));
assign C3mhy6 = (~(Au1nz6[7] & S3mhy6));
assign Cnlhy6 = (~(Klo7z6[2] & A4mhy6));
assign A4mhy6 = (~(I4mhy6 & Q4mhy6));
assign Q4mhy6 = (Y4mhy6 & G5mhy6);
assign G5mhy6 = (O5mhy6 & W5mhy6);
assign W5mhy6 = (~(Fpo7z6[5] & H9kiw6));
assign O5mhy6 = (E6mhy6 & A8khy6);
assign A8khy6 = (~(Pfuyx6 & M6mhy6));
assign E6mhy6 = (~(Nqo7z6[5] & M8kiw6));
assign Y4mhy6 = (U6mhy6 & C7mhy6);
assign C7mhy6 = (~(Hxo7z6[5] & W6kiw6));
assign U6mhy6 = (K7mhy6 & S7mhy6);
assign S7mhy6 = (~(Tetet6 & S4kiw6));
assign K7mhy6 = (~(Ouo7z6[5] & K7kiw6));
assign I4mhy6 = (A8mhy6 & I8mhy6);
assign I8mhy6 = (Q8mhy6 & Y8mhy6);
assign Y8mhy6 = (~(W3p7z6[7] & G5kiw6));
assign Q8mhy6 = (G9mhy6 & O9mhy6);
assign O9mhy6 = (~(Vro7z6[5] & Y7kiw6));
assign G9mhy6 = (~(T2p7z6[7] & U5kiw6));
assign A8mhy6 = (Tlyyx6 & W9mhy6);
assign W9mhy6 = (~(A0p7z6[5] & I6kiw6));
assign Tlyyx6 = (~(Z6ryx6 | Eamhy6));
assign Eamhy6 = (Mamhy6 & M6mhy6);
assign Mamhy6 = (Uamhy6 & R2syx6);
assign Z6ryx6 = (Cbmhy6 & Z4p7z6[2]);
assign Cbmhy6 = (Z4p7z6[1] & M6mhy6);
assign M6mhy6 = (~(Hfuyx6 | Ruzyx6));
assign Ruzyx6 = (~(Kbmhy6 & Z4p7z6[5]));
assign Kbmhy6 = (Z4p7z6[3] & Upeiw6);
assign Upeiw6 = (!Z4p7z6[4]);
assign Mmlhy6 = (Sbmhy6 & Acmhy6);
assign Acmhy6 = (~(N41zx6 & Klo7z6[0]));
assign N41zx6 = (Icmhy6 & V41zx6);
assign V41zx6 = (~(Hnryx6 | Pruyx6));
assign Hnryx6 = (Tt4yx6 | Zauyx6);
assign Zauyx6 = (~(Qcmhy6 & Zfs7z6[8]));
assign Qcmhy6 = (Mm27v6 & Zfs7z6[7]);
assign Icmhy6 = (Or27v6 & Ap27v6);
assign Sbmhy6 = (~(Ies7z6[7] & Tltyx6));
assign Uekhy6 = (~(Zmoyx6 & Rfe7x6));
assign Rfe7x6 = (~(Ycmhy6 & Gdmhy6));
assign Gdmhy6 = (~(Yca7z6 & Xnoyx6));
assign Xnoyx6 = (~(Odmhy6 & Wdmhy6));
assign Odmhy6 = (~(Eemhy6 & Memhy6));
assign Yca7z6 = (~(Uemhy6 & Cfmhy6));
assign Cfmhy6 = (~(HRDATAD[7] & Qln7z6[0]));
assign Uemhy6 = (~(HRDATAS[7] & Qln7z6[1]));
assign Ycmhy6 = (~(Tim7z6[7] & Tpoyx6));
assign Tpoyx6 = (~(Memhy6 | Kfmhy6));
assign Memhy6 = (~(Sfmhy6 & Yxixx6));
assign Sfmhy6 = (~(Jkqnv6 | Ven7z6[0]));
assign Eekhy6 = (Agmhy6 & Igmhy6);
assign Igmhy6 = (~(HRDATAS[7] & Ad47x6));
assign Agmhy6 = (~(HRDATAD[7] & Mc47x6));
assign Odkhy6 = (~(Lpryx6 & Kwp7x6));
assign Moo7v6 = (~(Qgmhy6 & Ygmhy6));
assign Ygmhy6 = (~(Jexmz6[8] & K94iw6));
assign Qgmhy6 = (Ghmhy6 & Ohmhy6);
assign Ohmhy6 = (~(Lloyx6 & Jf9ov6));
assign Jf9ov6 = (~(Whmhy6 & Eimhy6));
assign Eimhy6 = (Mimhy6 & Uimhy6);
assign Uimhy6 = (Bqoyx6 | Xaf7x6);
assign Xaf7x6 = (Cjmhy6 & Kjmhy6);
assign Kjmhy6 = (Sjmhy6 & Akmhy6);
assign Akmhy6 = (Ikmhy6 & Qkmhy6);
assign Qkmhy6 = (~(Rmzyx6 & Ykmhy6));
assign Ykmhy6 = (~(Glmhy6 & Olmhy6));
assign Olmhy6 = (Wlmhy6 & Emmhy6);
assign Emmhy6 = (Mmmhy6 & Ummhy6);
assign Ummhy6 = (~(Hyj7z6[0] & Dfk7z6[8]));
assign Mmmhy6 = (~(Hyj7z6[1] & Lpk7z6[8]));
assign Wlmhy6 = (Cnmhy6 & Knmhy6);
assign Knmhy6 = (~(Hyj7z6[2] & Tzk7z6[8]));
assign Cnmhy6 = (~(Hyj7z6[3] & Bal7z6[8]));
assign Glmhy6 = (Snmhy6 & Aomhy6);
assign Aomhy6 = (Iomhy6 & Qomhy6);
assign Qomhy6 = (~(Hyj7z6[4] & Jkl7z6[8]));
assign Iomhy6 = (~(Hyj7z6[5] & Rul7z6[8]));
assign Snmhy6 = (Yomhy6 & Gpmhy6);
assign Gpmhy6 = (~(Hyj7z6[6] & Z4m7z6[8]));
assign Yomhy6 = (~(Hyj7z6[7] & Hfm7z6[8]));
assign Ikmhy6 = (~(Xbzyx6 & Opmhy6));
assign Opmhy6 = (~(Wpmhy6 & Eqmhy6));
assign Eqmhy6 = (Mqmhy6 & Uqmhy6);
assign Uqmhy6 = (Crmhy6 & Krmhy6);
assign Krmhy6 = (~(Hyj7z6[0] & Rbk7z6[6]));
assign Crmhy6 = (~(Hyj7z6[1] & Zlk7z6[6]));
assign Mqmhy6 = (Srmhy6 & Asmhy6);
assign Asmhy6 = (~(Hyj7z6[2] & Hwk7z6[6]));
assign Srmhy6 = (~(Hyj7z6[3] & P6l7z6[6]));
assign Wpmhy6 = (Ismhy6 & Qsmhy6);
assign Qsmhy6 = (Ysmhy6 & Gtmhy6);
assign Gtmhy6 = (~(Hyj7z6[4] & Xgl7z6[6]));
assign Ysmhy6 = (~(Hyj7z6[5] & Frl7z6[6]));
assign Ismhy6 = (Otmhy6 & Wtmhy6);
assign Wtmhy6 = (~(Hyj7z6[6] & N1m7z6[6]));
assign Otmhy6 = (~(Hyj7z6[7] & Vbm7z6[6]));
assign Sjmhy6 = (Eumhy6 & Mumhy6);
assign Mumhy6 = (~(Uumhy6 & Ngqyx6));
assign Uumhy6 = (~(Cvmhy6 & Kvmhy6));
assign Kvmhy6 = (Svmhy6 & Awmhy6);
assign Awmhy6 = (Iwmhy6 & Qwmhy6);
assign Qwmhy6 = (Ywmhy6 & Gxmhy6);
assign Gxmhy6 = (~(Hnqyx6 & Fuadt6));
assign Ywmhy6 = (Dhsyx6 & Bqyyx6);
assign Iwmhy6 = (Oxmhy6 & Wxmhy6);
assign Wxmhy6 = (~(H1j7z6[8] & Rqqyx6));
assign Oxmhy6 = (Eymhy6 & Mymhy6);
assign Mymhy6 = (~(Prqyx6 & Z3j7z6[8]));
assign Eymhy6 = (~(A0j7z6[8] & Xrqyx6));
assign Svmhy6 = (Uymhy6 & Czmhy6);
assign Czmhy6 = (Kzmhy6 & Szmhy6);
assign Szmhy6 = (~(Dxqyx6 & Nob7z6[8]));
assign Kzmhy6 = (A0nhy6 & I0nhy6);
assign I0nhy6 = (~(Yydet6 & Ttqyx6));
assign A0nhy6 = (~(Bzi7z6[8] & Vsqyx6));
assign Uymhy6 = (Q0nhy6 & Y0nhy6);
assign Y0nhy6 = (~(Wui7z6[8] & Lxqyx6));
assign Q0nhy6 = (~(Dri7z6[8] & Fwqyx6));
assign Cvmhy6 = (G1nhy6 & O1nhy6);
assign O1nhy6 = (W1nhy6 & E2nhy6);
assign E2nhy6 = (M2nhy6 & U2nhy6);
assign U2nhy6 = (~(Pzqyx6 & G5j7z6[40]));
assign M2nhy6 = (C3nhy6 & K3nhy6);
assign K3nhy6 = (~(Bwi7z6[8] & Hzqyx6));
assign C3nhy6 = (~(Qti7z6[8] & Svkhy6));
assign W1nhy6 = (S3nhy6 & A4nhy6);
assign A4nhy6 = (~(Jyqyx6 & G5j7z6[8]));
assign S3nhy6 = (~(B2ryx6 & M6j7z6[40]));
assign G1nhy6 = (I4nhy6 & Q4nhy6);
assign Q4nhy6 = (Y4nhy6 & G5nhy6);
assign G5nhy6 = (~(O5nhy6 & Hsi7z6[0]));
assign Y4nhy6 = (W5nhy6 & E6nhy6);
assign E6nhy6 = (~(J2ryx6 & M6j7z6[8]));
assign W5nhy6 = (~(D1ryx6 & Ohj7z6[40]));
assign I4nhy6 = (M6nhy6 & U6nhy6);
assign U6nhy6 = (~(X3ryx6 & Ohj7z6[8]));
assign M6nhy6 = (~(STCALIB[8] & F4ryx6));
assign Eumhy6 = (~(Klo7z6[1] & C7nhy6));
assign C7nhy6 = (~(K7nhy6 & S7nhy6));
assign S7nhy6 = (A8nhy6 & I8nhy6);
assign I8nhy6 = (Q8nhy6 & Y8nhy6);
assign Y8nhy6 = (~(X9q7z6[3] & B6qyx6));
assign Q8nhy6 = (G9nhy6 & Ravyx6);
assign G9nhy6 = (~(T9tyx6 & Wt77z6));
assign A8nhy6 = (O9nhy6 & W9nhy6);
assign W9nhy6 = (~(D5qyx6 & Bqp7z6[8]));
assign O9nhy6 = (~(L9qyx6 & E6p7z6[8]));
assign K7nhy6 = (Eanhy6 & Manhy6);
assign Manhy6 = (Uanhy6 & Cbnhy6);
assign Cbnhy6 = (~(Fcqyx6 & B2q7z6[8]));
assign Uanhy6 = (~(Q0a8x6 & Cq2ft6));
assign Eanhy6 = (Kbnhy6 & Sbnhy6);
assign Sbnhy6 = (~(Tdqyx6 & Mkp7z6[8]));
assign Kbnhy6 = (~(U9p7z6[8] & Hfqyx6));
assign Cjmhy6 = (Acnhy6 & Icnhy6);
assign Icnhy6 = (Qcnhy6 & Ycnhy6);
assign Ycnhy6 = (~(Klo7z6[3] & Gdnhy6));
assign Gdnhy6 = (~(Odnhy6 & Wdnhy6));
assign Wdnhy6 = (Eenhy6 & Menhy6);
assign Menhy6 = (Uenhy6 & Cfnhy6);
assign Cfnhy6 = (~(Pk1nz6[8] & A8jhy6));
assign Uenhy6 = (Kfnhy6 & Sfnhy6);
assign Sfnhy6 = (~(Agnhy6 & Ignhy6));
assign Agnhy6 = (Mphiw6 & Tah7v6);
assign Kfnhy6 = (Jasyx6 | Qgnhy6);
assign Jasyx6 = (~(Ygnhy6 & Rgiiw6));
assign Rgiiw6 = (Ghnhy6 & Ohnhy6);
assign Ghnhy6 = (B6wyx6 & J02nz6[9]);
assign B6wyx6 = (~(Czlhy6 | J02nz6[4]));
assign Ygnhy6 = (J02nz6[2] & Jke7v6);
assign Eenhy6 = (Whnhy6 & Einhy6);
assign Einhy6 = (~(Ojymz6[5] & Minhy6));
assign Whnhy6 = (~(Unymz6[5] & Uinhy6));
assign Odnhy6 = (Cjnhy6 & Kjnhy6);
assign Kjnhy6 = (Sjnhy6 & Aknhy6);
assign Aknhy6 = (~(T077v6 & Iknhy6));
assign Sjnhy6 = (Qknhy6 & Yknhy6);
assign Yknhy6 = (~(Sgymz6[5] & Glnhy6));
assign Qknhy6 = (~(Biymz6[8] & Olnhy6));
assign Cjnhy6 = (Wlnhy6 & Emnhy6);
assign Emnhy6 = (~(Zs1nz6[0] & S3mhy6));
assign Wlnhy6 = (~(Nn1nz6[0] & U2mhy6));
assign Qcnhy6 = (~(Klo7z6[2] & Mmnhy6));
assign Mmnhy6 = (~(Umnhy6 & Cnnhy6));
assign Cnnhy6 = (Knnhy6 & Snnhy6);
assign Snnhy6 = (Aonhy6 & Ionhy6);
assign Ionhy6 = (~(Sctet6 & S4kiw6));
assign Aonhy6 = (Qonhy6 & Yonhy6);
assign Yonhy6 = (~(Nqo7z6[6] & M8kiw6));
assign Qonhy6 = (~(Fpo7z6[6] & H9kiw6));
assign Knnhy6 = (Gpnhy6 & Opnhy6);
assign Opnhy6 = (~(Ouo7z6[6] & K7kiw6));
assign Gpnhy6 = (~(Hxo7z6[6] & W6kiw6));
assign Umnhy6 = (Wpnhy6 & Eqnhy6);
assign Eqnhy6 = (Mqnhy6 & Uqnhy6);
assign Uqnhy6 = (~(Vro7z6[6] & Y7kiw6));
assign Mqnhy6 = (~(T2p7z6[8] & U5kiw6));
assign Wpnhy6 = (Crnhy6 & Krnhy6);
assign Krnhy6 = (~(W3p7z6[8] & G5kiw6));
assign Crnhy6 = (~(A0p7z6[6] & I6kiw6));
assign Acnhy6 = (Srnhy6 & Asnhy6);
assign Asnhy6 = (~(H56ft6 & Lltyx6));
assign Srnhy6 = (~(Ies7z6[8] & Tltyx6));
assign Mimhy6 = (~(Zmoyx6 & Ebf7x6));
assign Ebf7x6 = (~(Isnhy6 & Qsnhy6));
assign Qsnhy6 = (~(Ysnhy6 & Qca7z6));
assign Qca7z6 = (~(Gtnhy6 & Otnhy6));
assign Otnhy6 = (~(HRDATAD[8] & Qln7z6[0]));
assign Gtnhy6 = (~(HRDATAS[8] & Qln7z6[1]));
assign Isnhy6 = (Wtnhy6 & Eunhy6);
assign Eunhy6 = (~(Munhy6 & S7n7z6[0]));
assign Wtnhy6 = (~(Tim7z6[8] & Uunhy6));
assign Whmhy6 = (Cvnhy6 & Kvnhy6);
assign Kvnhy6 = (~(HRDATAS[8] & Ad47x6));
assign Cvnhy6 = (~(HRDATAD[8] & Mc47x6));
assign Ghmhy6 = (~(Lpryx6 & Kqonv6));
assign Foo7v6 = (~(Svnhy6 & Awnhy6));
assign Awnhy6 = (~(Jexmz6[9] & K94iw6));
assign Svnhy6 = (Iwnhy6 & Qwnhy6);
assign Qwnhy6 = (~(Lloyx6 & Ab67x6));
assign Ab67x6 = (~(Ywnhy6 & Gxnhy6));
assign Gxnhy6 = (Oxnhy6 & Wxnhy6);
assign Wxnhy6 = (Bqoyx6 | Kme7x6);
assign Kme7x6 = (Eynhy6 & Mynhy6);
assign Mynhy6 = (Uynhy6 & Cznhy6);
assign Cznhy6 = (Kznhy6 & Sznhy6);
assign Sznhy6 = (~(Rmzyx6 & A0ohy6));
assign A0ohy6 = (~(I0ohy6 & Q0ohy6));
assign Q0ohy6 = (Y0ohy6 & G1ohy6);
assign G1ohy6 = (O1ohy6 & W1ohy6);
assign W1ohy6 = (~(Hyj7z6[3] & Sybiw6));
assign O1ohy6 = (~(Hyj7z6[2] & Lybiw6));
assign Y0ohy6 = (E2ohy6 & M2ohy6);
assign M2ohy6 = (~(Hyj7z6[1] & Eybiw6));
assign E2ohy6 = (~(Hyj7z6[5] & Zybiw6));
assign I0ohy6 = (U2ohy6 & C3ohy6);
assign C3ohy6 = (K3ohy6 & S3ohy6);
assign S3ohy6 = (~(Hyj7z6[6] & Gzbiw6));
assign K3ohy6 = (~(Hyj7z6[7] & Nzbiw6));
assign U2ohy6 = (A4ohy6 & I4ohy6);
assign I4ohy6 = (~(Hyj7z6[0] & Dfk7z6[9]));
assign A4ohy6 = (~(Hyj7z6[4] & Jkl7z6[9]));
assign Kznhy6 = (Q4ohy6 & Y4ohy6);
assign Y4ohy6 = (~(D1pyx6 & G5ohy6));
assign G5ohy6 = (~(O5ohy6 & W5ohy6));
assign W5ohy6 = (E6ohy6 & Z6yyx6);
assign E6ohy6 = (~(M6ohy6 & C5rnv6));
assign M6ohy6 = (Unymz6[4] & Thpyx6);
assign O5ohy6 = (U6ohy6 & C7ohy6);
assign C7ohy6 = (~(Blsnv6 & Ngpyx6));
assign U6ohy6 = (~(Hl4xx6 & Hfpyx6));
assign Q4ohy6 = (~(Klo7z6[3] & K7ohy6));
assign K7ohy6 = (~(S7ohy6 & A8ohy6));
assign A8ohy6 = (~(W177v6 & Iknhy6));
assign S7ohy6 = (I8ohy6 & Q8ohy6);
assign Q8ohy6 = (~(Pk1nz6[9] & A8jhy6));
assign I8ohy6 = (~(Biymz6[9] & Olnhy6));
assign Uynhy6 = (Y8ohy6 & G9ohy6);
assign G9ohy6 = (~(Klo7z6[1] & O9ohy6));
assign O9ohy6 = (~(W9ohy6 & Eaohy6));
assign Eaohy6 = (Maohy6 & Uaohy6);
assign Uaohy6 = (Cbohy6 & Kbohy6);
assign Kbohy6 = (~(T9tyx6 & Ot77z6));
assign Cbohy6 = (Ravyx6 & Sbohy6);
assign Sbohy6 = (!Q0a8x6);
assign Maohy6 = (Acohy6 & Icohy6);
assign Icohy6 = (~(Id4ft6 & B6qyx6));
assign Acohy6 = (~(D5qyx6 & Bqp7z6[9]));
assign W9ohy6 = (Qcohy6 & Ycohy6);
assign Ycohy6 = (Gdohy6 & Odohy6);
assign Odohy6 = (~(L9qyx6 & E6p7z6[9]));
assign Gdohy6 = (~(Fcqyx6 & B2q7z6[9]));
assign Qcohy6 = (Wdohy6 & Eeohy6);
assign Eeohy6 = (~(Tdqyx6 & Mkp7z6[9]));
assign Wdohy6 = (~(U9p7z6[9] & Hfqyx6));
assign Y8ohy6 = (Meohy6 & Ueohy6);
assign Ueohy6 = (~(Xbzyx6 & Cfohy6));
assign Cfohy6 = (~(Kfohy6 & Sfohy6));
assign Sfohy6 = (Agohy6 & Igohy6);
assign Igohy6 = (Qgohy6 & Ygohy6);
assign Ygohy6 = (~(Hyj7z6[0] & Rbk7z6[7]));
assign Qgohy6 = (~(Hyj7z6[1] & Zlk7z6[7]));
assign Agohy6 = (Ghohy6 & Ohohy6);
assign Ohohy6 = (~(Hyj7z6[2] & Hwk7z6[7]));
assign Ghohy6 = (~(Hyj7z6[3] & P6l7z6[7]));
assign Kfohy6 = (Whohy6 & Eiohy6);
assign Eiohy6 = (Miohy6 & Uiohy6);
assign Uiohy6 = (~(Hyj7z6[4] & Xgl7z6[7]));
assign Miohy6 = (~(Hyj7z6[5] & Frl7z6[7]));
assign Whohy6 = (Cjohy6 & Kjohy6);
assign Kjohy6 = (~(Hyj7z6[6] & N1m7z6[7]));
assign Cjohy6 = (~(Hyj7z6[7] & Vbm7z6[7]));
assign Meohy6 = (~(Sjohy6 & Ngqyx6));
assign Sjohy6 = (~(Akohy6 & Ikohy6));
assign Ikohy6 = (Qkohy6 & Ykohy6);
assign Ykohy6 = (Glohy6 & Olohy6);
assign Olohy6 = (Wlohy6 & Emohy6);
assign Emohy6 = (~(A0j7z6[9] & Xrqyx6));
assign Wlohy6 = (Mmohy6 & Umohy6);
assign Umohy6 = (~(Cnohy6 & Fs0zx6));
assign Cnohy6 = (Lpyyx6 & Tpyyx6);
assign Mmohy6 = (~(Dtadt6 & Hnqyx6));
assign Hnqyx6 = (~(Tlqyx6 | Knohy6));
assign Glohy6 = (Snohy6 & Aoohy6);
assign Aoohy6 = (~(H1j7z6[9] & Rqqyx6));
assign Snohy6 = (~(X0eet6 & Ttqyx6));
assign Qkohy6 = (Ioohy6 & Qoohy6);
assign Qoohy6 = (Yoohy6 & Gpohy6);
assign Gpohy6 = (~(Dri7z6[9] & Fwqyx6));
assign Yoohy6 = (Opohy6 & Wpohy6);
assign Wpohy6 = (~(Bzi7z6[9] & Vsqyx6));
assign Opohy6 = (~(Wui7z6[9] & Lxqyx6));
assign Ioohy6 = (Eqohy6 & Mqohy6);
assign Mqohy6 = (~(Bwi7z6[9] & Hzqyx6));
assign Eqohy6 = (~(Svkhy6 & Qti7z6[9]));
assign Akohy6 = (Uqohy6 & Crohy6);
assign Crohy6 = (Krohy6 & Srohy6);
assign Srohy6 = (Asohy6 & Isohy6);
assign Isohy6 = (~(B2ryx6 & M6j7z6[41]));
assign Asohy6 = (Qsohy6 & Ysohy6);
assign Ysohy6 = (~(Pzqyx6 & G5j7z6[41]));
assign Qsohy6 = (~(Jyqyx6 & G5j7z6[9]));
assign Krohy6 = (Gtohy6 & Otohy6);
assign Otohy6 = (~(J2ryx6 & M6j7z6[9]));
assign Gtohy6 = (~(D1ryx6 & Ohj7z6[41]));
assign Uqohy6 = (Wtohy6 & Euohy6);
assign Euohy6 = (Muohy6 & Uuohy6);
assign Uuohy6 = (~(O5nhy6 & Hsi7z6[1]));
assign Muohy6 = (~(X3ryx6 & Ohj7z6[9]));
assign Wtohy6 = (Z2ryx6 & Cvohy6);
assign Cvohy6 = (~(STCALIB[9] & F4ryx6));
assign Eynhy6 = (Kvohy6 & Svohy6);
assign Svohy6 = (Awohy6 & Iwohy6);
assign Iwohy6 = (~(Zs1nz6[1] & Xjtyx6));
assign Awohy6 = (Qwohy6 & Ywohy6);
assign Ywohy6 = (~(Klo7z6[2] & Gxohy6));
assign Gxohy6 = (~(Oxohy6 & Wxohy6));
assign Wxohy6 = (Eyohy6 & Myohy6);
assign Myohy6 = (Uyohy6 & Czohy6);
assign Czohy6 = (~(Fpo7z6[7] & H9kiw6));
assign Uyohy6 = (Kzohy6 & S7khy6);
assign S7khy6 = (!Q3kiw6);
assign Q3kiw6 = (Szohy6 & A0phy6);
assign Szohy6 = (Hfuyx6 & Uamhy6);
assign Kzohy6 = (~(Nqo7z6[7] & M8kiw6));
assign Eyohy6 = (I0phy6 & Q0phy6);
assign Q0phy6 = (~(Ratet6 & S4kiw6));
assign I0phy6 = (~(Ouo7z6[7] & K7kiw6));
assign Oxohy6 = (Y0phy6 & G1phy6);
assign G1phy6 = (O1phy6 & W1phy6);
assign W1phy6 = (~(T2p7z6[9] & U5kiw6));
assign O1phy6 = (E2phy6 & M2phy6);
assign M2phy6 = (~(Hxo7z6[7] & W6kiw6));
assign E2phy6 = (~(Vro7z6[7] & Y7kiw6));
assign Y0phy6 = (U2phy6 & C3phy6);
assign C3phy6 = (~(W3p7z6[9] & G5kiw6));
assign U2phy6 = (~(A0p7z6[7] & I6kiw6));
assign Qwohy6 = (~(Nn1nz6[1] & Pjtyx6));
assign Kvohy6 = (K3phy6 & S3phy6);
assign S3phy6 = (~(Zm37v6 & Lltyx6));
assign K3phy6 = (~(Ies7z6[9] & Tltyx6));
assign Oxnhy6 = (~(Zmoyx6 & Rme7x6));
assign Rme7x6 = (~(A4phy6 & I4phy6));
assign I4phy6 = (~(Ysnhy6 & Ica7z6));
assign Ica7z6 = (~(Q4phy6 & Y4phy6));
assign Y4phy6 = (~(HRDATAD[9] & Qln7z6[0]));
assign Q4phy6 = (~(HRDATAS[9] & Qln7z6[1]));
assign A4phy6 = (~(Tim7z6[9] & Uunhy6));
assign Ywnhy6 = (G5phy6 & O5phy6);
assign O5phy6 = (~(HRDATAS[9] & Ad47x6));
assign G5phy6 = (~(HRDATAD[9] & Mc47x6));
assign Iwnhy6 = (~(Lpryx6 & H5q7x6));
assign Yno7v6 = (~(W5phy6 & E6phy6));
assign E6phy6 = (~(Jexmz6[10] & K94iw6));
assign W5phy6 = (M6phy6 & U6phy6);
assign U6phy6 = (~(Lloyx6 & Kdfov6));
assign Kdfov6 = (~(C7phy6 & K7phy6));
assign K7phy6 = (S7phy6 & A8phy6);
assign A8phy6 = (Bqoyx6 | Xpe7x6);
assign Xpe7x6 = (I8phy6 & Q8phy6);
assign Q8phy6 = (Y8phy6 & G9phy6);
assign G9phy6 = (O9phy6 & W9phy6);
assign W9phy6 = (~(Rmzyx6 & Eaphy6));
assign Eaphy6 = (~(Maphy6 & Uaphy6));
assign Uaphy6 = (Cbphy6 & Kbphy6);
assign Kbphy6 = (Sbphy6 & Acphy6);
assign Acphy6 = (~(Hyj7z6[3] & I0ciw6));
assign Sbphy6 = (~(Hyj7z6[2] & B0ciw6));
assign Cbphy6 = (Icphy6 & Qcphy6);
assign Qcphy6 = (~(Hyj7z6[1] & Uzbiw6));
assign Icphy6 = (~(Hyj7z6[5] & P0ciw6));
assign Maphy6 = (Ycphy6 & Gdphy6);
assign Gdphy6 = (Odphy6 & Wdphy6);
assign Wdphy6 = (~(Hyj7z6[6] & W0ciw6));
assign Odphy6 = (~(Hyj7z6[7] & D1ciw6));
assign Ycphy6 = (Eephy6 & Mephy6);
assign Mephy6 = (~(Hyj7z6[0] & Dfk7z6[10]));
assign Eephy6 = (~(Hyj7z6[4] & Jkl7z6[10]));
assign O9phy6 = (~(Xbzyx6 & Uephy6));
assign Uephy6 = (~(Cfphy6 & Kfphy6));
assign Kfphy6 = (Sfphy6 & Agphy6);
assign Agphy6 = (Igphy6 & Qgphy6);
assign Qgphy6 = (~(Hyj7z6[0] & Rbk7z6[8]));
assign Igphy6 = (~(Hyj7z6[1] & Zlk7z6[8]));
assign Sfphy6 = (Ygphy6 & Ghphy6);
assign Ghphy6 = (~(Hyj7z6[2] & Hwk7z6[8]));
assign Ygphy6 = (~(Hyj7z6[3] & P6l7z6[8]));
assign Cfphy6 = (Ohphy6 & Whphy6);
assign Whphy6 = (Eiphy6 & Miphy6);
assign Miphy6 = (~(Hyj7z6[4] & Xgl7z6[8]));
assign Eiphy6 = (~(Hyj7z6[5] & Frl7z6[8]));
assign Ohphy6 = (Uiphy6 & Cjphy6);
assign Cjphy6 = (~(Hyj7z6[6] & N1m7z6[8]));
assign Uiphy6 = (~(Hyj7z6[7] & Vbm7z6[8]));
assign Y8phy6 = (Kjphy6 & Sjphy6);
assign Sjphy6 = (~(Akphy6 & Ngqyx6));
assign Akphy6 = (~(Ikphy6 & Qkphy6));
assign Qkphy6 = (Ykphy6 & Glphy6);
assign Glphy6 = (Olphy6 & Wlphy6);
assign Wlphy6 = (Emphy6 & Mmphy6);
assign Mmphy6 = (~(H1j7z6[10] & Rqqyx6));
assign Emphy6 = (Umphy6 & Cnphy6);
assign Cnphy6 = (~(Prqyx6 & Z3j7z6[10]));
assign Umphy6 = (~(A0j7z6[10] & Xrqyx6));
assign Olphy6 = (Knphy6 & Snphy6);
assign Snphy6 = (~(W2eet6 & Ttqyx6));
assign Knphy6 = (~(Bzi7z6[10] & Vsqyx6));
assign Ykphy6 = (Aophy6 & Iophy6);
assign Iophy6 = (Qophy6 & Yophy6);
assign Yophy6 = (~(Wui7z6[10] & Lxqyx6));
assign Qophy6 = (~(Dri7z6[10] & Fwqyx6));
assign Aophy6 = (Gpphy6 & Opphy6);
assign Opphy6 = (~(Bwi7z6[10] & Hzqyx6));
assign Gpphy6 = (~(Svkhy6 & Pnb7z6[10]));
assign Ikphy6 = (Wpphy6 & Eqphy6);
assign Eqphy6 = (Mqphy6 & Uqphy6);
assign Uqphy6 = (Crphy6 & Krphy6);
assign Krphy6 = (~(Pzqyx6 & G5j7z6[42]));
assign Crphy6 = (~(Jyqyx6 & G5j7z6[10]));
assign Mqphy6 = (Srphy6 & Asphy6);
assign Asphy6 = (~(B2ryx6 & M6j7z6[42]));
assign Srphy6 = (~(J2ryx6 & M6j7z6[10]));
assign Wpphy6 = (Isphy6 & Qsphy6);
assign Qsphy6 = (Ysphy6 & Gtphy6);
assign Gtphy6 = (~(D1ryx6 & Ohj7z6[42]));
assign Ysphy6 = (~(Hsi7z6[2] & O5nhy6));
assign Isphy6 = (Otphy6 & Wtphy6);
assign Wtphy6 = (~(X3ryx6 & Ohj7z6[10]));
assign Otphy6 = (~(STCALIB[10] & F4ryx6));
assign Kjphy6 = (~(Klo7z6[1] & Euphy6));
assign Euphy6 = (~(Muphy6 & Uuphy6));
assign Uuphy6 = (Cvphy6 & Kvphy6);
assign Kvphy6 = (Svphy6 & Awphy6);
assign Awphy6 = (~(W5q7z6[0] & B6qyx6));
assign Svphy6 = (Iwphy6 & Ravyx6);
assign Iwphy6 = (~(T9tyx6 & Gt77z6));
assign Cvphy6 = (Qwphy6 & Ywphy6);
assign Ywphy6 = (~(D5qyx6 & Bqp7z6[10]));
assign Qwphy6 = (~(L9qyx6 & E6p7z6[10]));
assign Muphy6 = (Gxphy6 & Oxphy6);
assign Oxphy6 = (Wxphy6 & Eyphy6);
assign Eyphy6 = (~(Fcqyx6 & B2q7z6[10]));
assign Wxphy6 = (~(Gwp7z6[0] & Q0a8x6));
assign Gxphy6 = (Myphy6 & Uyphy6);
assign Uyphy6 = (~(Tdqyx6 & Mkp7z6[10]));
assign Myphy6 = (~(U9p7z6[10] & Hfqyx6));
assign I8phy6 = (Czphy6 & Kzphy6);
assign Kzphy6 = (Szphy6 & A0qhy6);
assign A0qhy6 = (~(Klo7z6[3] & I0qhy6));
assign I0qhy6 = (~(Q0qhy6 & Y0qhy6));
assign Y0qhy6 = (G1qhy6 & O1qhy6);
assign O1qhy6 = (W1qhy6 & E2qhy6);
assign E2qhy6 = (~(Blsnv6 & Glnhy6));
assign W1qhy6 = (M2qhy6 & U2qhy6);
assign M2qhy6 = (~(Mphiw6 & C3qhy6));
assign C3qhy6 = (~(K3qhy6 & S3qhy6));
assign S3qhy6 = (~(A4qhy6 & I4qhy6));
assign I4qhy6 = (Q4qhy6 & Y4qhy6);
assign Y4qhy6 = (~(Feymz6[2] | Feymz6[3]));
assign Q4qhy6 = (~(Bfymz6[2] | Feymz6[1]));
assign A4qhy6 = (G5qhy6 & O5qhy6);
assign O5qhy6 = (~(Bfymz6[0] | Bfymz6[1]));
assign G5qhy6 = (Feymz6[0] & Ignhy6);
assign Ignhy6 = (!L5pyx6);
assign K3qhy6 = (~(D9pyx6 & W5qhy6));
assign G1qhy6 = (E6qhy6 & M6qhy6);
assign M6qhy6 = (~(Hl4xx6 & Minhy6));
assign Q0qhy6 = (U6qhy6 & C7qhy6);
assign C7qhy6 = (K7qhy6 & S7qhy6);
assign S7qhy6 = (~(C477v6 & Iknhy6));
assign K7qhy6 = (A8qhy6 & I8qhy6);
assign I8qhy6 = (~(Pk1nz6[10] & A8jhy6));
assign A8qhy6 = (~(Biymz6[10] & Olnhy6));
assign U6qhy6 = (Q8qhy6 & Y8qhy6);
assign Y8qhy6 = (~(Zs1nz6[2] & S3mhy6));
assign Q8qhy6 = (~(Nn1nz6[2] & U2mhy6));
assign Szphy6 = (~(Klo7z6[2] & G9qhy6));
assign G9qhy6 = (~(O9qhy6 & W9qhy6));
assign W9qhy6 = (Eaqhy6 & Maqhy6);
assign Maqhy6 = (Uaqhy6 & Cbqhy6);
assign Cbqhy6 = (~(Q8tet6 & S4kiw6));
assign Uaqhy6 = (Kbqhy6 & Sbqhy6);
assign Sbqhy6 = (~(Nqo7z6[8] & M8kiw6));
assign Kbqhy6 = (~(Fpo7z6[8] & H9kiw6));
assign Eaqhy6 = (Acqhy6 & Icqhy6);
assign Icqhy6 = (~(Ouo7z6[8] & K7kiw6));
assign Acqhy6 = (~(Hxo7z6[8] & W6kiw6));
assign O9qhy6 = (Qcqhy6 & Ycqhy6);
assign Ycqhy6 = (Gdqhy6 & Odqhy6);
assign Odqhy6 = (~(Vro7z6[8] & Y7kiw6));
assign Gdqhy6 = (~(T2p7z6[10] & U5kiw6));
assign Qcqhy6 = (Wdqhy6 & Eeqhy6);
assign Eeqhy6 = (~(W3p7z6[10] & G5kiw6));
assign Wdqhy6 = (~(A0p7z6[8] & I6kiw6));
assign Czphy6 = (Meqhy6 & Ueqhy6);
assign Ueqhy6 = (~(Lltyx6 & R8s7z6[0]));
assign Meqhy6 = (~(Ies7z6[10] & Tltyx6));
assign S7phy6 = (~(Zmoyx6 & Eqe7x6));
assign Eqe7x6 = (~(Cfqhy6 & Kfqhy6));
assign Kfqhy6 = (~(Ysnhy6 & Aca7z6));
assign Aca7z6 = (~(Sfqhy6 & Agqhy6));
assign Agqhy6 = (~(HRDATAD[10] & Qln7z6[0]));
assign Sfqhy6 = (~(HRDATAS[10] & Qln7z6[1]));
assign Cfqhy6 = (~(Tim7z6[10] & Uunhy6));
assign C7phy6 = (Igqhy6 & Qgqhy6);
assign Qgqhy6 = (~(HRDATAS[10] & Ad47x6));
assign Igqhy6 = (~(HRDATAD[10] & Mc47x6));
assign M6phy6 = (~(Lpryx6 & Raq7x6));
assign Rno7v6 = (~(Ygqhy6 & Ghqhy6));
assign Ghqhy6 = (~(Jexmz6[11] & K94iw6));
assign Ygqhy6 = (Ohqhy6 & Whqhy6);
assign Whqhy6 = (~(Lloyx6 & Onlov6));
assign Onlov6 = (~(Eiqhy6 & Miqhy6));
assign Miqhy6 = (Uiqhy6 & Cjqhy6);
assign Cjqhy6 = (Bqoyx6 | Kte7x6);
assign Kte7x6 = (Kjqhy6 & Sjqhy6);
assign Sjqhy6 = (Akqhy6 & Ikqhy6);
assign Ikqhy6 = (Qkqhy6 & Ykqhy6);
assign Ykqhy6 = (~(Rmzyx6 & Glqhy6));
assign Glqhy6 = (~(Olqhy6 & Wlqhy6));
assign Wlqhy6 = (Emqhy6 & Mmqhy6);
assign Mmqhy6 = (Umqhy6 & Cnqhy6);
assign Cnqhy6 = (~(Hyj7z6[3] & A3ciw6));
assign Umqhy6 = (~(Hyj7z6[2] & M2ciw6));
assign Emqhy6 = (Knqhy6 & Snqhy6);
assign Snqhy6 = (~(Hyj7z6[1] & Y1ciw6));
assign Knqhy6 = (~(Hyj7z6[5] & V3ciw6));
assign Olqhy6 = (Aoqhy6 & Ioqhy6);
assign Ioqhy6 = (Qoqhy6 & Yoqhy6);
assign Yoqhy6 = (~(Hyj7z6[6] & Q4ciw6));
assign Qoqhy6 = (~(Hyj7z6[7] & X4ciw6));
assign Aoqhy6 = (Gpqhy6 & Opqhy6);
assign Opqhy6 = (~(Hyj7z6[0] & Dfk7z6[11]));
assign Gpqhy6 = (~(Hyj7z6[4] & Jkl7z6[11]));
assign Qkqhy6 = (Wpqhy6 & Eqqhy6);
assign Eqqhy6 = (~(Mqqhy6 & Uqqhy6));
assign Uqqhy6 = (~(Dtj7z6[2] | Dtj7z6[3]));
assign Mqqhy6 = (X7uyx6 & Dtj7z6[4]);
assign X7uyx6 = (Crqhy6 & Rmget6);
assign Crqhy6 = (Klo7z6[5] & T59iw6);
assign Wpqhy6 = (~(Xbzyx6 & Krqhy6));
assign Krqhy6 = (~(Srqhy6 & Asqhy6));
assign Asqhy6 = (Isqhy6 & Qsqhy6);
assign Qsqhy6 = (Ysqhy6 & Gtqhy6);
assign Gtqhy6 = (~(Hyj7z6[0] & Rbk7z6[9]));
assign Ysqhy6 = (~(Hyj7z6[1] & Zlk7z6[9]));
assign Isqhy6 = (Otqhy6 & Wtqhy6);
assign Wtqhy6 = (~(Hyj7z6[2] & Hwk7z6[9]));
assign Otqhy6 = (~(Hyj7z6[3] & P6l7z6[9]));
assign Srqhy6 = (Euqhy6 & Muqhy6);
assign Muqhy6 = (Uuqhy6 & Cvqhy6);
assign Cvqhy6 = (~(Hyj7z6[4] & Xgl7z6[9]));
assign Uuqhy6 = (~(Hyj7z6[5] & Frl7z6[9]));
assign Euqhy6 = (Kvqhy6 & Svqhy6);
assign Svqhy6 = (~(Hyj7z6[6] & N1m7z6[9]));
assign Kvqhy6 = (~(Hyj7z6[7] & Vbm7z6[9]));
assign Akqhy6 = (Awqhy6 & Iwqhy6);
assign Iwqhy6 = (~(Qwqhy6 & Ngqyx6));
assign Qwqhy6 = (~(Ywqhy6 & Gxqhy6));
assign Gxqhy6 = (Oxqhy6 & Wxqhy6);
assign Wxqhy6 = (Eyqhy6 & Myqhy6);
assign Myqhy6 = (Uyqhy6 & Czqhy6);
assign Czqhy6 = (~(Prqyx6 & Z3j7z6[11]));
assign Uyqhy6 = (~(A0j7z6[11] & Xrqyx6));
assign Eyqhy6 = (Kzqhy6 & Szqhy6);
assign Szqhy6 = (~(H1j7z6[11] & Rqqyx6));
assign Kzqhy6 = (~(Bzi7z6[11] & Vsqyx6));
assign Oxqhy6 = (A0rhy6 & I0rhy6);
assign I0rhy6 = (Q0rhy6 & Y0rhy6);
assign Y0rhy6 = (~(Wbcet6 & Dxqyx6));
assign Q0rhy6 = (~(Wui7z6[11] & Lxqyx6));
assign A0rhy6 = (G1rhy6 & O1rhy6);
assign O1rhy6 = (~(Dri7z6[11] & Fwqyx6));
assign G1rhy6 = (~(Bwi7z6[11] & Hzqyx6));
assign Ywqhy6 = (W1rhy6 & E2rhy6);
assign E2rhy6 = (M2rhy6 & U2rhy6);
assign U2rhy6 = (C3rhy6 & K3rhy6);
assign K3rhy6 = (~(Svkhy6 & Pnb7z6[11]));
assign C3rhy6 = (~(Pzqyx6 & G5j7z6[43]));
assign M2rhy6 = (S3rhy6 & A4rhy6);
assign A4rhy6 = (~(Jyqyx6 & G5j7z6[11]));
assign S3rhy6 = (~(B2ryx6 & M6j7z6[43]));
assign W1rhy6 = (I4rhy6 & Q4rhy6);
assign Q4rhy6 = (Y4rhy6 & G5rhy6);
assign G5rhy6 = (~(J2ryx6 & M6j7z6[11]));
assign Y4rhy6 = (~(D1ryx6 & Ohj7z6[43]));
assign I4rhy6 = (O5rhy6 & W5rhy6);
assign W5rhy6 = (~(X3ryx6 & Ohj7z6[11]));
assign O5rhy6 = (~(STCALIB[11] & F4ryx6));
assign Awqhy6 = (~(Klo7z6[3] & E6rhy6));
assign E6rhy6 = (~(M6rhy6 & U6rhy6));
assign U6rhy6 = (C7rhy6 & K7rhy6);
assign K7rhy6 = (S7rhy6 & A8rhy6);
assign A8rhy6 = (~(Mphiw6 & I8rhy6));
assign I8rhy6 = (~(Q8rhy6 & Y8rhy6));
assign Y8rhy6 = (~(G9rhy6 & O9rhy6));
assign O9rhy6 = (~(Bfymz6[1] | Bfymz6[2]));
assign G9rhy6 = (~(L5pyx6 | Bfymz6[0]));
assign S7rhy6 = (W9rhy6 & Earhy6);
assign Earhy6 = (~(Marhy6 & Blsnv6));
assign Blsnv6 = (Uarhy6 & Sgymz6[7]);
assign Uarhy6 = (Sgymz6[4] & Sgymz6[5]);
assign Marhy6 = (~(Cbrhy6 | Sgymz6[6]));
assign W9rhy6 = (~(Kbrhy6 & Hl4xx6));
assign Hl4xx6 = (Sbrhy6 & Ojymz6[7]);
assign Sbrhy6 = (Ojymz6[4] & Ojymz6[5]);
assign Kbrhy6 = (~(Acrhy6 | Ojymz6[6]));
assign C7rhy6 = (E6qhy6 & Icrhy6);
assign Icrhy6 = (U2qhy6 | Unymz6[6]);
assign U2qhy6 = (~(Qcrhy6 & C5rnv6));
assign C5rnv6 = (Unymz6[7] & Unymz6[5]);
assign Qcrhy6 = (Unymz6[4] & Uinhy6);
assign E6qhy6 = (Eylhy6 | Qgnhy6);
assign Eylhy6 = (~(Ycrhy6 & Gdrhy6));
assign Gdrhy6 = (Odrhy6 & Xvxyx6);
assign Odrhy6 = (J02nz6[8] & L9syx6);
assign Ycrhy6 = (Hrpyx6 & J02nz6[3]);
assign Hrpyx6 = (~(J02nz6[2] | J02nz6[4]));
assign M6rhy6 = (Wdrhy6 & Eerhy6);
assign Eerhy6 = (Merhy6 & Uerhy6);
assign Uerhy6 = (~(Ue77z6 & Iknhy6));
assign Merhy6 = (Cfrhy6 & Kfrhy6);
assign Kfrhy6 = (~(Pk1nz6[11] & A8jhy6));
assign Cfrhy6 = (~(Biymz6[11] & Olnhy6));
assign Wdrhy6 = (Sfrhy6 & Agrhy6);
assign Agrhy6 = (~(Zs1nz6[3] & S3mhy6));
assign Sfrhy6 = (~(Nn1nz6[3] & U2mhy6));
assign Kjqhy6 = (Igrhy6 & Qgrhy6);
assign Qgrhy6 = (Ygrhy6 & Ghrhy6);
assign Ghrhy6 = (~(Klo7z6[1] & Ohrhy6));
assign Ohrhy6 = (~(Whrhy6 & Eirhy6));
assign Eirhy6 = (Mirhy6 & Uirhy6);
assign Uirhy6 = (Cjrhy6 & Kjrhy6);
assign Kjrhy6 = (~(W5q7z6[1] & B6qyx6));
assign Cjrhy6 = (Sjrhy6 & Ravyx6);
assign Sjrhy6 = (~(T9tyx6 & Ys77z6));
assign Mirhy6 = (Akrhy6 & Ikrhy6);
assign Ikrhy6 = (~(D5qyx6 & Bqp7z6[11]));
assign Akrhy6 = (~(L9qyx6 & E6p7z6[11]));
assign Whrhy6 = (Qkrhy6 & Ykrhy6);
assign Ykrhy6 = (Glrhy6 & Olrhy6);
assign Olrhy6 = (~(Fcqyx6 & B2q7z6[11]));
assign Glrhy6 = (~(Gwp7z6[1] & Q0a8x6));
assign Qkrhy6 = (Wlrhy6 & Emrhy6);
assign Emrhy6 = (~(Tdqyx6 & Mkp7z6[11]));
assign Wlrhy6 = (~(U9p7z6[11] & Hfqyx6));
assign Ygrhy6 = (~(Klo7z6[2] & Mmrhy6));
assign Mmrhy6 = (~(Umrhy6 & Cnrhy6));
assign Cnrhy6 = (Knrhy6 & Snrhy6);
assign Snrhy6 = (Aorhy6 & Iorhy6);
assign Iorhy6 = (~(P6tet6 & S4kiw6));
assign Aorhy6 = (Qorhy6 & Yorhy6);
assign Yorhy6 = (~(Nqo7z6[9] & M8kiw6));
assign Qorhy6 = (~(Fpo7z6[9] & H9kiw6));
assign Knrhy6 = (Gprhy6 & Oprhy6);
assign Oprhy6 = (~(Ouo7z6[9] & K7kiw6));
assign Gprhy6 = (~(Hxo7z6[9] & W6kiw6));
assign Umrhy6 = (Wprhy6 & Eqrhy6);
assign Eqrhy6 = (Mqrhy6 & Uqrhy6);
assign Uqrhy6 = (~(Vro7z6[9] & Y7kiw6));
assign Mqrhy6 = (~(T2p7z6[11] & U5kiw6));
assign Wprhy6 = (Crrhy6 & Krrhy6);
assign Krrhy6 = (~(W3p7z6[11] & G5kiw6));
assign Crrhy6 = (~(A0p7z6[9] & I6kiw6));
assign Igrhy6 = (Srrhy6 & Asrhy6);
assign Asrhy6 = (~(R8s7z6[1] & Lltyx6));
assign Srrhy6 = (~(Ies7z6[11] & Tltyx6));
assign Uiqhy6 = (~(Zmoyx6 & Rte7x6));
assign Rte7x6 = (~(Isrhy6 & Qsrhy6));
assign Qsrhy6 = (~(Ysnhy6 & Sba7z6));
assign Sba7z6 = (~(Ysrhy6 & Gtrhy6));
assign Gtrhy6 = (~(HRDATAD[11] & Qln7z6[0]));
assign Ysrhy6 = (~(HRDATAS[11] & Qln7z6[1]));
assign Isrhy6 = (~(Tim7z6[11] & Uunhy6));
assign Eiqhy6 = (Otrhy6 & Wtrhy6);
assign Wtrhy6 = (~(HRDATAS[11] & Ad47x6));
assign Otrhy6 = (~(HRDATAD[11] & Mc47x6));
assign Ohqhy6 = (~(Lpryx6 & Bgq7x6));
assign Kno7v6 = (~(Eurhy6 & Murhy6));
assign Murhy6 = (~(Jexmz6[12] & K94iw6));
assign Eurhy6 = (Uurhy6 & Cvrhy6);
assign Cvrhy6 = (~(Lloyx6 & Tw57x6));
assign Tw57x6 = (~(Kvrhy6 & Svrhy6));
assign Svrhy6 = (Awrhy6 & Iwrhy6);
assign Iwrhy6 = (Bqoyx6 | Xwe7x6);
assign Xwe7x6 = (Qwrhy6 & Ywrhy6);
assign Ywrhy6 = (Gxrhy6 & Oxrhy6);
assign Oxrhy6 = (Wxrhy6 & Eyrhy6);
assign Eyrhy6 = (~(Rmzyx6 & Myrhy6));
assign Myrhy6 = (~(Uyrhy6 & Czrhy6));
assign Czrhy6 = (Kzrhy6 & Szrhy6);
assign Szrhy6 = (A0shy6 & I0shy6);
assign I0shy6 = (~(Hyj7z6[3] & N6ciw6));
assign A0shy6 = (~(Hyj7z6[2] & Z5ciw6));
assign Kzrhy6 = (Q0shy6 & Y0shy6);
assign Y0shy6 = (~(Hyj7z6[1] & L5ciw6));
assign Q0shy6 = (~(Hyj7z6[5] & I7ciw6));
assign Uyrhy6 = (G1shy6 & O1shy6);
assign O1shy6 = (W1shy6 & E2shy6);
assign E2shy6 = (~(Hyj7z6[6] & P7ciw6));
assign W1shy6 = (~(Hyj7z6[7] & D8ciw6));
assign G1shy6 = (M2shy6 & U2shy6);
assign U2shy6 = (~(Hyj7z6[0] & Dfk7z6[12]));
assign M2shy6 = (~(Hyj7z6[4] & Jkl7z6[12]));
assign Wxrhy6 = (~(Xbzyx6 & C3shy6));
assign C3shy6 = (~(K3shy6 & S3shy6));
assign S3shy6 = (A4shy6 & I4shy6);
assign I4shy6 = (Q4shy6 & Y4shy6);
assign Y4shy6 = (~(Hyj7z6[0] & Rbk7z6[10]));
assign Q4shy6 = (~(Hyj7z6[1] & Zlk7z6[10]));
assign A4shy6 = (G5shy6 & O5shy6);
assign O5shy6 = (~(Hyj7z6[2] & Hwk7z6[10]));
assign G5shy6 = (~(Hyj7z6[3] & P6l7z6[10]));
assign K3shy6 = (W5shy6 & E6shy6);
assign E6shy6 = (M6shy6 & U6shy6);
assign U6shy6 = (~(Hyj7z6[4] & Xgl7z6[10]));
assign M6shy6 = (~(Hyj7z6[5] & Frl7z6[10]));
assign W5shy6 = (C7shy6 & K7shy6);
assign K7shy6 = (~(Hyj7z6[6] & N1m7z6[10]));
assign C7shy6 = (~(Hyj7z6[7] & Vbm7z6[10]));
assign Gxrhy6 = (S7shy6 & A8shy6);
assign A8shy6 = (~(I8shy6 & Ngqyx6));
assign I8shy6 = (~(Q8shy6 & Y8shy6));
assign Y8shy6 = (G9shy6 & O9shy6);
assign O9shy6 = (W9shy6 & Eashy6);
assign Eashy6 = (Mashy6 & Uashy6);
assign Uashy6 = (~(H1j7z6[12] & Rqqyx6));
assign Mashy6 = (Cbshy6 & Kbshy6);
assign Kbshy6 = (~(Prqyx6 & Z3j7z6[12]));
assign Cbshy6 = (~(A0j7z6[12] & Xrqyx6));
assign W9shy6 = (Sbshy6 & Acshy6);
assign Acshy6 = (~(Bzi7z6[12] & Vsqyx6));
assign Sbshy6 = (~(Dxqyx6 & P2j7z6[0]));
assign G9shy6 = (Icshy6 & Qcshy6);
assign Qcshy6 = (Ycshy6 & Gdshy6);
assign Gdshy6 = (~(Wui7z6[12] & Lxqyx6));
assign Ycshy6 = (~(Dri7z6[12] & Fwqyx6));
assign Icshy6 = (Odshy6 & Wdshy6);
assign Wdshy6 = (~(Bwi7z6[12] & Hzqyx6));
assign Odshy6 = (~(Svkhy6 & Pnb7z6[12]));
assign Q8shy6 = (Eeshy6 & Meshy6);
assign Meshy6 = (Ueshy6 & Cfshy6);
assign Cfshy6 = (Kfshy6 & Sfshy6);
assign Sfshy6 = (~(Pzqyx6 & G5j7z6[44]));
assign Kfshy6 = (~(Jyqyx6 & G5j7z6[12]));
assign Ueshy6 = (Agshy6 & Igshy6);
assign Igshy6 = (~(B2ryx6 & M6j7z6[44]));
assign Agshy6 = (~(J2ryx6 & M6j7z6[12]));
assign Eeshy6 = (Qgshy6 & Ygshy6);
assign Ygshy6 = (Ghshy6 & Ohshy6);
assign Ohshy6 = (~(D1ryx6 & Ohj7z6[44]));
assign Ghshy6 = (~(X3ryx6 & Ohj7z6[12]));
assign Qgshy6 = (Whshy6 & Eishy6);
assign Eishy6 = (~(STCALIB[12] & F4ryx6));
assign S7shy6 = (~(Klo7z6[1] & Mishy6));
assign Mishy6 = (~(Uishy6 & Cjshy6));
assign Cjshy6 = (Kjshy6 & Sjshy6);
assign Sjshy6 = (Akshy6 & Ikshy6);
assign Ikshy6 = (~(Xkq7z6[12] & B6qyx6));
assign Akshy6 = (Qkshy6 & Ravyx6);
assign Qkshy6 = (~(T9tyx6 & Qs77z6));
assign Kjshy6 = (Ykshy6 & Glshy6);
assign Glshy6 = (~(D5qyx6 & Bqp7z6[12]));
assign Ykshy6 = (~(L9qyx6 & E6p7z6[12]));
assign Uishy6 = (Olshy6 & Wlshy6);
assign Wlshy6 = (Emshy6 & Mmshy6);
assign Mmshy6 = (~(Fcqyx6 & B2q7z6[12]));
assign Emshy6 = (~(Q0a8x6 & Bup7z6[0]));
assign Olshy6 = (Umshy6 & Cnshy6);
assign Cnshy6 = (~(Tdqyx6 & Mkp7z6[12]));
assign Umshy6 = (~(U9p7z6[12] & Hfqyx6));
assign Qwrhy6 = (Knshy6 & Snshy6);
assign Snshy6 = (~(Ies7z6[12] & Tltyx6));
assign Knshy6 = (Aoshy6 & Ioshy6);
assign Ioshy6 = (~(Klo7z6[3] & Qoshy6));
assign Qoshy6 = (~(Yoshy6 & Gpshy6));
assign Gpshy6 = (Opshy6 & Wpshy6);
assign Wpshy6 = (Eqshy6 & Mqshy6);
assign Mqshy6 = (~(Pk1nz6[12] & A8jhy6));
assign A8jhy6 = (Xvpyx6 & Kniiw6);
assign Xvpyx6 = (Yvhiw6 & Z2wyx6);
assign Z2wyx6 = (Iuhiw6 & Jke7v6);
assign Iuhiw6 = (Uqshy6 & Ohnhy6);
assign Ohnhy6 = (Crshy6 & Krshy6);
assign Krshy6 = (Srshy6 & L9syx6);
assign L9syx6 = (!J02nz6[5]);
assign Srshy6 = (~(J02nz6[6] | J02nz6[7]));
assign Crshy6 = (Asshy6 & H7syx6);
assign H7syx6 = (!J02nz6[10]);
assign Asshy6 = (~(J02nz6[11] | J02nz6[3]));
assign Uqshy6 = (~(J02nz6[8] | J02nz6[9]));
assign Yvhiw6 = (~(Puhiw6 | J02nz6[2]));
assign Eqshy6 = (Isshy6 & Qsshy6);
assign Qsshy6 = (~(Kzlhy6 & Ysshy6));
assign Ysshy6 = (~(Xntyx6 & Gtshy6));
assign Isshy6 = (Otshy6 | Wtshy6);
assign Opshy6 = (Eushy6 & Mushy6);
assign Mushy6 = (~(Ojymz6[6] & Minhy6));
assign Eushy6 = (~(Unymz6[6] & Uinhy6));
assign Yoshy6 = (Uushy6 & Cvshy6);
assign Cvshy6 = (Kvshy6 & Svshy6);
assign Svshy6 = (~(Sgymz6[6] & Glnhy6));
assign Kvshy6 = (~(Biymz6[12] & Olnhy6));
assign Uushy6 = (Awshy6 & Iwshy6);
assign Iwshy6 = (~(Zs1nz6[4] & S3mhy6));
assign Awshy6 = (~(Nn1nz6[4] & U2mhy6));
assign Aoshy6 = (~(Klo7z6[2] & Qwshy6));
assign Qwshy6 = (~(Ywshy6 & Gxshy6));
assign Gxshy6 = (Oxshy6 & Wxshy6);
assign Wxshy6 = (Eyshy6 & Myshy6);
assign Myshy6 = (~(O4tet6 & S4kiw6));
assign Eyshy6 = (Uyshy6 & Czshy6);
assign Czshy6 = (~(Nqo7z6[10] & M8kiw6));
assign Uyshy6 = (~(Fpo7z6[10] & H9kiw6));
assign Oxshy6 = (Kzshy6 & Szshy6);
assign Szshy6 = (~(Ouo7z6[10] & K7kiw6));
assign Kzshy6 = (~(Hxo7z6[10] & W6kiw6));
assign Ywshy6 = (A0thy6 & I0thy6);
assign I0thy6 = (Q0thy6 & Y0thy6);
assign Y0thy6 = (~(Vro7z6[10] & Y7kiw6));
assign Q0thy6 = (~(T2p7z6[12] & U5kiw6));
assign A0thy6 = (G1thy6 & O1thy6);
assign O1thy6 = (~(W3p7z6[12] & G5kiw6));
assign G1thy6 = (~(A0p7z6[10] & I6kiw6));
assign Awrhy6 = (~(Zmoyx6 & Exe7x6));
assign Exe7x6 = (~(W1thy6 & E2thy6));
assign E2thy6 = (~(Jco7v6 & Ysnhy6));
assign W1thy6 = (~(Tim7z6[12] & Uunhy6));
assign Kvrhy6 = (M2thy6 & U2thy6);
assign U2thy6 = (~(HRDATAS[12] & Ad47x6));
assign M2thy6 = (~(HRDATAD[12] & Mc47x6));
assign Uurhy6 = (~(Lpryx6 & Llq7x6));
assign Dno7v6 = (~(C3thy6 & K3thy6));
assign K3thy6 = (~(Jexmz6[13] & K94iw6));
assign C3thy6 = (S3thy6 & A4thy6);
assign A4thy6 = (~(Lloyx6 & Qr57x6));
assign Qr57x6 = (~(I4thy6 & Q4thy6));
assign Q4thy6 = (Y4thy6 & G5thy6);
assign G5thy6 = (Bqoyx6 | K0f7x6);
assign K0f7x6 = (O5thy6 & W5thy6);
assign W5thy6 = (E6thy6 & M6thy6);
assign M6thy6 = (U6thy6 & C7thy6);
assign C7thy6 = (~(Rmzyx6 & K7thy6));
assign K7thy6 = (~(S7thy6 & A8thy6));
assign A8thy6 = (I8thy6 & Q8thy6);
assign Q8thy6 = (Y8thy6 & G9thy6);
assign G9thy6 = (~(Hyj7z6[3] & Y8ciw6));
assign Y8thy6 = (~(Hyj7z6[2] & R8ciw6));
assign I8thy6 = (O9thy6 & W9thy6);
assign W9thy6 = (~(Hyj7z6[1] & K8ciw6));
assign O9thy6 = (~(Hyj7z6[5] & F9ciw6));
assign S7thy6 = (Eathy6 & Mathy6);
assign Mathy6 = (Uathy6 & Cbthy6);
assign Cbthy6 = (~(Hyj7z6[6] & M9ciw6));
assign Uathy6 = (~(Hyj7z6[7] & T9ciw6));
assign Eathy6 = (Kbthy6 & Sbthy6);
assign Sbthy6 = (~(Hyj7z6[0] & Dfk7z6[13]));
assign Kbthy6 = (~(Hyj7z6[4] & Jkl7z6[13]));
assign U6thy6 = (~(Xbzyx6 & Acthy6));
assign Acthy6 = (~(Icthy6 & Qcthy6));
assign Qcthy6 = (Ycthy6 & Gdthy6);
assign Gdthy6 = (Odthy6 & Wdthy6);
assign Wdthy6 = (~(Hyj7z6[0] & Rbk7z6[11]));
assign Odthy6 = (~(Hyj7z6[1] & Zlk7z6[11]));
assign Ycthy6 = (Eethy6 & Methy6);
assign Methy6 = (~(Hyj7z6[2] & Hwk7z6[11]));
assign Eethy6 = (~(Hyj7z6[3] & P6l7z6[11]));
assign Icthy6 = (Uethy6 & Cfthy6);
assign Cfthy6 = (Kfthy6 & Sfthy6);
assign Sfthy6 = (~(Hyj7z6[4] & Xgl7z6[11]));
assign Kfthy6 = (~(Hyj7z6[5] & Frl7z6[11]));
assign Uethy6 = (Agthy6 & Igthy6);
assign Igthy6 = (~(Hyj7z6[6] & N1m7z6[11]));
assign Agthy6 = (~(Hyj7z6[7] & Vbm7z6[11]));
assign E6thy6 = (Qgthy6 & Ygthy6);
assign Ygthy6 = (~(Ghthy6 & Ngqyx6));
assign Ghthy6 = (~(Ohthy6 & Whthy6));
assign Whthy6 = (Eithy6 & Mithy6);
assign Mithy6 = (Uithy6 & Cjthy6);
assign Cjthy6 = (Kjthy6 & Sjthy6);
assign Sjthy6 = (Akthy6 & Ikthy6);
assign Ikthy6 = (~(V40zx6 & Zdj7z6[0]));
assign Akthy6 = (Qkthy6 & Ykthy6);
assign Qkthy6 = (~(Prqyx6 & Z3j7z6[13]));
assign Kjthy6 = (Glthy6 & Olthy6);
assign Olthy6 = (~(A0j7z6[13] & Xrqyx6));
assign Glthy6 = (~(H1j7z6[13] & Rqqyx6));
assign Uithy6 = (Wlthy6 & Emthy6);
assign Emthy6 = (Mmthy6 & 1'b1);
assign Mmthy6 = (~(Dxqyx6 & P2j7z6[1]));
assign Wlthy6 = (Umthy6 & Cnthy6);
assign Cnthy6 = (~(Wui7z6[13] & Lxqyx6));
assign Umthy6 = (~(Dri7z6[13] & Fwqyx6));
assign Eithy6 = (Knthy6 & Snthy6);
assign Snthy6 = (Aothy6 & Iothy6);
assign Iothy6 = (Qothy6 & Yothy6);
assign Yothy6 = (~(Bwi7z6[13] & Hzqyx6));
assign Qothy6 = (~(Svkhy6 & Pnb7z6[13]));
assign Aothy6 = (Gpthy6 & Opthy6);
assign Opthy6 = (~(D90zx6 & Lgj7z6[183]));
assign Gpthy6 = (~(Za0zx6 & Lgj7z6[171]));
assign Knthy6 = (Wpthy6 & Eqthy6);
assign Eqthy6 = (Mqthy6 & Uqthy6);
assign Uqthy6 = (~(Hb0zx6 & Lgj7z6[159]));
assign Mqthy6 = (~(Vc0zx6 & Lgj7z6[147]));
assign Wpthy6 = (Crthy6 & Krthy6);
assign Krthy6 = (~(Dd0zx6 & Lgj7z6[135]));
assign Crthy6 = (~(Be0zx6 & Lgj7z6[123]));
assign Ohthy6 = (Srthy6 & Asthy6);
assign Asthy6 = (Isthy6 & Qsthy6);
assign Qsthy6 = (Ysthy6 & Gtthy6);
assign Gtthy6 = (Otthy6 & Wtthy6);
assign Wtthy6 = (~(Ji0zx6 & Lgj7z6[87]));
assign Otthy6 = (Euthy6 & Muthy6);
assign Muthy6 = (~(Je0zx6 & Lgj7z6[111]));
assign Euthy6 = (~(Bi0zx6 & Lgj7z6[99]));
assign Ysthy6 = (Uuthy6 & Cvthy6);
assign Cvthy6 = (~(Dh0zx6 & Lgj7z6[75]));
assign Uuthy6 = (~(Hj0zx6 & Lgj7z6[63]));
assign Isthy6 = (Kvthy6 & Svthy6);
assign Svthy6 = (Awthy6 & Iwthy6);
assign Iwthy6 = (~(Pj0zx6 & Lgj7z6[51]));
assign Awthy6 = (~(Dl0zx6 & Lgj7z6[39]));
assign Kvthy6 = (Qwthy6 & Ywthy6);
assign Ywthy6 = (~(Ll0zx6 & Lgj7z6[27]));
assign Qwthy6 = (~(Jm0zx6 & Lgj7z6[15]));
assign Srthy6 = (Gxthy6 & Oxthy6);
assign Oxthy6 = (Wxthy6 & Eythy6);
assign Eythy6 = (Mythy6 & Uythy6);
assign Uythy6 = (~(Rm0zx6 & Lgj7z6[3]));
assign Mythy6 = (~(Pzqyx6 & G5j7z6[45]));
assign Wxthy6 = (Czthy6 & Kzthy6);
assign Kzthy6 = (~(Jyqyx6 & G5j7z6[13]));
assign Czthy6 = (~(B2ryx6 & M6j7z6[45]));
assign Gxthy6 = (Szthy6 & A0uhy6);
assign A0uhy6 = (I0uhy6 & Q0uhy6);
assign Q0uhy6 = (~(J2ryx6 & M6j7z6[13]));
assign I0uhy6 = (~(D1ryx6 & Ohj7z6[45]));
assign Szthy6 = (Y0uhy6 & G1uhy6);
assign G1uhy6 = (~(X3ryx6 & Ohj7z6[13]));
assign Y0uhy6 = (~(STCALIB[13] & F4ryx6));
assign Qgthy6 = (~(Klo7z6[1] & O1uhy6));
assign O1uhy6 = (~(W1uhy6 & E2uhy6));
assign E2uhy6 = (M2uhy6 & U2uhy6);
assign U2uhy6 = (C3uhy6 & K3uhy6);
assign K3uhy6 = (~(Xkq7z6[13] & B6qyx6));
assign C3uhy6 = (S3uhy6 & Ravyx6);
assign S3uhy6 = (~(T9tyx6 & Is77z6));
assign M2uhy6 = (A4uhy6 & I4uhy6);
assign I4uhy6 = (~(D5qyx6 & Bqp7z6[13]));
assign A4uhy6 = (~(L9qyx6 & E6p7z6[13]));
assign W1uhy6 = (Q4uhy6 & Y4uhy6);
assign Y4uhy6 = (G5uhy6 & O5uhy6);
assign O5uhy6 = (~(Fcqyx6 & B2q7z6[13]));
assign G5uhy6 = (~(Q0a8x6 & Bup7z6[1]));
assign Q4uhy6 = (W5uhy6 & E6uhy6);
assign E6uhy6 = (~(Tdqyx6 & Mkp7z6[13]));
assign W5uhy6 = (~(U9p7z6[13] & Hfqyx6));
assign O5thy6 = (M6uhy6 & U6uhy6);
assign U6uhy6 = (~(Ies7z6[13] & Tltyx6));
assign M6uhy6 = (C7uhy6 & K7uhy6);
assign K7uhy6 = (~(Klo7z6[3] & S7uhy6));
assign S7uhy6 = (~(A8uhy6 & I8uhy6));
assign I8uhy6 = (Q8uhy6 & Y8uhy6);
assign Y8uhy6 = (G9uhy6 & O9uhy6);
assign O9uhy6 = (~(Unymz6[7] & Uinhy6));
assign G9uhy6 = (W9uhy6 & Eauhy6);
assign Eauhy6 = (~(Mphiw6 & Mauhy6));
assign Mauhy6 = (~(Z6yyx6 & Uauhy6));
assign Uauhy6 = (~(P3xyx6 & J2xyx6));
assign W9uhy6 = (~(Ojymz6[7] & Minhy6));
assign Q8uhy6 = (Cbuhy6 & Kbuhy6);
assign Kbuhy6 = (~(Sgymz6[7] & Glnhy6));
assign Cbuhy6 = (~(Biymz6[13] & Olnhy6));
assign A8uhy6 = (Sbuhy6 & Acuhy6);
assign Acuhy6 = (Icuhy6 & Qcuhy6);
assign Qcuhy6 = (~(Bfymz6[2] & Iknhy6));
assign Icuhy6 = (~(Zs1nz6[5] & S3mhy6));
assign Sbuhy6 = (Ycuhy6 & Gduhy6);
assign Gduhy6 = (~(Nn1nz6[5] & U2mhy6));
assign Ycuhy6 = (Oduhy6 | Pntyx6);
assign C7uhy6 = (~(Klo7z6[2] & Wduhy6));
assign Wduhy6 = (~(Eeuhy6 & Meuhy6));
assign Meuhy6 = (Ueuhy6 & Cfuhy6);
assign Cfuhy6 = (Kfuhy6 & Sfuhy6);
assign Sfuhy6 = (~(N2tet6 & S4kiw6));
assign Kfuhy6 = (Aguhy6 & Iguhy6);
assign Iguhy6 = (~(Nqo7z6[11] & M8kiw6));
assign Aguhy6 = (~(Fpo7z6[11] & H9kiw6));
assign Ueuhy6 = (Qguhy6 & Yguhy6);
assign Yguhy6 = (~(Ouo7z6[11] & K7kiw6));
assign Qguhy6 = (~(Hxo7z6[11] & W6kiw6));
assign Eeuhy6 = (Ghuhy6 & Ohuhy6);
assign Ohuhy6 = (Whuhy6 & Eiuhy6);
assign Eiuhy6 = (~(Vro7z6[11] & Y7kiw6));
assign Whuhy6 = (~(T2p7z6[13] & U5kiw6));
assign Ghuhy6 = (Miuhy6 & Uiuhy6);
assign Uiuhy6 = (~(W3p7z6[13] & G5kiw6));
assign Miuhy6 = (~(A0p7z6[11] & I6kiw6));
assign Y4thy6 = (~(Zmoyx6 & R0f7x6));
assign R0f7x6 = (~(Cjuhy6 & Kjuhy6));
assign Kjuhy6 = (~(Ysnhy6 & Kba7z6));
assign Kba7z6 = (~(Sjuhy6 & Akuhy6));
assign Akuhy6 = (~(HRDATAD[13] & Qln7z6[0]));
assign Sjuhy6 = (~(HRDATAS[13] & Qln7z6[1]));
assign Cjuhy6 = (~(Tim7z6[13] & Uunhy6));
assign I4thy6 = (Ikuhy6 & Qkuhy6);
assign Qkuhy6 = (~(HRDATAS[13] & Ad47x6));
assign Ikuhy6 = (~(HRDATAD[13] & Mc47x6));
assign S3thy6 = (~(Lpryx6 & Vqq7x6));
assign Wmo7v6 = (~(Ykuhy6 & Gluhy6));
assign Gluhy6 = (~(Jexmz6[14] & K94iw6));
assign Ykuhy6 = (Oluhy6 & Wluhy6);
assign Wluhy6 = (~(Lloyx6 & Nm57x6));
assign Nm57x6 = (~(Emuhy6 & Mmuhy6));
assign Mmuhy6 = (Umuhy6 & Cnuhy6);
assign Cnuhy6 = (Bqoyx6 | X3f7x6);
assign X3f7x6 = (Knuhy6 & Snuhy6);
assign Snuhy6 = (Aouhy6 & Iouhy6);
assign Iouhy6 = (Qouhy6 & Youhy6);
assign Youhy6 = (~(Rmzyx6 & Gpuhy6));
assign Gpuhy6 = (~(Opuhy6 & Wpuhy6));
assign Wpuhy6 = (Equhy6 & Mquhy6);
assign Mquhy6 = (Uquhy6 & Cruhy6);
assign Cruhy6 = (~(Hyj7z6[3] & Oaciw6));
assign Uquhy6 = (~(Hyj7z6[2] & Haciw6));
assign Equhy6 = (Kruhy6 & Sruhy6);
assign Sruhy6 = (~(Hyj7z6[1] & Aaciw6));
assign Kruhy6 = (~(Hyj7z6[5] & Vaciw6));
assign Opuhy6 = (Asuhy6 & Isuhy6);
assign Isuhy6 = (Qsuhy6 & Ysuhy6);
assign Ysuhy6 = (~(Hyj7z6[6] & Cbciw6));
assign Qsuhy6 = (~(Hyj7z6[7] & Jbciw6));
assign Asuhy6 = (Gtuhy6 & Otuhy6);
assign Otuhy6 = (~(Hyj7z6[0] & Dfk7z6[14]));
assign Gtuhy6 = (~(Hyj7z6[4] & Jkl7z6[14]));
assign Qouhy6 = (~(Xbzyx6 & Wtuhy6));
assign Wtuhy6 = (~(Euuhy6 & Muuhy6));
assign Muuhy6 = (Uuuhy6 & Cvuhy6);
assign Cvuhy6 = (Kvuhy6 & Svuhy6);
assign Svuhy6 = (~(Hyj7z6[0] & Rbk7z6[12]));
assign Kvuhy6 = (~(Hyj7z6[1] & Zlk7z6[12]));
assign Uuuhy6 = (Awuhy6 & Iwuhy6);
assign Iwuhy6 = (~(Hyj7z6[2] & Hwk7z6[12]));
assign Awuhy6 = (~(Hyj7z6[3] & P6l7z6[12]));
assign Euuhy6 = (Qwuhy6 & Ywuhy6);
assign Ywuhy6 = (Gxuhy6 & Oxuhy6);
assign Oxuhy6 = (~(Hyj7z6[4] & Xgl7z6[12]));
assign Gxuhy6 = (~(Hyj7z6[5] & Frl7z6[12]));
assign Qwuhy6 = (Wxuhy6 & Eyuhy6);
assign Eyuhy6 = (~(Hyj7z6[6] & N1m7z6[12]));
assign Wxuhy6 = (~(Hyj7z6[7] & Vbm7z6[12]));
assign Aouhy6 = (Myuhy6 & Uyuhy6);
assign Uyuhy6 = (~(Czuhy6 & Ngqyx6));
assign Czuhy6 = (~(Kzuhy6 & Szuhy6));
assign Szuhy6 = (A0vhy6 & I0vhy6);
assign I0vhy6 = (Q0vhy6 & Y0vhy6);
assign Y0vhy6 = (G1vhy6 & O1vhy6);
assign O1vhy6 = (W1vhy6 & E2vhy6);
assign E2vhy6 = (~(V40zx6 & Zdj7z6[1]));
assign W1vhy6 = (M2vhy6 & U2vhy6);
assign M2vhy6 = (~(Prqyx6 & Z3j7z6[14]));
assign G1vhy6 = (C3vhy6 & K3vhy6);
assign K3vhy6 = (~(A0j7z6[14] & Xrqyx6));
assign C3vhy6 = (~(H1j7z6[14] & Rqqyx6));
assign Q0vhy6 = (S3vhy6 & A4vhy6);
assign A4vhy6 = (I4vhy6 & Q4vhy6);
assign Q4vhy6 = (~(Dxqyx6 & P2j7z6[2]));
assign I4vhy6 = (~(Wui7z6[14] & Lxqyx6));
assign S3vhy6 = (Y4vhy6 & G5vhy6);
assign G5vhy6 = (~(Dri7z6[14] & Fwqyx6));
assign Y4vhy6 = (~(Bwi7z6[14] & Hzqyx6));
assign A0vhy6 = (O5vhy6 & W5vhy6);
assign W5vhy6 = (E6vhy6 & M6vhy6);
assign M6vhy6 = (U6vhy6 & C7vhy6);
assign C7vhy6 = (~(Svkhy6 & Pnb7z6[14]));
assign U6vhy6 = (~(D90zx6 & Lgj7z6[184]));
assign E6vhy6 = (K7vhy6 & S7vhy6);
assign S7vhy6 = (~(Za0zx6 & Lgj7z6[172]));
assign K7vhy6 = (~(Hb0zx6 & Lgj7z6[160]));
assign O5vhy6 = (A8vhy6 & I8vhy6);
assign I8vhy6 = (Q8vhy6 & Y8vhy6);
assign Y8vhy6 = (~(Vc0zx6 & Lgj7z6[148]));
assign Q8vhy6 = (~(Dd0zx6 & Lgj7z6[136]));
assign A8vhy6 = (G9vhy6 & O9vhy6);
assign O9vhy6 = (~(Be0zx6 & Lgj7z6[124]));
assign G9vhy6 = (~(Je0zx6 & Lgj7z6[112]));
assign Kzuhy6 = (W9vhy6 & Eavhy6);
assign Eavhy6 = (Mavhy6 & Uavhy6);
assign Uavhy6 = (Cbvhy6 & Kbvhy6);
assign Kbvhy6 = (Sbvhy6 & Acvhy6);
assign Acvhy6 = (~(Bi0zx6 & Lgj7z6[100]));
assign Sbvhy6 = (~(Ji0zx6 & Lgj7z6[88]));
assign Cbvhy6 = (Icvhy6 & Qcvhy6);
assign Qcvhy6 = (~(Dh0zx6 & Lgj7z6[76]));
assign Icvhy6 = (~(Hj0zx6 & Lgj7z6[64]));
assign Mavhy6 = (Ycvhy6 & Gdvhy6);
assign Gdvhy6 = (Odvhy6 & Wdvhy6);
assign Wdvhy6 = (~(Pj0zx6 & Lgj7z6[52]));
assign Odvhy6 = (~(Dl0zx6 & Lgj7z6[40]));
assign Ycvhy6 = (Eevhy6 & Mevhy6);
assign Mevhy6 = (~(Ll0zx6 & Lgj7z6[28]));
assign Eevhy6 = (~(Jm0zx6 & Lgj7z6[16]));
assign W9vhy6 = (Uevhy6 & Cfvhy6);
assign Cfvhy6 = (Kfvhy6 & Sfvhy6);
assign Sfvhy6 = (Agvhy6 & Igvhy6);
assign Igvhy6 = (~(Rm0zx6 & Lgj7z6[4]));
assign Agvhy6 = (~(Pzqyx6 & G5j7z6[46]));
assign Kfvhy6 = (Qgvhy6 & Ygvhy6);
assign Ygvhy6 = (~(Jyqyx6 & G5j7z6[14]));
assign Qgvhy6 = (~(B2ryx6 & M6j7z6[46]));
assign Uevhy6 = (Ghvhy6 & Ohvhy6);
assign Ohvhy6 = (Whvhy6 & Eivhy6);
assign Eivhy6 = (~(J2ryx6 & M6j7z6[14]));
assign Whvhy6 = (~(D1ryx6 & Ohj7z6[46]));
assign Ghvhy6 = (Mivhy6 & Uivhy6);
assign Uivhy6 = (~(X3ryx6 & Ohj7z6[14]));
assign Mivhy6 = (~(STCALIB[14] & F4ryx6));
assign Myuhy6 = (~(Klo7z6[1] & Cjvhy6));
assign Cjvhy6 = (~(Kjvhy6 & Sjvhy6));
assign Sjvhy6 = (Akvhy6 & Ikvhy6);
assign Ikvhy6 = (Qkvhy6 & Ravyx6);
assign Qkvhy6 = (~(T9tyx6 & As77z6));
assign Akvhy6 = (Ykvhy6 & Glvhy6);
assign Glvhy6 = (~(Xkq7z6[14] & B6qyx6));
assign Ykvhy6 = (~(D5qyx6 & Bqp7z6[14]));
assign Kjvhy6 = (Olvhy6 & Wlvhy6);
assign Wlvhy6 = (Emvhy6 & Mmvhy6);
assign Mmvhy6 = (~(L9qyx6 & E6p7z6[14]));
assign Emvhy6 = (~(Fcqyx6 & B2q7z6[14]));
assign Olvhy6 = (Umvhy6 & Cnvhy6);
assign Cnvhy6 = (~(Tdqyx6 & Mkp7z6[14]));
assign Umvhy6 = (~(U9p7z6[14] & Hfqyx6));
assign Knuhy6 = (Knvhy6 & Snvhy6);
assign Snvhy6 = (~(Ies7z6[14] & Tltyx6));
assign Knvhy6 = (Aovhy6 & Iovhy6);
assign Iovhy6 = (~(Klo7z6[3] & Qovhy6));
assign Qovhy6 = (~(Yovhy6 & Gpvhy6));
assign Gpvhy6 = (Opvhy6 & Wpvhy6);
assign Wpvhy6 = (Eqvhy6 & Mqvhy6);
assign Mqvhy6 = (~(Ojymz6[8] & Minhy6));
assign Eqvhy6 = (~(Unymz6[8] & Uinhy6));
assign Opvhy6 = (Uqvhy6 & Crvhy6);
assign Crvhy6 = (Kfsnv6 | Cbrhy6);
assign Kfsnv6 = (!Sgymz6[8]);
assign Uqvhy6 = (~(Biymz6[14] & Olnhy6));
assign Yovhy6 = (Krvhy6 & Srvhy6);
assign Krvhy6 = (Asvhy6 & Isvhy6);
assign Isvhy6 = (~(Zs1nz6[6] & S3mhy6));
assign Asvhy6 = (~(Nn1nz6[6] & U2mhy6));
assign Aovhy6 = (~(Klo7z6[2] & Qsvhy6));
assign Qsvhy6 = (~(Ysvhy6 & Gtvhy6));
assign Gtvhy6 = (Otvhy6 & Wtvhy6);
assign Wtvhy6 = (Euvhy6 & Muvhy6);
assign Muvhy6 = (~(M0tet6 & S4kiw6));
assign Euvhy6 = (Uuvhy6 & Cvvhy6);
assign Cvvhy6 = (~(Nqo7z6[12] & M8kiw6));
assign Uuvhy6 = (~(Fpo7z6[12] & H9kiw6));
assign Otvhy6 = (Kvvhy6 & Svvhy6);
assign Svvhy6 = (~(Ouo7z6[12] & K7kiw6));
assign Kvvhy6 = (~(Hxo7z6[12] & W6kiw6));
assign Ysvhy6 = (Awvhy6 & Iwvhy6);
assign Iwvhy6 = (Qwvhy6 & Ywvhy6);
assign Ywvhy6 = (~(Vro7z6[12] & Y7kiw6));
assign Qwvhy6 = (~(T2p7z6[14] & U5kiw6));
assign Awvhy6 = (Gxvhy6 & Oxvhy6);
assign Oxvhy6 = (~(W3p7z6[14] & G5kiw6));
assign Gxvhy6 = (~(A0p7z6[12] & I6kiw6));
assign Umuhy6 = (~(Zmoyx6 & E4f7x6));
assign Emuhy6 = (Wxvhy6 & Eyvhy6);
assign Eyvhy6 = (~(HRDATAS[14] & Ad47x6));
assign Wxvhy6 = (~(HRDATAD[14] & Mc47x6));
assign Oluhy6 = (~(Lpryx6 & Twq7x6));
assign Pmo7v6 = (~(Myvhy6 & Uyvhy6));
assign Uyvhy6 = (~(Jexmz6[15] & K94iw6));
assign Myvhy6 = (Czvhy6 & Kzvhy6);
assign Kzvhy6 = (~(Lloyx6 & Dh57x6));
assign Dh57x6 = (~(Szvhy6 & A0why6));
assign A0why6 = (I0why6 & Q0why6);
assign Q0why6 = (Bqoyx6 | K7f7x6);
assign K7f7x6 = (Y0why6 & G1why6);
assign G1why6 = (O1why6 & W1why6);
assign W1why6 = (E2why6 & M2why6);
assign M2why6 = (~(Rmzyx6 & U2why6));
assign U2why6 = (~(C3why6 & K3why6));
assign K3why6 = (S3why6 & A4why6);
assign A4why6 = (I4why6 & Q4why6);
assign Q4why6 = (~(Hyj7z6[3] & Lcciw6));
assign I4why6 = (~(Hyj7z6[2] & Ecciw6));
assign S3why6 = (Y4why6 & G5why6);
assign G5why6 = (~(Hyj7z6[1] & Xbciw6));
assign Y4why6 = (~(Hyj7z6[5] & Zcciw6));
assign C3why6 = (O5why6 & W5why6);
assign W5why6 = (E6why6 & M6why6);
assign M6why6 = (~(Hyj7z6[6] & Ndciw6));
assign E6why6 = (~(Hyj7z6[7] & Udciw6));
assign O5why6 = (U6why6 & C7why6);
assign C7why6 = (~(Hyj7z6[0] & Dfk7z6[15]));
assign U6why6 = (~(Hyj7z6[4] & Jkl7z6[15]));
assign E2why6 = (~(Xbzyx6 & K7why6));
assign K7why6 = (~(S7why6 & A8why6));
assign A8why6 = (I8why6 & Q8why6);
assign Q8why6 = (Y8why6 & G9why6);
assign G9why6 = (~(Hyj7z6[0] & Rbk7z6[13]));
assign Y8why6 = (~(Hyj7z6[1] & Zlk7z6[13]));
assign I8why6 = (O9why6 & W9why6);
assign W9why6 = (~(Hyj7z6[2] & Hwk7z6[13]));
assign O9why6 = (~(Hyj7z6[3] & P6l7z6[13]));
assign S7why6 = (Eawhy6 & Mawhy6);
assign Mawhy6 = (Uawhy6 & Cbwhy6);
assign Cbwhy6 = (~(Hyj7z6[4] & Xgl7z6[13]));
assign Uawhy6 = (~(Hyj7z6[5] & Frl7z6[13]));
assign Eawhy6 = (Kbwhy6 & Sbwhy6);
assign Sbwhy6 = (~(Hyj7z6[6] & N1m7z6[13]));
assign Kbwhy6 = (~(Hyj7z6[7] & Vbm7z6[13]));
assign O1why6 = (Acwhy6 & Icwhy6);
assign Icwhy6 = (~(Qcwhy6 & Ngqyx6));
assign Qcwhy6 = (~(Ycwhy6 & Gdwhy6));
assign Gdwhy6 = (Odwhy6 & Wdwhy6);
assign Wdwhy6 = (Eewhy6 & Mewhy6);
assign Mewhy6 = (Uewhy6 & Cfwhy6);
assign Cfwhy6 = (Kfwhy6 & Sfwhy6);
assign Sfwhy6 = (~(V40zx6 & Zdj7z6[2]));
assign Kfwhy6 = (Agwhy6 & U2vhy6);
assign Agwhy6 = (~(Prqyx6 & Z3j7z6[15]));
assign Uewhy6 = (Igwhy6 & Qgwhy6);
assign Qgwhy6 = (~(A0j7z6[15] & Xrqyx6));
assign Igwhy6 = (~(H1j7z6[15] & Rqqyx6));
assign Eewhy6 = (Ygwhy6 & Ghwhy6);
assign Ghwhy6 = (Ohwhy6 & Whwhy6);
assign Whwhy6 = (~(Bzi7z6[15] & Vsqyx6));
assign Ohwhy6 = (~(Dxqyx6 & P2j7z6[3]));
assign Ygwhy6 = (Eiwhy6 & Miwhy6);
assign Miwhy6 = (~(Wui7z6[15] & Lxqyx6));
assign Eiwhy6 = (~(Dri7z6[15] & Fwqyx6));
assign Odwhy6 = (Uiwhy6 & Cjwhy6);
assign Cjwhy6 = (Kjwhy6 & Sjwhy6);
assign Sjwhy6 = (Akwhy6 & Ikwhy6);
assign Ikwhy6 = (~(D90zx6 & Lgj7z6[185]));
assign Akwhy6 = (Qkwhy6 & Ykwhy6);
assign Ykwhy6 = (~(Bwi7z6[15] & Hzqyx6));
assign Qkwhy6 = (~(Svkhy6 & Pnb7z6[15]));
assign Kjwhy6 = (Glwhy6 & Olwhy6);
assign Olwhy6 = (~(Za0zx6 & Lgj7z6[173]));
assign Glwhy6 = (~(Hb0zx6 & Lgj7z6[161]));
assign Uiwhy6 = (Wlwhy6 & Emwhy6);
assign Emwhy6 = (Mmwhy6 & Umwhy6);
assign Umwhy6 = (~(Vc0zx6 & Lgj7z6[149]));
assign Mmwhy6 = (~(Dd0zx6 & Lgj7z6[137]));
assign Wlwhy6 = (Cnwhy6 & Knwhy6);
assign Knwhy6 = (~(Be0zx6 & Lgj7z6[125]));
assign Cnwhy6 = (~(Je0zx6 & Lgj7z6[113]));
assign Ycwhy6 = (Snwhy6 & Aowhy6);
assign Aowhy6 = (Iowhy6 & Qowhy6);
assign Qowhy6 = (Yowhy6 & Gpwhy6);
assign Gpwhy6 = (Opwhy6 & Wpwhy6);
assign Wpwhy6 = (~(Dh0zx6 & Lgj7z6[77]));
assign Opwhy6 = (Eqwhy6 & Mqwhy6);
assign Mqwhy6 = (~(Bi0zx6 & Lgj7z6[101]));
assign Eqwhy6 = (~(Ji0zx6 & Lgj7z6[89]));
assign Yowhy6 = (Uqwhy6 & Crwhy6);
assign Crwhy6 = (~(Hj0zx6 & Lgj7z6[65]));
assign Uqwhy6 = (~(Pj0zx6 & Lgj7z6[53]));
assign Iowhy6 = (Krwhy6 & Srwhy6);
assign Srwhy6 = (Aswhy6 & Iswhy6);
assign Iswhy6 = (~(Dl0zx6 & Lgj7z6[41]));
assign Aswhy6 = (~(Ll0zx6 & Lgj7z6[29]));
assign Krwhy6 = (Qswhy6 & Yswhy6);
assign Yswhy6 = (~(Jm0zx6 & Lgj7z6[17]));
assign Qswhy6 = (~(Rm0zx6 & Lgj7z6[5]));
assign Snwhy6 = (Gtwhy6 & Otwhy6);
assign Otwhy6 = (Wtwhy6 & Euwhy6);
assign Euwhy6 = (Muwhy6 & Uuwhy6);
assign Uuwhy6 = (~(Pzqyx6 & G5j7z6[47]));
assign Muwhy6 = (~(Jyqyx6 & G5j7z6[15]));
assign Wtwhy6 = (Cvwhy6 & Kvwhy6);
assign Kvwhy6 = (~(B2ryx6 & M6j7z6[47]));
assign Cvwhy6 = (~(J2ryx6 & M6j7z6[15]));
assign Gtwhy6 = (Svwhy6 & Awwhy6);
assign Awwhy6 = (Iwwhy6 & Qwwhy6);
assign Qwwhy6 = (~(D1ryx6 & Ohj7z6[47]));
assign Iwwhy6 = (~(O5nhy6 & Evadt6));
assign O5nhy6 = (!Ywwhy6);
assign Svwhy6 = (Gxwhy6 & Oxwhy6);
assign Oxwhy6 = (~(X3ryx6 & Ohj7z6[15]));
assign Gxwhy6 = (~(STCALIB[15] & F4ryx6));
assign Acwhy6 = (~(Klo7z6[1] & Wxwhy6));
assign Wxwhy6 = (~(Eywhy6 & Mywhy6));
assign Mywhy6 = (Uywhy6 & Czwhy6);
assign Czwhy6 = (Kzwhy6 & Ravyx6);
assign Kzwhy6 = (~(T9tyx6 & Sr77z6));
assign Uywhy6 = (Szwhy6 & A0xhy6);
assign A0xhy6 = (~(Xkq7z6[15] & B6qyx6));
assign Szwhy6 = (~(Bqp7z6[15] & D5qyx6));
assign Eywhy6 = (I0xhy6 & Q0xhy6);
assign Q0xhy6 = (Y0xhy6 & G1xhy6);
assign G1xhy6 = (~(E6p7z6[15] & L9qyx6));
assign Y0xhy6 = (~(B2q7z6[15] & Fcqyx6));
assign I0xhy6 = (O1xhy6 & W1xhy6);
assign W1xhy6 = (~(Mkp7z6[15] & Tdqyx6));
assign O1xhy6 = (~(Hfqyx6 & U9p7z6[15]));
assign Y0why6 = (E2xhy6 & M2xhy6);
assign M2xhy6 = (~(Ies7z6[15] & Tltyx6));
assign E2xhy6 = (U2xhy6 & C3xhy6);
assign C3xhy6 = (~(Klo7z6[3] & K3xhy6));
assign K3xhy6 = (~(S3xhy6 & A4xhy6));
assign A4xhy6 = (I4xhy6 & Q4xhy6);
assign Q4xhy6 = (Y4xhy6 & G5xhy6);
assign G5xhy6 = (~(Ojymz6[9] & Minhy6));
assign Minhy6 = (!Acrhy6);
assign Acrhy6 = (~(Hfpyx6 & Mphiw6));
assign Y4xhy6 = (~(Unymz6[9] & Uinhy6));
assign Uinhy6 = (Thpyx6 & Mphiw6);
assign I4xhy6 = (O5xhy6 & W5xhy6);
assign W5xhy6 = (~(Sgymz6[9] & Glnhy6));
assign Glnhy6 = (!Cbrhy6);
assign Cbrhy6 = (~(Ngpyx6 & Mphiw6));
assign O5xhy6 = (~(Biymz6[15] & Olnhy6));
assign Olnhy6 = (Ddpyx6 & Mphiw6);
assign S3xhy6 = (E6xhy6 & Srvhy6);
assign Srvhy6 = (M6xhy6 & U6xhy6);
assign U6xhy6 = (~(C7xhy6 & Mphiw6));
assign M6xhy6 = (~(K7xhy6 & O1mhy6));
assign K7xhy6 = (~(S7xhy6 | Oduhy6));
assign E6xhy6 = (A8xhy6 & I8xhy6);
assign I8xhy6 = (~(Zs1nz6[7] & S3mhy6));
assign A8xhy6 = (~(Nn1nz6[7] & U2mhy6));
assign U2xhy6 = (~(Klo7z6[2] & Q8xhy6));
assign Q8xhy6 = (~(Y8xhy6 & G9xhy6));
assign G9xhy6 = (O9xhy6 & W9xhy6);
assign W9xhy6 = (Eaxhy6 & Maxhy6);
assign Maxhy6 = (~(Lyset6 & S4kiw6));
assign Eaxhy6 = (Uaxhy6 & Cbxhy6);
assign Cbxhy6 = (~(Nqo7z6[13] & M8kiw6));
assign Uaxhy6 = (~(Fpo7z6[13] & H9kiw6));
assign O9xhy6 = (Kbxhy6 & Sbxhy6);
assign Sbxhy6 = (~(Ouo7z6[13] & K7kiw6));
assign Kbxhy6 = (~(Hxo7z6[13] & W6kiw6));
assign Y8xhy6 = (Acxhy6 & Icxhy6);
assign Icxhy6 = (Qcxhy6 & Ycxhy6);
assign Ycxhy6 = (~(Vro7z6[13] & Y7kiw6));
assign Qcxhy6 = (~(T2p7z6[15] & U5kiw6));
assign Acxhy6 = (Gdxhy6 & Odxhy6);
assign Odxhy6 = (~(W3p7z6[15] & G5kiw6));
assign Gdxhy6 = (~(A0p7z6[13] & I6kiw6));
assign I0why6 = (~(Zmoyx6 & R7f7x6));
assign Szvhy6 = (Wdxhy6 & Eexhy6);
assign Eexhy6 = (~(HRDATAS[15] & Ad47x6));
assign Wdxhy6 = (~(HRDATAD[15] & Mc47x6));
assign Czvhy6 = (~(Lpryx6 & Oyp7x6));
assign Imo7v6 = (~(Mexhy6 & Uexhy6));
assign Uexhy6 = (~(Jexmz6[16] & K94iw6));
assign Mexhy6 = (Cfxhy6 & Kfxhy6);
assign Kfxhy6 = (~(Lloyx6 & Ve9ov6));
assign Ve9ov6 = (~(Sfxhy6 & Agxhy6));
assign Agxhy6 = (Igxhy6 & Qgxhy6);
assign Qgxhy6 = (Bqoyx6 | G4g7x6);
assign G4g7x6 = (Ygxhy6 & Ghxhy6);
assign Ghxhy6 = (Ohxhy6 & Whxhy6);
assign Whxhy6 = (Eixhy6 & Mixhy6);
assign Mixhy6 = (~(Xbzyx6 & Uixhy6));
assign Uixhy6 = (~(Cjxhy6 & Kjxhy6));
assign Kjxhy6 = (Sjxhy6 & Akxhy6);
assign Akxhy6 = (Ikxhy6 & Qkxhy6);
assign Qkxhy6 = (~(Hyj7z6[0] & Rbk7z6[14]));
assign Ikxhy6 = (~(Hyj7z6[1] & Zlk7z6[14]));
assign Sjxhy6 = (Ykxhy6 & Glxhy6);
assign Glxhy6 = (~(Hyj7z6[2] & Hwk7z6[14]));
assign Ykxhy6 = (~(Hyj7z6[3] & P6l7z6[14]));
assign Cjxhy6 = (Olxhy6 & Wlxhy6);
assign Wlxhy6 = (Emxhy6 & Mmxhy6);
assign Mmxhy6 = (~(Hyj7z6[4] & Xgl7z6[14]));
assign Emxhy6 = (~(Hyj7z6[5] & Frl7z6[14]));
assign Olxhy6 = (Umxhy6 & Cnxhy6);
assign Cnxhy6 = (~(Hyj7z6[6] & N1m7z6[14]));
assign Umxhy6 = (~(Hyj7z6[7] & Vbm7z6[14]));
assign Eixhy6 = (Knxhy6 & Snxhy6);
assign Snxhy6 = (~(D1pyx6 & Aoxhy6));
assign Aoxhy6 = (~(Ioxhy6 & Qoxhy6));
assign Qoxhy6 = (Yoxhy6 & Gpxhy6);
assign Gpxhy6 = (~(Ojymz6[10] & Hfpyx6));
assign Yoxhy6 = (Opxhy6 & Wpxhy6);
assign Wpxhy6 = (~(Bfymz6[0] & Fgpyx6));
assign Opxhy6 = (~(Sgymz6[10] & Ngpyx6));
assign Ioxhy6 = (Eqxhy6 & Mqxhy6);
assign Mqxhy6 = (~(Blymz6[0] & Lhpyx6));
assign Eqxhy6 = (~(Unymz6[10] & Thpyx6));
assign Knxhy6 = (~(Rmzyx6 & Uqxhy6));
assign Uqxhy6 = (~(Crxhy6 & Krxhy6));
assign Krxhy6 = (Srxhy6 & Asxhy6);
assign Asxhy6 = (Isxhy6 & Qsxhy6);
assign Qsxhy6 = (~(Hyj7z6[0] & Dfk7z6[16]));
assign Isxhy6 = (~(Hyj7z6[1] & Lpk7z6[16]));
assign Srxhy6 = (Ysxhy6 & Gtxhy6);
assign Gtxhy6 = (~(Hyj7z6[2] & Tzk7z6[16]));
assign Ysxhy6 = (~(Hyj7z6[3] & Bal7z6[16]));
assign Crxhy6 = (Otxhy6 & Wtxhy6);
assign Wtxhy6 = (Euxhy6 & Muxhy6);
assign Muxhy6 = (~(Hyj7z6[4] & Jkl7z6[16]));
assign Euxhy6 = (~(Hyj7z6[5] & Rul7z6[16]));
assign Otxhy6 = (Uuxhy6 & Cvxhy6);
assign Cvxhy6 = (~(Hyj7z6[6] & Z4m7z6[16]));
assign Uuxhy6 = (~(Hyj7z6[7] & Hfm7z6[16]));
assign Ohxhy6 = (Kvxhy6 & Svxhy6);
assign Svxhy6 = (~(Klo7z6[1] & Awxhy6));
assign Awxhy6 = (~(Iwxhy6 & Qwxhy6));
assign Qwxhy6 = (Ywxhy6 & Gxxhy6);
assign Gxxhy6 = (Oxxhy6 & Wxxhy6);
assign Wxxhy6 = (~(Xkq7z6[16] & B6qyx6));
assign Oxxhy6 = (Eyxhy6 & Ravyx6);
assign Eyxhy6 = (~(T9tyx6 & Kr77z6));
assign Ywxhy6 = (Myxhy6 & Uyxhy6);
assign Uyxhy6 = (~(Bqp7z6[16] & D5qyx6));
assign Myxhy6 = (~(E6p7z6[16] & L9qyx6));
assign Iwxhy6 = (Czxhy6 & Kzxhy6);
assign Kzxhy6 = (Szxhy6 & A0yhy6);
assign A0yhy6 = (~(B2q7z6[16] & Fcqyx6));
assign Szxhy6 = (~(Q0a8x6 & Wrp7z6[0]));
assign Czxhy6 = (I0yhy6 & Q0yhy6);
assign Q0yhy6 = (~(Mkp7z6[16] & Tdqyx6));
assign I0yhy6 = (~(Hfqyx6 & U9p7z6[16]));
assign Kvxhy6 = (~(Y0yhy6 & Ngqyx6));
assign Y0yhy6 = (~(G1yhy6 & O1yhy6));
assign O1yhy6 = (W1yhy6 & E2yhy6);
assign E2yhy6 = (M2yhy6 & U2yhy6);
assign U2yhy6 = (C3yhy6 & K3yhy6);
assign K3yhy6 = (~(Prqyx6 & Ykcet6));
assign C3yhy6 = (S3yhy6 & A4yhy6);
assign A4yhy6 = (~(I4yhy6 & Buqyx6));
assign I4yhy6 = (Kdadt6 & V9lov6);
assign V9lov6 = (~(Cwadt6 & X6eet6));
assign S3yhy6 = (~(Q4yhy6 & Macet6));
assign Q4yhy6 = (~(Lxuyx6 | Hzuyx6));
assign M2yhy6 = (Y4yhy6 & G5yhy6);
assign G5yhy6 = (~(Ttqyx6 & E1cet6));
assign Y4yhy6 = (O5yhy6 & W5yhy6);
assign W5yhy6 = (~(A0j7z6[16] & Xrqyx6));
assign O5yhy6 = (~(H1j7z6[16] & Rqqyx6));
assign W1yhy6 = (E6yhy6 & M6yhy6);
assign M6yhy6 = (U6yhy6 & C7yhy6);
assign C7yhy6 = (~(Dxqyx6 & P2j7z6[4]));
assign U6yhy6 = (K7yhy6 & S7yhy6);
assign S7yhy6 = (~(Bzi7z6[16] & Vsqyx6));
assign K7yhy6 = (~(Hjsyx6 & A8yhy6));
assign E6yhy6 = (I8yhy6 & Q8yhy6);
assign Q8yhy6 = (~(Wui7z6[16] & Lxqyx6));
assign I8yhy6 = (~(Dri7z6[16] & Fwqyx6));
assign G1yhy6 = (Y8yhy6 & G9yhy6);
assign G9yhy6 = (O9yhy6 & W9yhy6);
assign W9yhy6 = (Eayhy6 & Mayhy6);
assign Mayhy6 = (~(Pzqyx6 & G5j7z6[48]));
assign Eayhy6 = (Uayhy6 & Cbyhy6);
assign Cbyhy6 = (~(Bwi7z6[16] & Hzqyx6));
assign Uayhy6 = (~(Svkhy6 & Pnb7z6[16]));
assign O9yhy6 = (Kbyhy6 & Sbyhy6);
assign Sbyhy6 = (~(J2ryx6 & M6j7z6[16]));
assign Kbyhy6 = (Acyhy6 & Icyhy6);
assign Icyhy6 = (~(Jyqyx6 & G5j7z6[16]));
assign Acyhy6 = (~(B2ryx6 & M6j7z6[48]));
assign Y8yhy6 = (Qcyhy6 & Ycyhy6);
assign Ycyhy6 = (Gdyhy6 & Odyhy6);
assign Odyhy6 = (~(STCALIB[16] & F4ryx6));
assign Gdyhy6 = (Wdyhy6 & Eeyhy6);
assign Eeyhy6 = (~(D1ryx6 & Ohj7z6[48]));
assign Wdyhy6 = (~(X3ryx6 & Ohj7z6[16]));
assign Qcyhy6 = (Pr0zx6 & Meyhy6);
assign Ygxhy6 = (Ueyhy6 & Cfyhy6);
assign Cfyhy6 = (Kfyhy6 & Sfyhy6);
assign Sfyhy6 = (~(Yr1nz6[0] & Xjtyx6));
assign Kfyhy6 = (Agyhy6 & Igyhy6);
assign Igyhy6 = (~(Klo7z6[2] & Qgyhy6));
assign Qgyhy6 = (~(Ygyhy6 & Ghyhy6));
assign Ghyhy6 = (Ohyhy6 & Whyhy6);
assign Whyhy6 = (Eiyhy6 & Miyhy6);
assign Miyhy6 = (~(Kwset6 & S4kiw6));
assign Eiyhy6 = (Uiyhy6 & Cjyhy6);
assign Cjyhy6 = (~(Nqo7z6[14] & M8kiw6));
assign Uiyhy6 = (~(Fpo7z6[14] & H9kiw6));
assign Ohyhy6 = (Kjyhy6 & Sjyhy6);
assign Sjyhy6 = (~(Ouo7z6[14] & K7kiw6));
assign Kjyhy6 = (~(Hxo7z6[14] & W6kiw6));
assign Ygyhy6 = (Akyhy6 & Ikyhy6);
assign Ikyhy6 = (Qkyhy6 & Ykyhy6);
assign Ykyhy6 = (~(Vro7z6[14] & Y7kiw6));
assign Qkyhy6 = (~(T2p7z6[16] & U5kiw6));
assign Akyhy6 = (Glyhy6 & Olyhy6);
assign Olyhy6 = (~(W3p7z6[16] & G5kiw6));
assign Glyhy6 = (~(A0p7z6[14] & I6kiw6));
assign Agyhy6 = (~(Mm1nz6[0] & Pjtyx6));
assign Ueyhy6 = (Wlyhy6 & Emyhy6);
assign Emyhy6 = (~(Mqb7z6[0] & Lltyx6));
assign Wlyhy6 = (~(Ies7z6[16] & Tltyx6));
assign Igxhy6 = (~(HRDATAS[16] & Ad47x6));
assign Sfxhy6 = (Mmyhy6 & Umyhy6);
assign Umyhy6 = (~(HRDATAD[16] & Mc47x6));
assign Mmyhy6 = (~(Zmoyx6 & N4g7x6));
assign Cfxhy6 = (~(Lpryx6 & V4r7x6));
assign Bmo7v6 = (~(Cnyhy6 & Knyhy6));
assign Knyhy6 = (~(Jexmz6[17] & K94iw6));
assign Cnyhy6 = (Snyhy6 & Aoyhy6);
assign Aoyhy6 = (~(Lloyx6 & Ob67x6));
assign Ob67x6 = (~(Ioyhy6 & Qoyhy6));
assign Qoyhy6 = (Yoyhy6 & Gpyhy6);
assign Gpyhy6 = (Bqoyx6 | Tff7x6);
assign Tff7x6 = (Opyhy6 & Wpyhy6);
assign Wpyhy6 = (Eqyhy6 & Mqyhy6);
assign Mqyhy6 = (Uqyhy6 & Cryhy6);
assign Cryhy6 = (~(Xbzyx6 & Kryhy6));
assign Kryhy6 = (~(Sryhy6 & Asyhy6));
assign Asyhy6 = (Isyhy6 & Qsyhy6);
assign Qsyhy6 = (Ysyhy6 & Gtyhy6);
assign Gtyhy6 = (~(Hyj7z6[0] & Rbk7z6[15]));
assign Ysyhy6 = (~(Hyj7z6[1] & Zlk7z6[15]));
assign Isyhy6 = (Otyhy6 & Wtyhy6);
assign Wtyhy6 = (~(Hyj7z6[2] & Hwk7z6[15]));
assign Otyhy6 = (~(Hyj7z6[3] & P6l7z6[15]));
assign Sryhy6 = (Euyhy6 & Muyhy6);
assign Muyhy6 = (Uuyhy6 & Cvyhy6);
assign Cvyhy6 = (~(Hyj7z6[4] & Xgl7z6[15]));
assign Uuyhy6 = (~(Hyj7z6[5] & Frl7z6[15]));
assign Euyhy6 = (Kvyhy6 & Svyhy6);
assign Svyhy6 = (~(Hyj7z6[6] & N1m7z6[15]));
assign Kvyhy6 = (~(Hyj7z6[7] & Vbm7z6[15]));
assign Uqyhy6 = (Awyhy6 & Iwyhy6);
assign Iwyhy6 = (~(D1pyx6 & Qwyhy6));
assign Qwyhy6 = (~(Ywyhy6 & Gxyhy6));
assign Gxyhy6 = (~(Blymz6[1] & Lhpyx6));
assign Ywyhy6 = (Oxyhy6 & L5pyx6);
assign L5pyx6 = (~(P3xyx6 & N8pyx6));
assign N8pyx6 = (Wxyhy6 & Xfymz6[4]);
assign Wxyhy6 = (Xfymz6[2] & Eyyhy6);
assign Oxyhy6 = (~(Bfymz6[1] & Fgpyx6));
assign Awyhy6 = (~(Rmzyx6 & Myyhy6));
assign Myyhy6 = (~(Uyyhy6 & Czyhy6));
assign Czyhy6 = (Kzyhy6 & Szyhy6);
assign Szyhy6 = (A0zhy6 & I0zhy6);
assign I0zhy6 = (~(Hyj7z6[3] & Ahciw6));
assign A0zhy6 = (~(Hyj7z6[2] & Tgciw6));
assign Kzyhy6 = (Q0zhy6 & Y0zhy6);
assign Y0zhy6 = (~(Hyj7z6[1] & Mgciw6));
assign Q0zhy6 = (~(Hyj7z6[5] & Hhciw6));
assign Uyyhy6 = (G1zhy6 & O1zhy6);
assign O1zhy6 = (W1zhy6 & E2zhy6);
assign E2zhy6 = (~(Hyj7z6[6] & Ohciw6));
assign W1zhy6 = (~(Hyj7z6[7] & Vhciw6));
assign G1zhy6 = (M2zhy6 & U2zhy6);
assign U2zhy6 = (~(Hyj7z6[0] & Dfk7z6[17]));
assign M2zhy6 = (~(Hyj7z6[4] & Jkl7z6[17]));
assign Eqyhy6 = (C3zhy6 & K3zhy6);
assign K3zhy6 = (~(Klo7z6[1] & S3zhy6));
assign S3zhy6 = (~(A4zhy6 & I4zhy6));
assign I4zhy6 = (Q4zhy6 & Y4zhy6);
assign Y4zhy6 = (G5zhy6 & O5zhy6);
assign O5zhy6 = (~(Xkq7z6[17] & B6qyx6));
assign G5zhy6 = (W5zhy6 & Ravyx6);
assign W5zhy6 = (~(T9tyx6 & Cr77z6));
assign Q4zhy6 = (E6zhy6 & M6zhy6);
assign M6zhy6 = (~(Bqp7z6[17] & D5qyx6));
assign E6zhy6 = (~(E6p7z6[17] & L9qyx6));
assign A4zhy6 = (U6zhy6 & C7zhy6);
assign C7zhy6 = (K7zhy6 & S7zhy6);
assign S7zhy6 = (~(B2q7z6[17] & Fcqyx6));
assign K7zhy6 = (~(Q0a8x6 & Wrp7z6[1]));
assign U6zhy6 = (A8zhy6 & I8zhy6);
assign I8zhy6 = (~(Mkp7z6[17] & Tdqyx6));
assign A8zhy6 = (~(Hfqyx6 & U9p7z6[17]));
assign C3zhy6 = (~(Q8zhy6 & Ngqyx6));
assign Q8zhy6 = (~(Y8zhy6 & G9zhy6));
assign G9zhy6 = (O9zhy6 & W9zhy6);
assign W9zhy6 = (Eazhy6 & Mazhy6);
assign Mazhy6 = (Uazhy6 & Cbzhy6);
assign Cbzhy6 = (~(A0j7z6[17] & Xrqyx6));
assign Uazhy6 = (Kbzhy6 & U2vhy6);
assign Kbzhy6 = (~(Prqyx6 & Sjcet6));
assign Eazhy6 = (Sbzhy6 & Aczhy6);
assign Aczhy6 = (~(H1j7z6[17] & Rqqyx6));
assign Sbzhy6 = (~(Ttqyx6 & Oecet6));
assign O9zhy6 = (Iczhy6 & Qczhy6);
assign Qczhy6 = (Yczhy6 & Gdzhy6);
assign Gdzhy6 = (~(Dxqyx6 & P2j7z6[5]));
assign Yczhy6 = (Odzhy6 & Wdzhy6);
assign Wdzhy6 = (~(Buqyx6 & F02nv6));
assign Odzhy6 = (~(Bzi7z6[17] & Vsqyx6));
assign Iczhy6 = (Eezhy6 & Mezhy6);
assign Mezhy6 = (~(Wui7z6[17] & Lxqyx6));
assign Eezhy6 = (~(Dri7z6[17] & Fwqyx6));
assign Y8zhy6 = (Uezhy6 & Cfzhy6);
assign Cfzhy6 = (Kfzhy6 & Sfzhy6);
assign Sfzhy6 = (Agzhy6 & Igzhy6);
assign Igzhy6 = (~(Pzqyx6 & G5j7z6[49]));
assign Agzhy6 = (Qgzhy6 & Ygzhy6);
assign Ygzhy6 = (~(Bwi7z6[17] & Hzqyx6));
assign Qgzhy6 = (~(Svkhy6 & Pnb7z6[17]));
assign Kfzhy6 = (Ghzhy6 & Ohzhy6);
assign Ohzhy6 = (~(Jyqyx6 & G5j7z6[17]));
assign Ghzhy6 = (~(B2ryx6 & M6j7z6[49]));
assign Uezhy6 = (Whzhy6 & Eizhy6);
assign Eizhy6 = (Mizhy6 & Uizhy6);
assign Uizhy6 = (~(J2ryx6 & M6j7z6[17]));
assign Mizhy6 = (~(D1ryx6 & Ohj7z6[49]));
assign Whzhy6 = (Cjzhy6 & Kjzhy6);
assign Kjzhy6 = (~(X3ryx6 & Ohj7z6[17]));
assign Cjzhy6 = (~(STCALIB[17] & F4ryx6));
assign Opyhy6 = (Sjzhy6 & Akzhy6);
assign Akzhy6 = (Ikzhy6 & Qkzhy6);
assign Qkzhy6 = (~(Yr1nz6[1] & Xjtyx6));
assign Ikzhy6 = (Ykzhy6 & Glzhy6);
assign Glzhy6 = (~(Klo7z6[2] & Olzhy6));
assign Olzhy6 = (~(Wlzhy6 & Emzhy6));
assign Emzhy6 = (Mmzhy6 & Umzhy6);
assign Umzhy6 = (Cnzhy6 & Knzhy6);
assign Knzhy6 = (~(Juset6 & S4kiw6));
assign Cnzhy6 = (Snzhy6 & Aozhy6);
assign Aozhy6 = (~(Nqo7z6[15] & M8kiw6));
assign Snzhy6 = (~(Fpo7z6[15] & H9kiw6));
assign Mmzhy6 = (Iozhy6 & Qozhy6);
assign Qozhy6 = (~(Ouo7z6[15] & K7kiw6));
assign Iozhy6 = (~(Hxo7z6[15] & W6kiw6));
assign Wlzhy6 = (Yozhy6 & Gpzhy6);
assign Gpzhy6 = (Opzhy6 & Wpzhy6);
assign Wpzhy6 = (~(Vro7z6[15] & Y7kiw6));
assign Opzhy6 = (~(T2p7z6[17] & U5kiw6));
assign Yozhy6 = (Eqzhy6 & Mqzhy6);
assign Mqzhy6 = (~(W3p7z6[17] & G5kiw6));
assign Eqzhy6 = (~(A0p7z6[15] & I6kiw6));
assign Ykzhy6 = (~(Mm1nz6[1] & Pjtyx6));
assign Sjzhy6 = (Uqzhy6 & Crzhy6);
assign Crzhy6 = (~(Mqb7z6[1] & Lltyx6));
assign Uqzhy6 = (~(Ies7z6[17] & Tltyx6));
assign Yoyhy6 = (~(Zmoyx6 & Agf7x6));
assign Agf7x6 = (~(Krzhy6 & Srzhy6));
assign Srzhy6 = (~(Aszhy6 & Eaa7z6));
assign Eaa7z6 = (~(Iszhy6 & Qszhy6));
assign Qszhy6 = (~(HRDATAD[17] & Qln7z6[0]));
assign Iszhy6 = (~(HRDATAS[17] & Qln7z6[1]));
assign Krzhy6 = (~(Tim7z6[17] & Yszhy6));
assign Ioyhy6 = (Gtzhy6 & Otzhy6);
assign Otzhy6 = (~(HRDATAS[17] & Ad47x6));
assign Gtzhy6 = (~(HRDATAD[17] & Mc47x6));
assign Snyhy6 = (~(Lpryx6 & Y3q7x6));
assign Ulo7v6 = (~(Wtzhy6 & Euzhy6));
assign Euzhy6 = (~(Jexmz6[18] & K94iw6));
assign Wtzhy6 = (Muzhy6 & Uuzhy6);
assign Uuzhy6 = (~(Lloyx6 & Ddfov6));
assign Ddfov6 = (~(Cvzhy6 & Kvzhy6));
assign Kvzhy6 = (Svzhy6 & Awzhy6);
assign Awzhy6 = (Bqoyx6 | Gjf7x6);
assign Gjf7x6 = (Iwzhy6 & Qwzhy6);
assign Qwzhy6 = (Ywzhy6 & Gxzhy6);
assign Gxzhy6 = (Oxzhy6 & Wxzhy6);
assign Wxzhy6 = (~(Rmzyx6 & Eyzhy6));
assign Eyzhy6 = (~(Myzhy6 & Uyzhy6));
assign Uyzhy6 = (Czzhy6 & Kzzhy6);
assign Kzzhy6 = (Szzhy6 & A00iy6);
assign A00iy6 = (~(Hyj7z6[7] & Ljciw6));
assign Szzhy6 = (~(Hyj7z6[3] & Qiciw6));
assign Czzhy6 = (I00iy6 & Q00iy6);
assign Q00iy6 = (~(Hyj7z6[2] & Jiciw6));
assign I00iy6 = (~(Hyj7z6[1] & Ciciw6));
assign Myzhy6 = (Y00iy6 & G10iy6);
assign G10iy6 = (O10iy6 & W10iy6);
assign W10iy6 = (~(Hyj7z6[5] & Xiciw6));
assign O10iy6 = (~(Hyj7z6[6] & Ejciw6));
assign Y00iy6 = (E20iy6 & M20iy6);
assign M20iy6 = (~(Hyj7z6[0] & Dfk7z6[18]));
assign E20iy6 = (~(Hyj7z6[4] & Jkl7z6[18]));
assign Oxzhy6 = (~(Xbzyx6 & U20iy6));
assign U20iy6 = (~(C30iy6 & K30iy6));
assign K30iy6 = (S30iy6 & A40iy6);
assign A40iy6 = (I40iy6 & Q40iy6);
assign Q40iy6 = (~(Rbk7z6[16] & Hyj7z6[0]));
assign I40iy6 = (~(Zlk7z6[16] & Hyj7z6[1]));
assign S30iy6 = (Y40iy6 & G50iy6);
assign G50iy6 = (~(Hwk7z6[16] & Hyj7z6[2]));
assign Y40iy6 = (~(P6l7z6[16] & Hyj7z6[3]));
assign C30iy6 = (O50iy6 & W50iy6);
assign W50iy6 = (E60iy6 & M60iy6);
assign M60iy6 = (~(Xgl7z6[16] & Hyj7z6[4]));
assign E60iy6 = (~(Frl7z6[16] & Hyj7z6[5]));
assign O50iy6 = (U60iy6 & C70iy6);
assign C70iy6 = (~(N1m7z6[16] & Hyj7z6[6]));
assign U60iy6 = (~(Vbm7z6[16] & Hyj7z6[7]));
assign Ywzhy6 = (K70iy6 & S70iy6);
assign S70iy6 = (~(A80iy6 & Ngqyx6));
assign A80iy6 = (~(I80iy6 & Q80iy6));
assign Q80iy6 = (Y80iy6 & G90iy6);
assign G90iy6 = (O90iy6 & W90iy6);
assign W90iy6 = (Ea0iy6 & Ma0iy6);
assign Ma0iy6 = (~(Prqyx6 & Micet6));
assign Prqyx6 = (~(Ua0iy6 | Tlqyx6));
assign O90iy6 = (Cb0iy6 & Kb0iy6);
assign Kb0iy6 = (~(A0j7z6[18] & Xrqyx6));
assign Cb0iy6 = (~(H1j7z6[18] & Rqqyx6));
assign Y80iy6 = (Sb0iy6 & Ac0iy6);
assign Ac0iy6 = (Ic0iy6 & Qc0iy6);
assign Qc0iy6 = (~(Bzi7z6[18] & Vsqyx6));
assign Ic0iy6 = (Yc0iy6 & Gd0iy6);
assign Gd0iy6 = (~(Vzbet6 & Ttqyx6));
assign Yc0iy6 = (~(Buqyx6 & Cqiiw6));
assign Cqiiw6 = (!K3jnv6);
assign Sb0iy6 = (Od0iy6 & Wd0iy6);
assign Wd0iy6 = (~(Dxqyx6 & P2j7z6[6]));
assign Od0iy6 = (~(Wui7z6[18] & Lxqyx6));
assign I80iy6 = (Ee0iy6 & Me0iy6);
assign Me0iy6 = (Ue0iy6 & Cf0iy6);
assign Cf0iy6 = (Kf0iy6 & Sf0iy6);
assign Sf0iy6 = (~(Svkhy6 & Pnb7z6[18]));
assign Kf0iy6 = (Ag0iy6 & Ig0iy6);
assign Ig0iy6 = (~(Dri7z6[18] & Fwqyx6));
assign Ag0iy6 = (~(Bwi7z6[18] & Hzqyx6));
assign Ue0iy6 = (Qg0iy6 & Yg0iy6);
assign Yg0iy6 = (~(Pzqyx6 & G5j7z6[50]));
assign Qg0iy6 = (~(Jyqyx6 & G5j7z6[18]));
assign Ee0iy6 = (Gh0iy6 & Oh0iy6);
assign Oh0iy6 = (Wh0iy6 & Ei0iy6);
assign Ei0iy6 = (~(D1ryx6 & Ohj7z6[50]));
assign Wh0iy6 = (Mi0iy6 & Ui0iy6);
assign Ui0iy6 = (~(B2ryx6 & M6j7z6[50]));
assign Mi0iy6 = (~(J2ryx6 & M6j7z6[18]));
assign Gh0iy6 = (Cj0iy6 & Kj0iy6);
assign Kj0iy6 = (~(X3ryx6 & Ohj7z6[18]));
assign Cj0iy6 = (~(STCALIB[18] & F4ryx6));
assign K70iy6 = (~(Klo7z6[1] & Sj0iy6));
assign Sj0iy6 = (~(Ak0iy6 & Ik0iy6));
assign Ik0iy6 = (Qk0iy6 & Yk0iy6);
assign Yk0iy6 = (Gl0iy6 & Ravyx6);
assign Gl0iy6 = (~(T9tyx6 & Uq77z6));
assign Qk0iy6 = (Ol0iy6 & Wl0iy6);
assign Wl0iy6 = (~(Xkq7z6[18] & B6qyx6));
assign Ol0iy6 = (~(Bqp7z6[18] & D5qyx6));
assign Ak0iy6 = (Em0iy6 & Mm0iy6);
assign Mm0iy6 = (Um0iy6 & Cn0iy6);
assign Cn0iy6 = (~(E6p7z6[18] & L9qyx6));
assign Um0iy6 = (~(B2q7z6[18] & Fcqyx6));
assign Em0iy6 = (Kn0iy6 & Sn0iy6);
assign Sn0iy6 = (~(Mkp7z6[18] & Tdqyx6));
assign Kn0iy6 = (~(Hfqyx6 & U9p7z6[18]));
assign Iwzhy6 = (Ao0iy6 & Io0iy6);
assign Io0iy6 = (Qo0iy6 & Yo0iy6);
assign Yo0iy6 = (~(Klo7z6[3] & Gp0iy6));
assign Gp0iy6 = (~(Op0iy6 & Wp0iy6));
assign Wp0iy6 = (Eq0iy6 & Mq0iy6);
assign Mq0iy6 = (~(Kzlhy6 & Uq0iy6));
assign Uq0iy6 = (~(Cr0iy6 & Kr0iy6));
assign Kzlhy6 = (!Oduhy6);
assign Eq0iy6 = (~(Mphiw6 & Sr0iy6));
assign Sr0iy6 = (~(As0iy6 & Wtshy6));
assign Wtshy6 = (Z6yyx6 & Q8rhy6);
assign Q8rhy6 = (~(Ied8x6 & W5qhy6));
assign Z6yyx6 = (!C7xhy6);
assign As0iy6 = (Is0iy6 & Qs0iy6);
assign Qs0iy6 = (~(Ys0iy6 & Dp77v6));
assign Is0iy6 = (~(Blymz6[2] & Lhpyx6));
assign Op0iy6 = (Gt0iy6 & Ot0iy6);
assign Ot0iy6 = (~(Yr1nz6[2] & S3mhy6));
assign Gt0iy6 = (~(Mm1nz6[2] & U2mhy6));
assign Qo0iy6 = (~(Klo7z6[2] & Wt0iy6));
assign Wt0iy6 = (~(Eu0iy6 & Mu0iy6));
assign Mu0iy6 = (Uu0iy6 & Cv0iy6);
assign Cv0iy6 = (Kv0iy6 & Sv0iy6);
assign Sv0iy6 = (~(Isset6 & S4kiw6));
assign Kv0iy6 = (Aw0iy6 & Iw0iy6);
assign Iw0iy6 = (~(Nqo7z6[16] & M8kiw6));
assign Aw0iy6 = (~(Fpo7z6[16] & H9kiw6));
assign Uu0iy6 = (Qw0iy6 & Yw0iy6);
assign Yw0iy6 = (~(Ouo7z6[16] & K7kiw6));
assign Qw0iy6 = (~(Hxo7z6[16] & W6kiw6));
assign Eu0iy6 = (Gx0iy6 & Ox0iy6);
assign Ox0iy6 = (Wx0iy6 & Ey0iy6);
assign Ey0iy6 = (~(Vro7z6[16] & Y7kiw6));
assign Wx0iy6 = (~(T2p7z6[18] & U5kiw6));
assign Gx0iy6 = (My0iy6 & Uy0iy6);
assign Uy0iy6 = (~(W3p7z6[18] & G5kiw6));
assign My0iy6 = (~(A0p7z6[16] & I6kiw6));
assign Ao0iy6 = (Cz0iy6 & Kz0iy6);
assign Kz0iy6 = (~(Mqb7z6[2] & Lltyx6));
assign Cz0iy6 = (~(Ies7z6[18] & Tltyx6));
assign Svzhy6 = (~(Zmoyx6 & Njf7x6));
assign Njf7x6 = (~(Sz0iy6 & A01iy6));
assign A01iy6 = (~(Aszhy6 & W9a7z6));
assign W9a7z6 = (~(I01iy6 & Q01iy6));
assign Q01iy6 = (~(HRDATAD[18] & Qln7z6[0]));
assign I01iy6 = (~(HRDATAS[18] & Qln7z6[1]));
assign Sz0iy6 = (~(Tim7z6[18] & Yszhy6));
assign Cvzhy6 = (Y01iy6 & G11iy6);
assign G11iy6 = (~(HRDATAS[18] & Ad47x6));
assign Y01iy6 = (~(HRDATAD[18] & Mc47x6));
assign Muzhy6 = (~(Lpryx6 & I9q7x6));
assign Nlo7v6 = (~(O11iy6 & W11iy6));
assign W11iy6 = (~(Jexmz6[19] & K94iw6));
assign O11iy6 = (E21iy6 & M21iy6);
assign M21iy6 = (~(Lloyx6 & Hnlov6));
assign Hnlov6 = (~(U21iy6 & C31iy6));
assign C31iy6 = (K31iy6 & S31iy6);
assign S31iy6 = (Bqoyx6 | Tmf7x6);
assign Tmf7x6 = (A41iy6 & I41iy6);
assign I41iy6 = (Q41iy6 & Y41iy6);
assign Y41iy6 = (G51iy6 & O51iy6);
assign O51iy6 = (~(Xbzyx6 & W51iy6));
assign W51iy6 = (~(E61iy6 & M61iy6));
assign M61iy6 = (U61iy6 & C71iy6);
assign C71iy6 = (K71iy6 & S71iy6);
assign S71iy6 = (~(Hyj7z6[0] & Rbk7z6[17]));
assign K71iy6 = (~(Hyj7z6[1] & Zlk7z6[17]));
assign U61iy6 = (A81iy6 & I81iy6);
assign I81iy6 = (~(Hyj7z6[2] & Hwk7z6[17]));
assign A81iy6 = (~(Hyj7z6[3] & P6l7z6[17]));
assign E61iy6 = (Q81iy6 & Y81iy6);
assign Y81iy6 = (G91iy6 & O91iy6);
assign O91iy6 = (~(Hyj7z6[4] & Xgl7z6[17]));
assign G91iy6 = (~(Hyj7z6[5] & Frl7z6[17]));
assign Q81iy6 = (W91iy6 & Ea1iy6);
assign Ea1iy6 = (~(Hyj7z6[6] & N1m7z6[17]));
assign W91iy6 = (~(Hyj7z6[7] & Vbm7z6[17]));
assign G51iy6 = (Ma1iy6 & Ua1iy6);
assign Ua1iy6 = (~(Cb1iy6 & Blymz6[3]));
assign Cb1iy6 = (D1pyx6 & Lhpyx6);
assign Ma1iy6 = (~(Rmzyx6 & Kb1iy6));
assign Kb1iy6 = (~(Sb1iy6 & Ac1iy6));
assign Ac1iy6 = (Ic1iy6 & Qc1iy6);
assign Qc1iy6 = (Yc1iy6 & Gd1iy6);
assign Gd1iy6 = (~(Hyj7z6[3] & Gkciw6));
assign Yc1iy6 = (~(Hyj7z6[2] & Zjciw6));
assign Ic1iy6 = (Od1iy6 & Wd1iy6);
assign Wd1iy6 = (~(Hyj7z6[1] & Sjciw6));
assign Od1iy6 = (~(Hyj7z6[5] & Nkciw6));
assign Sb1iy6 = (Ee1iy6 & Me1iy6);
assign Me1iy6 = (Ue1iy6 & Cf1iy6);
assign Cf1iy6 = (~(Hyj7z6[6] & Ukciw6));
assign Ue1iy6 = (~(Hyj7z6[7] & Blciw6));
assign Ee1iy6 = (Kf1iy6 & Sf1iy6);
assign Sf1iy6 = (~(Hyj7z6[0] & Dfk7z6[19]));
assign Kf1iy6 = (~(Hyj7z6[4] & Jkl7z6[19]));
assign Q41iy6 = (Ag1iy6 & Ig1iy6);
assign Ig1iy6 = (~(Klo7z6[1] & Qg1iy6));
assign Qg1iy6 = (~(Yg1iy6 & Gh1iy6));
assign Gh1iy6 = (Oh1iy6 & Wh1iy6);
assign Wh1iy6 = (Ei1iy6 & Ravyx6);
assign Ei1iy6 = (~(T9tyx6 & Mq77z6));
assign Oh1iy6 = (Mi1iy6 & Ui1iy6);
assign Ui1iy6 = (~(Xkq7z6[19] & B6qyx6));
assign Mi1iy6 = (~(Bqp7z6[19] & D5qyx6));
assign Yg1iy6 = (Cj1iy6 & Kj1iy6);
assign Kj1iy6 = (Sj1iy6 & Ak1iy6);
assign Ak1iy6 = (~(E6p7z6[19] & L9qyx6));
assign Sj1iy6 = (~(B2q7z6[19] & Fcqyx6));
assign Cj1iy6 = (Ik1iy6 & Qk1iy6);
assign Qk1iy6 = (~(Mkp7z6[19] & Tdqyx6));
assign Ik1iy6 = (~(Hfqyx6 & U9p7z6[19]));
assign Ag1iy6 = (~(Yk1iy6 & Ngqyx6));
assign Yk1iy6 = (~(Gl1iy6 & Ol1iy6));
assign Ol1iy6 = (Wl1iy6 & Em1iy6);
assign Em1iy6 = (Mm1iy6 & Um1iy6);
assign Um1iy6 = (Cn1iy6 & Kn1iy6);
assign Kn1iy6 = (~(H1j7z6[19] & Rqqyx6));
assign Cn1iy6 = (Sn1iy6 & U2vhy6);
assign Sn1iy6 = (~(A0j7z6[19] & Xrqyx6));
assign Mm1iy6 = (Ao1iy6 & Io1iy6);
assign Io1iy6 = (~(Nybet6 & Ttqyx6));
assign Ao1iy6 = (~(Buqyx6 & Lua7x6));
assign Lua7x6 = (!Mhh7v6);
assign Wl1iy6 = (Qo1iy6 & Yo1iy6);
assign Yo1iy6 = (Gp1iy6 & Op1iy6);
assign Op1iy6 = (~(Bzi7z6[19] & Vsqyx6));
assign Gp1iy6 = (~(Wui7z6[19] & Lxqyx6));
assign Qo1iy6 = (Wp1iy6 & Eq1iy6);
assign Eq1iy6 = (~(Dri7z6[19] & Fwqyx6));
assign Wp1iy6 = (~(Bwi7z6[19] & Hzqyx6));
assign Gl1iy6 = (Mq1iy6 & Uq1iy6);
assign Uq1iy6 = (Cr1iy6 & Kr1iy6);
assign Kr1iy6 = (Sr1iy6 & As1iy6);
assign As1iy6 = (~(Svkhy6 & Pnb7z6[19]));
assign Sr1iy6 = (~(Pzqyx6 & G5j7z6[51]));
assign Cr1iy6 = (Is1iy6 & Qs1iy6);
assign Qs1iy6 = (~(Jyqyx6 & G5j7z6[19]));
assign Is1iy6 = (~(B2ryx6 & M6j7z6[51]));
assign Mq1iy6 = (Ys1iy6 & Gt1iy6);
assign Gt1iy6 = (Ot1iy6 & Wt1iy6);
assign Wt1iy6 = (~(J2ryx6 & M6j7z6[19]));
assign Ot1iy6 = (~(D1ryx6 & Ohj7z6[51]));
assign Ys1iy6 = (Eu1iy6 & Mu1iy6);
assign Mu1iy6 = (~(X3ryx6 & Ohj7z6[19]));
assign Eu1iy6 = (~(STCALIB[19] & F4ryx6));
assign A41iy6 = (Uu1iy6 & Cv1iy6);
assign Cv1iy6 = (Kv1iy6 & Sv1iy6);
assign Sv1iy6 = (~(Yr1nz6[3] & Xjtyx6));
assign Kv1iy6 = (Aw1iy6 & Iw1iy6);
assign Iw1iy6 = (~(Klo7z6[2] & Qw1iy6));
assign Qw1iy6 = (~(Yw1iy6 & Gx1iy6));
assign Gx1iy6 = (Ox1iy6 & Wx1iy6);
assign Wx1iy6 = (Ey1iy6 & My1iy6);
assign My1iy6 = (~(Hqset6 & S4kiw6));
assign Ey1iy6 = (Uy1iy6 & Cz1iy6);
assign Cz1iy6 = (~(Nqo7z6[17] & M8kiw6));
assign Uy1iy6 = (~(Fpo7z6[17] & H9kiw6));
assign Ox1iy6 = (Kz1iy6 & Sz1iy6);
assign Sz1iy6 = (~(Ouo7z6[17] & K7kiw6));
assign Kz1iy6 = (~(Hxo7z6[17] & W6kiw6));
assign Yw1iy6 = (A02iy6 & I02iy6);
assign I02iy6 = (Q02iy6 & Y02iy6);
assign Y02iy6 = (~(Vro7z6[17] & Y7kiw6));
assign Q02iy6 = (~(T2p7z6[19] & U5kiw6));
assign A02iy6 = (G12iy6 & O12iy6);
assign O12iy6 = (~(W3p7z6[19] & G5kiw6));
assign G12iy6 = (~(A0p7z6[17] & I6kiw6));
assign Aw1iy6 = (~(Mm1nz6[3] & Pjtyx6));
assign Uu1iy6 = (W12iy6 & E22iy6);
assign E22iy6 = (~(Mqb7z6[3] & Lltyx6));
assign W12iy6 = (~(Ies7z6[19] & Tltyx6));
assign K31iy6 = (~(Zmoyx6 & Anf7x6));
assign Anf7x6 = (~(M22iy6 & U22iy6));
assign U22iy6 = (~(Aszhy6 & O9a7z6));
assign O9a7z6 = (~(C32iy6 & K32iy6));
assign K32iy6 = (~(HRDATAD[19] & Qln7z6[0]));
assign C32iy6 = (~(HRDATAS[19] & Qln7z6[1]));
assign M22iy6 = (~(Tim7z6[19] & Yszhy6));
assign U21iy6 = (S32iy6 & A42iy6);
assign A42iy6 = (~(HRDATAS[19] & Ad47x6));
assign S32iy6 = (~(HRDATAD[19] & Mc47x6));
assign E21iy6 = (~(Lpryx6 & Seq7x6));
assign Glo7v6 = (~(I42iy6 & Q42iy6));
assign Q42iy6 = (~(Jexmz6[20] & K94iw6));
assign I42iy6 = (Y42iy6 & G52iy6);
assign G52iy6 = (~(Lloyx6 & Ax57x6));
assign Ax57x6 = (~(O52iy6 & W52iy6));
assign W52iy6 = (E62iy6 & M62iy6);
assign M62iy6 = (Bqoyx6 | Gqf7x6);
assign Gqf7x6 = (U62iy6 & C72iy6);
assign C72iy6 = (K72iy6 & S72iy6);
assign S72iy6 = (A82iy6 & I82iy6);
assign I82iy6 = (~(Klo7z6[1] & Q82iy6));
assign Q82iy6 = (~(Y82iy6 & G92iy6));
assign G92iy6 = (O92iy6 & W92iy6);
assign W92iy6 = (Ea2iy6 & Ravyx6);
assign Ea2iy6 = (~(T9tyx6 & Eq77z6));
assign O92iy6 = (Ma2iy6 & Ua2iy6);
assign Ua2iy6 = (~(Xkq7z6[20] & B6qyx6));
assign Ma2iy6 = (~(Bqp7z6[20] & D5qyx6));
assign Y82iy6 = (Cb2iy6 & Kb2iy6);
assign Kb2iy6 = (Sb2iy6 & Ac2iy6);
assign Ac2iy6 = (~(E6p7z6[20] & L9qyx6));
assign Sb2iy6 = (~(B2q7z6[20] & Fcqyx6));
assign Cb2iy6 = (Ic2iy6 & Qc2iy6);
assign Qc2iy6 = (~(Mkp7z6[20] & Tdqyx6));
assign Ic2iy6 = (~(Hfqyx6 & U9p7z6[20]));
assign A82iy6 = (Yc2iy6 & Gd2iy6);
assign Yc2iy6 = (~(Rmzyx6 & Od2iy6));
assign Od2iy6 = (~(Wd2iy6 & Ee2iy6));
assign Ee2iy6 = (Me2iy6 & Ue2iy6);
assign Ue2iy6 = (Cf2iy6 & Kf2iy6);
assign Kf2iy6 = (~(Hyj7z6[3] & Wlciw6));
assign Cf2iy6 = (~(Hyj7z6[2] & Plciw6));
assign Me2iy6 = (Sf2iy6 & Ag2iy6);
assign Ag2iy6 = (~(Hyj7z6[1] & Ilciw6));
assign Sf2iy6 = (~(Hyj7z6[5] & Dmciw6));
assign Wd2iy6 = (Ig2iy6 & Qg2iy6);
assign Qg2iy6 = (Yg2iy6 & Gh2iy6);
assign Gh2iy6 = (~(Hyj7z6[6] & Kmciw6));
assign Yg2iy6 = (~(Hyj7z6[7] & Rmciw6));
assign Ig2iy6 = (Oh2iy6 & Wh2iy6);
assign Wh2iy6 = (~(Hyj7z6[0] & Dfk7z6[20]));
assign Oh2iy6 = (~(Hyj7z6[4] & Jkl7z6[20]));
assign K72iy6 = (Ei2iy6 & Mi2iy6);
assign Mi2iy6 = (~(Klo7z6[2] & Ui2iy6));
assign Ui2iy6 = (~(Cj2iy6 & Kj2iy6));
assign Kj2iy6 = (Sj2iy6 & Ak2iy6);
assign Ak2iy6 = (Ik2iy6 & Qk2iy6);
assign Qk2iy6 = (~(Goset6 & S4kiw6));
assign Ik2iy6 = (Yk2iy6 & Gl2iy6);
assign Gl2iy6 = (~(Nqo7z6[18] & M8kiw6));
assign Yk2iy6 = (~(Fpo7z6[18] & H9kiw6));
assign Sj2iy6 = (Ol2iy6 & Wl2iy6);
assign Wl2iy6 = (~(Ouo7z6[18] & K7kiw6));
assign Ol2iy6 = (~(Hxo7z6[18] & W6kiw6));
assign Cj2iy6 = (Em2iy6 & Mm2iy6);
assign Mm2iy6 = (Um2iy6 & Cn2iy6);
assign Cn2iy6 = (~(Vro7z6[18] & Y7kiw6));
assign Um2iy6 = (~(T2p7z6[20] & U5kiw6));
assign Em2iy6 = (Kn2iy6 & Sn2iy6);
assign Sn2iy6 = (~(W3p7z6[20] & G5kiw6));
assign Kn2iy6 = (~(A0p7z6[18] & I6kiw6));
assign Ei2iy6 = (Ao2iy6 & Io2iy6);
assign Io2iy6 = (~(Xbzyx6 & Qo2iy6));
assign Qo2iy6 = (~(Yo2iy6 & Gp2iy6));
assign Gp2iy6 = (Op2iy6 & Wp2iy6);
assign Wp2iy6 = (Eq2iy6 & Mq2iy6);
assign Mq2iy6 = (~(Hyj7z6[0] & Rbk7z6[18]));
assign Eq2iy6 = (~(Hyj7z6[1] & Zlk7z6[18]));
assign Op2iy6 = (Uq2iy6 & Cr2iy6);
assign Cr2iy6 = (~(Hyj7z6[2] & Hwk7z6[18]));
assign Uq2iy6 = (~(Hyj7z6[3] & P6l7z6[18]));
assign Yo2iy6 = (Kr2iy6 & Sr2iy6);
assign Sr2iy6 = (As2iy6 & Is2iy6);
assign Is2iy6 = (~(Hyj7z6[4] & Xgl7z6[18]));
assign As2iy6 = (~(Hyj7z6[5] & Frl7z6[18]));
assign Kr2iy6 = (Qs2iy6 & Ys2iy6);
assign Ys2iy6 = (~(Hyj7z6[6] & N1m7z6[18]));
assign Qs2iy6 = (~(Hyj7z6[7] & Vbm7z6[18]));
assign Ao2iy6 = (~(Gt2iy6 & Ngqyx6));
assign Gt2iy6 = (~(Ot2iy6 & Wt2iy6));
assign Wt2iy6 = (Eu2iy6 & Mu2iy6);
assign Mu2iy6 = (Uu2iy6 & Cv2iy6);
assign Cv2iy6 = (Kv2iy6 & Sv2iy6);
assign Sv2iy6 = (~(Dpwyx6 & Fs0zx6));
assign Dpwyx6 = (Jmqyx6 & Tpyyx6);
assign Kv2iy6 = (Aw2iy6 & Ykthy6);
assign Aw2iy6 = (~(Iw2iy6 & Qw2iy6));
assign Iw2iy6 = (Voqyx6 & D2k7x6);
assign Uu2iy6 = (Yw2iy6 & Gx2iy6);
assign Gx2iy6 = (~(A0j7z6[20] & Xrqyx6));
assign Yw2iy6 = (~(H1j7z6[20] & Rqqyx6));
assign Eu2iy6 = (Ox2iy6 & Wx2iy6);
assign Wx2iy6 = (Ey2iy6 & My2iy6);
assign My2iy6 = (~(Wui7z6[20] & Lxqyx6));
assign Ey2iy6 = (~(Dri7z6[20] & Fwqyx6));
assign Ox2iy6 = (Uy2iy6 & Cz2iy6);
assign Cz2iy6 = (~(Bwi7z6[20] & Hzqyx6));
assign Uy2iy6 = (~(Svkhy6 & Pnb7z6[20]));
assign Ot2iy6 = (Kz2iy6 & Sz2iy6);
assign Sz2iy6 = (A03iy6 & I03iy6);
assign I03iy6 = (Q03iy6 & Y03iy6);
assign Y03iy6 = (~(Pzqyx6 & G5j7z6[52]));
assign Q03iy6 = (~(Jyqyx6 & G5j7z6[20]));
assign A03iy6 = (G13iy6 & O13iy6);
assign O13iy6 = (~(B2ryx6 & M6j7z6[52]));
assign G13iy6 = (~(J2ryx6 & M6j7z6[20]));
assign Kz2iy6 = (W13iy6 & E23iy6);
assign E23iy6 = (M23iy6 & U23iy6);
assign U23iy6 = (~(D1ryx6 & Ohj7z6[52]));
assign M23iy6 = (~(X3ryx6 & Ohj7z6[20]));
assign W13iy6 = (Whshy6 & C33iy6);
assign C33iy6 = (~(STCALIB[20] & F4ryx6));
assign Whshy6 = (Bqyyx6 & K33iy6);
assign U62iy6 = (S33iy6 & A43iy6);
assign A43iy6 = (I43iy6 & Q43iy6);
assign Q43iy6 = (~(Mqb7z6[4] & Lltyx6));
assign I43iy6 = (Y43iy6 & G53iy6);
assign G53iy6 = (~(Mm1nz6[4] & Pjtyx6));
assign Y43iy6 = (~(Yr1nz6[4] & Xjtyx6));
assign S33iy6 = (O53iy6 & W53iy6);
assign W53iy6 = (~(Ies7z6[20] & Tltyx6));
assign E62iy6 = (~(Zmoyx6 & Nqf7x6));
assign Nqf7x6 = (~(E63iy6 & M63iy6));
assign M63iy6 = (~(Cco7v6 & Aszhy6));
assign E63iy6 = (~(Tim7z6[20] & Yszhy6));
assign O52iy6 = (U63iy6 & C73iy6);
assign C73iy6 = (~(HRDATAS[20] & Ad47x6));
assign U63iy6 = (~(HRDATAD[20] & Mc47x6));
assign Y42iy6 = (~(Lpryx6 & Ckq7x6));
assign Zko7v6 = (~(K73iy6 & S73iy6));
assign S73iy6 = (~(Jexmz6[21] & K94iw6));
assign K73iy6 = (A83iy6 & I83iy6);
assign I83iy6 = (~(Lloyx6 & Xr57x6));
assign Xr57x6 = (~(Q83iy6 & Y83iy6));
assign Y83iy6 = (G93iy6 & O93iy6);
assign O93iy6 = (Bqoyx6 | Ttf7x6);
assign Ttf7x6 = (W93iy6 & Ea3iy6);
assign Ea3iy6 = (Ma3iy6 & Ua3iy6);
assign Ua3iy6 = (Cb3iy6 & Kb3iy6);
assign Kb3iy6 = (~(Xbzyx6 & Sb3iy6));
assign Sb3iy6 = (~(Ac3iy6 & Ic3iy6));
assign Ic3iy6 = (Qc3iy6 & Yc3iy6);
assign Yc3iy6 = (Gd3iy6 & Od3iy6);
assign Od3iy6 = (~(Hyj7z6[0] & Rbk7z6[19]));
assign Gd3iy6 = (~(Hyj7z6[1] & Zlk7z6[19]));
assign Qc3iy6 = (Wd3iy6 & Ee3iy6);
assign Ee3iy6 = (~(Hyj7z6[2] & Hwk7z6[19]));
assign Wd3iy6 = (~(Hyj7z6[3] & P6l7z6[19]));
assign Ac3iy6 = (Me3iy6 & Ue3iy6);
assign Ue3iy6 = (Cf3iy6 & Kf3iy6);
assign Kf3iy6 = (~(Hyj7z6[4] & Xgl7z6[19]));
assign Cf3iy6 = (~(Hyj7z6[5] & Frl7z6[19]));
assign Me3iy6 = (Sf3iy6 & Ag3iy6);
assign Ag3iy6 = (~(Hyj7z6[6] & N1m7z6[19]));
assign Sf3iy6 = (~(Hyj7z6[7] & Vbm7z6[19]));
assign Cb3iy6 = (Ig3iy6 & Qg3iy6);
assign Ig3iy6 = (~(Yg3iy6 & Feymz6[3]));
assign Ma3iy6 = (Gh3iy6 & Oh3iy6);
assign Oh3iy6 = (~(Wh3iy6 & Ngqyx6));
assign Wh3iy6 = (~(Ei3iy6 & Mi3iy6));
assign Mi3iy6 = (Ui3iy6 & Cj3iy6);
assign Cj3iy6 = (Kj3iy6 & Sj3iy6);
assign Sj3iy6 = (Ak3iy6 & Ik3iy6);
assign Ik3iy6 = (Qk3iy6 & Yk3iy6);
assign Yk3iy6 = (~(V40zx6 & Tcj7z6[0]));
assign Qk3iy6 = (U2vhy6 & Dhsyx6);
assign Ak3iy6 = (Gl3iy6 & Ol3iy6);
assign Ol3iy6 = (~(A0j7z6[21] & Xrqyx6));
assign Gl3iy6 = (~(H1j7z6[21] & Rqqyx6));
assign Kj3iy6 = (Wl3iy6 & Em3iy6);
assign Em3iy6 = (Mm3iy6 & Um3iy6);
assign Um3iy6 = (~(Wui7z6[21] & Lxqyx6));
assign Mm3iy6 = (~(Dri7z6[21] & Fwqyx6));
assign Wl3iy6 = (Cn3iy6 & Kn3iy6);
assign Kn3iy6 = (~(Bwi7z6[21] & Hzqyx6));
assign Cn3iy6 = (~(Ba0zx6 & Z8j7z6[0]));
assign Ui3iy6 = (Sn3iy6 & Ao3iy6);
assign Ao3iy6 = (Io3iy6 & Qo3iy6);
assign Qo3iy6 = (Yo3iy6 & Gp3iy6);
assign Gp3iy6 = (~(Svkhy6 & Pnb7z6[21]));
assign Yo3iy6 = (~(D90zx6 & Lgj7z6[186]));
assign Io3iy6 = (Op3iy6 & Wp3iy6);
assign Wp3iy6 = (~(Za0zx6 & Lgj7z6[174]));
assign Op3iy6 = (~(Hb0zx6 & Lgj7z6[162]));
assign Sn3iy6 = (Eq3iy6 & Mq3iy6);
assign Mq3iy6 = (Uq3iy6 & Cr3iy6);
assign Cr3iy6 = (~(Vc0zx6 & Lgj7z6[150]));
assign Uq3iy6 = (~(Dd0zx6 & Lgj7z6[138]));
assign Eq3iy6 = (Kr3iy6 & Sr3iy6);
assign Sr3iy6 = (~(Be0zx6 & Lgj7z6[126]));
assign Kr3iy6 = (~(Je0zx6 & Lgj7z6[114]));
assign Ei3iy6 = (As3iy6 & Is3iy6);
assign Is3iy6 = (Qs3iy6 & Ys3iy6);
assign Ys3iy6 = (Gt3iy6 & Ot3iy6);
assign Ot3iy6 = (Wt3iy6 & Eu3iy6);
assign Eu3iy6 = (~(Bi0zx6 & Lgj7z6[102]));
assign Wt3iy6 = (~(Ji0zx6 & Lgj7z6[90]));
assign Gt3iy6 = (Mu3iy6 & Uu3iy6);
assign Uu3iy6 = (~(Dh0zx6 & Lgj7z6[78]));
assign Mu3iy6 = (~(Hj0zx6 & Lgj7z6[66]));
assign Qs3iy6 = (Cv3iy6 & Kv3iy6);
assign Kv3iy6 = (Sv3iy6 & Aw3iy6);
assign Aw3iy6 = (~(Pj0zx6 & Lgj7z6[54]));
assign Sv3iy6 = (~(Dl0zx6 & Lgj7z6[42]));
assign Cv3iy6 = (Iw3iy6 & Qw3iy6);
assign Qw3iy6 = (~(Ll0zx6 & Lgj7z6[30]));
assign Iw3iy6 = (~(Jm0zx6 & Lgj7z6[18]));
assign As3iy6 = (Yw3iy6 & Gx3iy6);
assign Gx3iy6 = (Ox3iy6 & Wx3iy6);
assign Wx3iy6 = (Ey3iy6 & My3iy6);
assign My3iy6 = (~(Rm0zx6 & Lgj7z6[6]));
assign Ey3iy6 = (~(Pzqyx6 & G5j7z6[53]));
assign Ox3iy6 = (Uy3iy6 & Cz3iy6);
assign Cz3iy6 = (~(Jyqyx6 & G5j7z6[21]));
assign Uy3iy6 = (~(B2ryx6 & M6j7z6[53]));
assign Yw3iy6 = (Kz3iy6 & Sz3iy6);
assign Sz3iy6 = (A04iy6 & I04iy6);
assign I04iy6 = (~(J2ryx6 & M6j7z6[21]));
assign A04iy6 = (~(D1ryx6 & Ohj7z6[53]));
assign Kz3iy6 = (Q04iy6 & Y04iy6);
assign Y04iy6 = (~(X3ryx6 & Ohj7z6[21]));
assign Q04iy6 = (~(STCALIB[21] & F4ryx6));
assign Gh3iy6 = (G14iy6 & O14iy6);
assign O14iy6 = (~(Rmzyx6 & W14iy6));
assign W14iy6 = (~(E24iy6 & M24iy6));
assign M24iy6 = (U24iy6 & C34iy6);
assign C34iy6 = (K34iy6 & S34iy6);
assign S34iy6 = (~(Hyj7z6[3] & Tnciw6));
assign K34iy6 = (~(Hyj7z6[2] & Mnciw6));
assign U24iy6 = (A44iy6 & I44iy6);
assign I44iy6 = (~(Hyj7z6[1] & Fnciw6));
assign A44iy6 = (~(Hyj7z6[5] & Aociw6));
assign E24iy6 = (Q44iy6 & Y44iy6);
assign Y44iy6 = (G54iy6 & O54iy6);
assign O54iy6 = (~(Hyj7z6[6] & Oociw6));
assign G54iy6 = (~(Hyj7z6[7] & Cpciw6));
assign Q44iy6 = (W54iy6 & E64iy6);
assign E64iy6 = (~(Hyj7z6[0] & Dfk7z6[21]));
assign W54iy6 = (~(Hyj7z6[4] & Jkl7z6[21]));
assign G14iy6 = (~(Klo7z6[2] & M64iy6));
assign M64iy6 = (~(U64iy6 & C74iy6));
assign C74iy6 = (K74iy6 & S74iy6);
assign S74iy6 = (A84iy6 & I84iy6);
assign I84iy6 = (~(Fmset6 & S4kiw6));
assign A84iy6 = (Q84iy6 & Y84iy6);
assign Y84iy6 = (~(Nqo7z6[19] & M8kiw6));
assign Q84iy6 = (~(Fpo7z6[19] & H9kiw6));
assign K74iy6 = (G94iy6 & O94iy6);
assign O94iy6 = (~(Ouo7z6[19] & K7kiw6));
assign G94iy6 = (~(Hxo7z6[19] & W6kiw6));
assign U64iy6 = (W94iy6 & Ea4iy6);
assign Ea4iy6 = (Ma4iy6 & Ua4iy6);
assign Ua4iy6 = (~(Vro7z6[19] & Y7kiw6));
assign Ma4iy6 = (~(T2p7z6[21] & U5kiw6));
assign W94iy6 = (Cb4iy6 & Kb4iy6);
assign Kb4iy6 = (~(W3p7z6[21] & G5kiw6));
assign Cb4iy6 = (~(A0p7z6[19] & I6kiw6));
assign W93iy6 = (Sb4iy6 & Ac4iy6);
assign Ac4iy6 = (Ic4iy6 & Qc4iy6);
assign Qc4iy6 = (~(Yr1nz6[5] & Xjtyx6));
assign Ic4iy6 = (Yc4iy6 & Gd4iy6);
assign Gd4iy6 = (~(Klo7z6[1] & Od4iy6));
assign Od4iy6 = (~(Wd4iy6 & Ee4iy6));
assign Ee4iy6 = (Me4iy6 & Ue4iy6);
assign Ue4iy6 = (Cf4iy6 & Ravyx6);
assign Cf4iy6 = (~(T9tyx6 & Wp77z6));
assign Me4iy6 = (Kf4iy6 & Sf4iy6);
assign Sf4iy6 = (~(Xkq7z6[21] & B6qyx6));
assign Kf4iy6 = (~(Bqp7z6[21] & D5qyx6));
assign Wd4iy6 = (Ag4iy6 & Ig4iy6);
assign Ig4iy6 = (Qg4iy6 & Yg4iy6);
assign Yg4iy6 = (~(E6p7z6[21] & L9qyx6));
assign Qg4iy6 = (~(B2q7z6[21] & Fcqyx6));
assign Ag4iy6 = (Gh4iy6 & Oh4iy6);
assign Oh4iy6 = (~(Mkp7z6[21] & Tdqyx6));
assign Gh4iy6 = (~(Hfqyx6 & U9p7z6[21]));
assign Yc4iy6 = (~(Mm1nz6[5] & Pjtyx6));
assign Sb4iy6 = (Wh4iy6 & Ei4iy6);
assign Ei4iy6 = (~(Mqb7z6[5] & Lltyx6));
assign Wh4iy6 = (~(Ies7z6[21] & Tltyx6));
assign G93iy6 = (~(Zmoyx6 & Auf7x6));
assign Auf7x6 = (~(Mi4iy6 & Ui4iy6));
assign Ui4iy6 = (~(Aszhy6 & G9a7z6));
assign G9a7z6 = (~(Cj4iy6 & Kj4iy6));
assign Kj4iy6 = (~(HRDATAD[21] & Qln7z6[0]));
assign Cj4iy6 = (~(HRDATAS[21] & Qln7z6[1]));
assign Mi4iy6 = (~(Tim7z6[21] & Yszhy6));
assign Q83iy6 = (Sj4iy6 & Ak4iy6);
assign Ak4iy6 = (~(HRDATAS[21] & Ad47x6));
assign Sj4iy6 = (~(HRDATAD[21] & Mc47x6));
assign A83iy6 = (~(Lpryx6 & Mpq7x6));
assign Sko7v6 = (~(Ik4iy6 & Qk4iy6));
assign Qk4iy6 = (~(Jexmz6[22] & K94iw6));
assign Ik4iy6 = (Yk4iy6 & Gl4iy6);
assign Gl4iy6 = (~(Lloyx6 & Um57x6));
assign Um57x6 = (~(Ol4iy6 & Wl4iy6));
assign Wl4iy6 = (Em4iy6 & Mm4iy6);
assign Mm4iy6 = (Bqoyx6 | Gxf7x6);
assign Gxf7x6 = (Um4iy6 & Cn4iy6);
assign Cn4iy6 = (Kn4iy6 & Sn4iy6);
assign Sn4iy6 = (Ao4iy6 & Io4iy6);
assign Io4iy6 = (~(Qo4iy6 & U2jhy6));
assign Qo4iy6 = (Yo4iy6 & K3jhy6);
assign Yo4iy6 = (~(Gp4iy6 & Op4iy6));
assign Op4iy6 = (Wp4iy6 & Eq4iy6);
assign Eq4iy6 = (Mq4iy6 & Uq4iy6);
assign Uq4iy6 = (~(Hyj7z6[3] & Xpciw6));
assign Mq4iy6 = (~(Hyj7z6[2] & Qpciw6));
assign Wp4iy6 = (Cr4iy6 & Kr4iy6);
assign Kr4iy6 = (~(Hyj7z6[1] & Jpciw6));
assign Cr4iy6 = (~(Hyj7z6[5] & Eqciw6));
assign Gp4iy6 = (Sr4iy6 & As4iy6);
assign As4iy6 = (Is4iy6 & Qs4iy6);
assign Qs4iy6 = (~(Hyj7z6[6] & Lqciw6));
assign Is4iy6 = (~(Hyj7z6[7] & Sqciw6));
assign Sr4iy6 = (Ys4iy6 & Gt4iy6);
assign Gt4iy6 = (~(Hyj7z6[0] & Dfk7z6[22]));
assign Ys4iy6 = (~(Hyj7z6[4] & Jkl7z6[22]));
assign Ao4iy6 = (Gd2iy6 & Qg3iy6);
assign Kn4iy6 = (Ot4iy6 & Wt4iy6);
assign Wt4iy6 = (~(Eu4iy6 & Ngqyx6));
assign Eu4iy6 = (~(Mu4iy6 & Uu4iy6));
assign Uu4iy6 = (Cv4iy6 & Kv4iy6);
assign Kv4iy6 = (Sv4iy6 & Aw4iy6);
assign Aw4iy6 = (Iw4iy6 & Qw4iy6);
assign Qw4iy6 = (Yw4iy6 & Gx4iy6);
assign Gx4iy6 = (~(Dxqyx6 & Ox4iy6));
assign Ox4iy6 = (~(Wx4iy6 & Ey4iy6));
assign Ey4iy6 = (My4iy6 & Uy4iy6);
assign Uy4iy6 = (Cz4iy6 & Kz4iy6);
assign Kz4iy6 = (Sz4iy6 & A05iy6);
assign A05iy6 = (I05iy6 & Q05iy6);
assign Q05iy6 = (E4eov6 & X3eov6);
assign X3eov6 = (!M6j7z6[9]);
assign E4eov6 = (!M6j7z6[8]);
assign I05iy6 = (Zpeov6 & Ageov6);
assign Ageov6 = (!M6j7z6[7]);
assign Zpeov6 = (!M6j7z6[6]);
assign Sz4iy6 = (Y05iy6 & G15iy6);
assign G15iy6 = (Rfdov6 & Sweov6);
assign Sweov6 = (!M6j7z6[63]);
assign Rfdov6 = (!M6j7z6[62]);
assign Y05iy6 = (Tgdov6 & Wedov6);
assign Wedov6 = (!M6j7z6[61]);
assign Tgdov6 = (!M6j7z6[60]);
assign Cz4iy6 = (O15iy6 & W15iy6);
assign W15iy6 = (E25iy6 & M25iy6);
assign M25iy6 = (Gkdov6 & Yeeov6);
assign Yeeov6 = (!M6j7z6[5]);
assign Gkdov6 = (!M6j7z6[59]);
assign E25iy6 = (Fndov6 & Nkdov6);
assign Nkdov6 = (!M6j7z6[58]);
assign Fndov6 = (!M6j7z6[57]);
assign O15iy6 = (U25iy6 & C35iy6);
assign C35iy6 = (Ahdov6 & Mndov6);
assign Mndov6 = (!M6j7z6[56]);
assign Ahdov6 = (!M6j7z6[55]);
assign U25iy6 = (Ljdov6 & Ejdov6);
assign Ejdov6 = (!M6j7z6[54]);
assign Ljdov6 = (!M6j7z6[53]);
assign My4iy6 = (K35iy6 & S35iy6);
assign S35iy6 = (A45iy6 & I45iy6);
assign I45iy6 = (Q45iy6 & Y45iy6);
assign Y45iy6 = (A9eov6 & Jidov6);
assign Jidov6 = (!M6j7z6[52]);
assign A9eov6 = (!M6j7z6[51]);
assign Q45iy6 = (Uqeov6 & Lieov6);
assign Lieov6 = (!M6j7z6[50]);
assign Uqeov6 = (!M6j7z6[4]);
assign A45iy6 = (G55iy6 & O55iy6);
assign O55iy6 = (Sieov6 & H9eov6);
assign H9eov6 = (!M6j7z6[49]);
assign Sieov6 = (!M6j7z6[48]);
assign G55iy6 = (Kmdov6 & Aueov6);
assign Aueov6 = (!M6j7z6[47]);
assign Kmdov6 = (!M6j7z6[46]);
assign K35iy6 = (W55iy6 & E65iy6);
assign E65iy6 = (M65iy6 & U65iy6);
assign U65iy6 = (Oodov6 & Hodov6);
assign Hodov6 = (!M6j7z6[45]);
assign Oodov6 = (!M6j7z6[44]);
assign M65iy6 = (Eqdov6 & Xpdov6);
assign Xpdov6 = (!M6j7z6[43]);
assign Eqdov6 = (!M6j7z6[42]);
assign W55iy6 = (C75iy6 & K75iy6);
assign K75iy6 = (Grdov6 & Zqdov6);
assign Zqdov6 = (!M6j7z6[41]);
assign Grdov6 = (!M6j7z6[40]);
assign C75iy6 = (F8eov6 & Vgeov6);
assign Vgeov6 = (!M6j7z6[3]);
assign F8eov6 = (!M6j7z6[39]);
assign Wx4iy6 = (S75iy6 & A85iy6);
assign A85iy6 = (I85iy6 & Q85iy6);
assign Q85iy6 = (Y85iy6 & G95iy6);
assign G95iy6 = (O95iy6 & W95iy6);
assign W95iy6 = (Caeov6 & Njeov6);
assign Njeov6 = (!M6j7z6[38]);
assign Caeov6 = (!M6j7z6[37]);
assign O95iy6 = (Jaeov6 & Ujeov6);
assign Ujeov6 = (!M6j7z6[36]);
assign Jaeov6 = (!M6j7z6[35]);
assign Y85iy6 = (Ea5iy6 & Ma5iy6);
assign Ma5iy6 = (Sbeov6 & Aneov6);
assign Aneov6 = (!M6j7z6[34]);
assign Sbeov6 = (!M6j7z6[33]);
assign Ea5iy6 = (Mudov6 & Hneov6);
assign Hneov6 = (!M6j7z6[32]);
assign Mudov6 = (!M6j7z6[31]);
assign I85iy6 = (Ua5iy6 & Cb5iy6);
assign Cb5iy6 = (Kb5iy6 & Sb5iy6);
assign Sb5iy6 = (Breov6 & Tudov6);
assign Tudov6 = (!M6j7z6[30]);
assign Breov6 = (!M6j7z6[2]);
assign Kb5iy6 = (Ovdov6 & Rtdov6);
assign Rtdov6 = (!M6j7z6[29]);
assign Ovdov6 = (!M6j7z6[28]);
assign Ua5iy6 = (Ac5iy6 & Ic5iy6);
assign Ic5iy6 = (Exdov6 & Vvdov6);
assign Vvdov6 = (!M6j7z6[27]);
assign Exdov6 = (!M6j7z6[26]);
assign Ac5iy6 = (Gydov6 & Lxdov6);
assign Lxdov6 = (!M6j7z6[25]);
assign Gydov6 = (!M6j7z6[24]);
assign S75iy6 = (Qc5iy6 & Yc5iy6);
assign Yc5iy6 = (Gd5iy6 & Od5iy6);
assign Od5iy6 = (Wd5iy6 & Ee5iy6);
assign Ee5iy6 = (Fmeov6 & Zbeov6);
assign Zbeov6 = (!M6j7z6[23]);
assign Fmeov6 = (!M6j7z6[22]);
assign Wd5iy6 = (Coeov6 & Uceov6);
assign Uceov6 = (!M6j7z6[21]);
assign Coeov6 = (!M6j7z6[20]);
assign Gd5iy6 = (Me5iy6 & Ue5iy6);
assign Ue5iy6 = (Bdeov6 & Cheov6);
assign Cheov6 = (!M6j7z6[1]);
assign Bdeov6 = (!M6j7z6[19]);
assign Me5iy6 = (Tfeov6 & Joeov6);
assign Joeov6 = (!M6j7z6[18]);
assign Tfeov6 = (!M6j7z6[17]);
assign Qc5iy6 = (Cf5iy6 & Kf5iy6);
assign Kf5iy6 = (Sf5iy6 & Ag5iy6);
assign Ag5iy6 = (Nydov6 & Speov6);
assign Speov6 = (!M6j7z6[16]);
assign Nydov6 = (!M6j7z6[15]);
assign Sf5iy6 = (M1eov6 & F1eov6);
assign F1eov6 = (!M6j7z6[14]);
assign M1eov6 = (!M6j7z6[13]);
assign Cf5iy6 = (Ig5iy6 & Qg5iy6);
assign Qg5iy6 = (H2eov6 & K0eov6);
assign K0eov6 = (!M6j7z6[12]);
assign H2eov6 = (!M6j7z6[11]);
assign Ig5iy6 = (Tteov6 & O2eov6);
assign O2eov6 = (!M6j7z6[10]);
assign Tteov6 = (!M6j7z6[0]);
assign Yw4iy6 = (~(V40zx6 & Tcj7z6[1]));
assign Iw4iy6 = (Yg5iy6 & Gh5iy6);
assign Gh5iy6 = (~(A0j7z6[22] & Xrqyx6));
assign Yg5iy6 = (~(H1j7z6[22] & Rqqyx6));
assign Sv4iy6 = (Oh5iy6 & Wh5iy6);
assign Wh5iy6 = (Ei5iy6 & Mi5iy6);
assign Mi5iy6 = (~(Wui7z6[22] & Lxqyx6));
assign Ei5iy6 = (~(Dri7z6[22] & Fwqyx6));
assign Oh5iy6 = (Ui5iy6 & Cj5iy6);
assign Cj5iy6 = (~(Bwi7z6[22] & Hzqyx6));
assign Ui5iy6 = (~(Ba0zx6 & Z8j7z6[1]));
assign Cv4iy6 = (Kj5iy6 & Sj5iy6);
assign Sj5iy6 = (Ak5iy6 & Ik5iy6);
assign Ik5iy6 = (Qk5iy6 & Yk5iy6);
assign Yk5iy6 = (~(Svkhy6 & Pnb7z6[22]));
assign Qk5iy6 = (~(D90zx6 & Lgj7z6[187]));
assign Ak5iy6 = (Gl5iy6 & Ol5iy6);
assign Ol5iy6 = (~(Za0zx6 & Lgj7z6[175]));
assign Gl5iy6 = (~(Hb0zx6 & Lgj7z6[163]));
assign Kj5iy6 = (Wl5iy6 & Em5iy6);
assign Em5iy6 = (Mm5iy6 & Um5iy6);
assign Um5iy6 = (~(Vc0zx6 & Lgj7z6[151]));
assign Mm5iy6 = (~(Dd0zx6 & Lgj7z6[139]));
assign Wl5iy6 = (Cn5iy6 & Kn5iy6);
assign Kn5iy6 = (~(Be0zx6 & Lgj7z6[127]));
assign Cn5iy6 = (~(Je0zx6 & Lgj7z6[115]));
assign Mu4iy6 = (Sn5iy6 & Ao5iy6);
assign Ao5iy6 = (Io5iy6 & Qo5iy6);
assign Qo5iy6 = (Yo5iy6 & Gp5iy6);
assign Gp5iy6 = (Op5iy6 & Wp5iy6);
assign Wp5iy6 = (~(Bi0zx6 & Lgj7z6[103]));
assign Op5iy6 = (~(Ji0zx6 & Lgj7z6[91]));
assign Yo5iy6 = (Eq5iy6 & Mq5iy6);
assign Mq5iy6 = (~(Dh0zx6 & Lgj7z6[79]));
assign Eq5iy6 = (~(Hj0zx6 & Lgj7z6[67]));
assign Io5iy6 = (Uq5iy6 & Cr5iy6);
assign Cr5iy6 = (Kr5iy6 & Sr5iy6);
assign Sr5iy6 = (~(Pj0zx6 & Lgj7z6[55]));
assign Kr5iy6 = (~(Dl0zx6 & Lgj7z6[43]));
assign Uq5iy6 = (As5iy6 & Is5iy6);
assign Is5iy6 = (~(Ll0zx6 & Lgj7z6[31]));
assign As5iy6 = (~(Jm0zx6 & Lgj7z6[19]));
assign Sn5iy6 = (Qs5iy6 & Ys5iy6);
assign Ys5iy6 = (Gt5iy6 & Ot5iy6);
assign Ot5iy6 = (Wt5iy6 & Eu5iy6);
assign Eu5iy6 = (~(Rm0zx6 & Lgj7z6[7]));
assign Wt5iy6 = (~(Pzqyx6 & G5j7z6[54]));
assign Gt5iy6 = (Mu5iy6 & Uu5iy6);
assign Uu5iy6 = (~(Jyqyx6 & G5j7z6[22]));
assign Mu5iy6 = (~(B2ryx6 & M6j7z6[54]));
assign Qs5iy6 = (Cv5iy6 & Kv5iy6);
assign Kv5iy6 = (Sv5iy6 & Aw5iy6);
assign Aw5iy6 = (~(J2ryx6 & M6j7z6[22]));
assign Sv5iy6 = (~(D1ryx6 & Ohj7z6[54]));
assign Cv5iy6 = (Iw5iy6 & Qw5iy6);
assign Qw5iy6 = (~(X3ryx6 & Ohj7z6[22]));
assign Iw5iy6 = (~(STCALIB[22] & F4ryx6));
assign Ot4iy6 = (~(Klo7z6[2] & Yw5iy6));
assign Yw5iy6 = (~(Gx5iy6 & Ox5iy6));
assign Ox5iy6 = (Wx5iy6 & Ey5iy6);
assign Ey5iy6 = (My5iy6 & Uy5iy6);
assign Uy5iy6 = (~(Ekset6 & S4kiw6));
assign My5iy6 = (Cz5iy6 & Kz5iy6);
assign Kz5iy6 = (~(Nqo7z6[20] & M8kiw6));
assign Cz5iy6 = (~(Fpo7z6[20] & H9kiw6));
assign Wx5iy6 = (Sz5iy6 & A06iy6);
assign A06iy6 = (~(Ouo7z6[20] & K7kiw6));
assign Sz5iy6 = (~(Hxo7z6[20] & W6kiw6));
assign Gx5iy6 = (I06iy6 & Q06iy6);
assign Q06iy6 = (Y06iy6 & G16iy6);
assign G16iy6 = (~(Vro7z6[20] & Y7kiw6));
assign Y06iy6 = (~(T2p7z6[22] & U5kiw6));
assign I06iy6 = (O16iy6 & W16iy6);
assign W16iy6 = (~(W3p7z6[22] & G5kiw6));
assign O16iy6 = (~(A0p7z6[20] & I6kiw6));
assign Um4iy6 = (E26iy6 & M26iy6);
assign M26iy6 = (U26iy6 & C36iy6);
assign C36iy6 = (~(Yr1nz6[6] & Xjtyx6));
assign U26iy6 = (K36iy6 & S36iy6);
assign S36iy6 = (~(Klo7z6[1] & A46iy6));
assign A46iy6 = (~(I46iy6 & Q46iy6));
assign Q46iy6 = (Y46iy6 & G56iy6);
assign G56iy6 = (O56iy6 & Ravyx6);
assign O56iy6 = (~(T9tyx6 & Op77z6));
assign Y46iy6 = (W56iy6 & E66iy6);
assign E66iy6 = (~(Xkq7z6[22] & B6qyx6));
assign W56iy6 = (~(Bqp7z6[22] & D5qyx6));
assign I46iy6 = (M66iy6 & U66iy6);
assign U66iy6 = (C76iy6 & K76iy6);
assign K76iy6 = (~(E6p7z6[22] & L9qyx6));
assign C76iy6 = (~(B2q7z6[22] & Fcqyx6));
assign M66iy6 = (S76iy6 & A86iy6);
assign A86iy6 = (~(Mkp7z6[22] & Tdqyx6));
assign S76iy6 = (~(Hfqyx6 & U9p7z6[22]));
assign K36iy6 = (~(Mm1nz6[6] & Pjtyx6));
assign E26iy6 = (I86iy6 & Q86iy6);
assign Q86iy6 = (~(Mqb7z6[6] & Lltyx6));
assign I86iy6 = (~(Ies7z6[22] & Tltyx6));
assign Em4iy6 = (~(Zmoyx6 & Nxf7x6));
assign Nxf7x6 = (~(Y86iy6 & G96iy6));
assign G96iy6 = (~(Aszhy6 & Y8a7z6));
assign Y8a7z6 = (~(O96iy6 & W96iy6));
assign W96iy6 = (~(HRDATAD[22] & Qln7z6[0]));
assign O96iy6 = (~(HRDATAS[22] & Qln7z6[1]));
assign Y86iy6 = (~(Tim7z6[22] & Yszhy6));
assign Ol4iy6 = (Ea6iy6 & Ma6iy6);
assign Ma6iy6 = (~(HRDATAS[22] & Ad47x6));
assign Ea6iy6 = (~(HRDATAD[22] & Mc47x6));
assign Yk4iy6 = (~(Lpryx6 & Wuq7x6));
assign Lko7v6 = (~(Ua6iy6 & Cb6iy6));
assign Cb6iy6 = (~(Jexmz6[23] & K94iw6));
assign Ua6iy6 = (Kb6iy6 & Sb6iy6);
assign Sb6iy6 = (~(Lloyx6 & Rh57x6));
assign Rh57x6 = (~(Ac6iy6 & Ic6iy6));
assign Ic6iy6 = (Qc6iy6 & Yc6iy6);
assign Yc6iy6 = (Bqoyx6 | T0g7x6);
assign T0g7x6 = (Gd6iy6 & Od6iy6);
assign Od6iy6 = (Wd6iy6 & Ee6iy6);
assign Ee6iy6 = (Me6iy6 & Ue6iy6);
assign Ue6iy6 = (~(Lltyx6 & Tp3yx6));
assign Tp3yx6 = (~(Cf6iy6 & Kf6iy6));
assign Kf6iy6 = (~(La6ft6 | I96ft6));
assign Cf6iy6 = (Pf5ov6 & N0hyx6);
assign N0hyx6 = (!Zygyx6);
assign Zygyx6 = (~(Sf6iy6 & Ag6iy6));
assign Ag6iy6 = (Ig6iy6 & Tw37v6);
assign Ig6iy6 = (Ly37v6 & D047v6);
assign Sf6iy6 = (~(D1gyx6 | Thfyx6));
assign Thfyx6 = (!Bv37v6);
assign D1gyx6 = (!Jt37v6);
assign Pf5ov6 = (!X3gyx6);
assign X3gyx6 = (~(Rqhyx6 & Dthyx6));
assign Dthyx6 = (C55ov6 & Vcgyx6);
assign Vcgyx6 = (!Fbxmz6[3]);
assign C55ov6 = (!Fbxmz6[2]);
assign Rqhyx6 = (Ncgyx6 & M35ov6);
assign M35ov6 = (!Fbxmz6[1]);
assign Ncgyx6 = (!Fbxmz6[0]);
assign Lltyx6 = (Qg6iy6 & Klo7z6[0]);
assign Qg6iy6 = (Zfs7z6[7] & Hfryx6);
assign Me6iy6 = (Yg6iy6 & Gh6iy6);
assign Gh6iy6 = (~(Oh6iy6 & U2jhy6));
assign Oh6iy6 = (Wh6iy6 & K3jhy6);
assign Wh6iy6 = (~(Ei6iy6 & Mi6iy6));
assign Mi6iy6 = (Ui6iy6 & Cj6iy6);
assign Cj6iy6 = (Kj6iy6 & Sj6iy6);
assign Sj6iy6 = (~(Hyj7z6[1] & Grciw6));
assign Kj6iy6 = (~(Hyj7z6[2] & Nrciw6));
assign Ui6iy6 = (Ak6iy6 & Ik6iy6);
assign Ik6iy6 = (~(Hyj7z6[3] & Urciw6));
assign Ak6iy6 = (~(Hyj7z6[5] & Bsciw6));
assign Ei6iy6 = (Qk6iy6 & Yk6iy6);
assign Yk6iy6 = (Gl6iy6 & Ol6iy6);
assign Ol6iy6 = (~(Hyj7z6[6] & Isciw6));
assign Gl6iy6 = (~(Hyj7z6[7] & Psciw6));
assign Qk6iy6 = (Wl6iy6 & Em6iy6);
assign Em6iy6 = (~(Hyj7z6[0] & Dfk7z6[23]));
assign Wl6iy6 = (~(Hyj7z6[4] & Jkl7z6[23]));
assign Yg6iy6 = (~(Klo7z6[1] & Mm6iy6));
assign Mm6iy6 = (~(Um6iy6 & Cn6iy6));
assign Cn6iy6 = (Kn6iy6 & Sn6iy6);
assign Sn6iy6 = (~(B2q7z6[23] & Fcqyx6));
assign Kn6iy6 = (Ao6iy6 & Io6iy6);
assign Io6iy6 = (~(Bqp7z6[23] & D5qyx6));
assign Ao6iy6 = (~(E6p7z6[23] & L9qyx6));
assign Um6iy6 = (Qo6iy6 & Yo6iy6);
assign Yo6iy6 = (~(Mkp7z6[23] & Tdqyx6));
assign Qo6iy6 = (~(Hfqyx6 & U9p7z6[23]));
assign Wd6iy6 = (Gp6iy6 & Op6iy6);
assign Op6iy6 = (~(Mm1nz6[7] & Pjtyx6));
assign Gp6iy6 = (~(Yr1nz6[7] & Xjtyx6));
assign Gd6iy6 = (Wp6iy6 & Eq6iy6);
assign Eq6iy6 = (Mq6iy6 & Uq6iy6);
assign Uq6iy6 = (~(Cr6iy6 & Gp77z6));
assign Mq6iy6 = (Kr6iy6 & Sr6iy6);
assign Sr6iy6 = (~(As6iy6 & Ngqyx6));
assign As6iy6 = (~(Is6iy6 & Qs6iy6));
assign Qs6iy6 = (Ys6iy6 & Gt6iy6);
assign Gt6iy6 = (Ot6iy6 & Wt6iy6);
assign Wt6iy6 = (Eu6iy6 & Mu6iy6);
assign Mu6iy6 = (Uu6iy6 & Cv6iy6);
assign Cv6iy6 = (~(Kv6iy6 & Dxqyx6));
assign Kv6iy6 = (Tnzdt6 & F02nv6);
assign Uu6iy6 = (~(V40zx6 & Tcj7z6[2]));
assign V40zx6 = (~(Knohy6 | Zyuyx6));
assign Eu6iy6 = (Sv6iy6 & Aw6iy6);
assign Aw6iy6 = (~(A0j7z6[23] & Xrqyx6));
assign Xrqyx6 = (~(Lxuyx6 | Zyuyx6));
assign Sv6iy6 = (~(H1j7z6[23] & Rqqyx6));
assign Rqqyx6 = (~(Tlqyx6 | Lxuyx6));
assign Ot6iy6 = (Iw6iy6 & Qw6iy6);
assign Qw6iy6 = (Yw6iy6 & Gx6iy6);
assign Gx6iy6 = (~(Wui7z6[23] & Lxqyx6));
assign Yw6iy6 = (~(Dri7z6[23] & Fwqyx6));
assign Iw6iy6 = (Ox6iy6 & Wx6iy6);
assign Wx6iy6 = (~(Bwi7z6[23] & Hzqyx6));
assign Ox6iy6 = (~(Ba0zx6 & Z8j7z6[2]));
assign Ys6iy6 = (Ey6iy6 & My6iy6);
assign My6iy6 = (Uy6iy6 & Cz6iy6);
assign Cz6iy6 = (Kz6iy6 & Sz6iy6);
assign Sz6iy6 = (~(Svkhy6 & Pnb7z6[23]));
assign Kz6iy6 = (~(D90zx6 & Lgj7z6[188]));
assign Uy6iy6 = (A07iy6 & I07iy6);
assign I07iy6 = (~(Za0zx6 & Lgj7z6[176]));
assign A07iy6 = (~(Hb0zx6 & Lgj7z6[164]));
assign Ey6iy6 = (Q07iy6 & Y07iy6);
assign Y07iy6 = (G17iy6 & O17iy6);
assign O17iy6 = (~(Vc0zx6 & Lgj7z6[152]));
assign G17iy6 = (~(Dd0zx6 & Lgj7z6[140]));
assign Q07iy6 = (W17iy6 & E27iy6);
assign E27iy6 = (~(Be0zx6 & Lgj7z6[128]));
assign W17iy6 = (~(Je0zx6 & Lgj7z6[116]));
assign Is6iy6 = (M27iy6 & U27iy6);
assign U27iy6 = (C37iy6 & K37iy6);
assign K37iy6 = (S37iy6 & A47iy6);
assign A47iy6 = (I47iy6 & Q47iy6);
assign Q47iy6 = (~(Bi0zx6 & Lgj7z6[104]));
assign I47iy6 = (~(Ji0zx6 & Lgj7z6[92]));
assign S37iy6 = (Y47iy6 & G57iy6);
assign G57iy6 = (~(Dh0zx6 & Lgj7z6[80]));
assign Y47iy6 = (~(Hj0zx6 & Lgj7z6[68]));
assign C37iy6 = (O57iy6 & W57iy6);
assign W57iy6 = (E67iy6 & M67iy6);
assign M67iy6 = (~(Pj0zx6 & Lgj7z6[56]));
assign E67iy6 = (~(Dl0zx6 & Lgj7z6[44]));
assign O57iy6 = (U67iy6 & C77iy6);
assign C77iy6 = (~(Ll0zx6 & Lgj7z6[32]));
assign U67iy6 = (~(Jm0zx6 & Lgj7z6[20]));
assign M27iy6 = (K77iy6 & S77iy6);
assign S77iy6 = (A87iy6 & I87iy6);
assign I87iy6 = (Q87iy6 & Y87iy6);
assign Y87iy6 = (~(Rm0zx6 & Lgj7z6[8]));
assign Q87iy6 = (~(Pzqyx6 & G5j7z6[55]));
assign A87iy6 = (G97iy6 & O97iy6);
assign O97iy6 = (~(Jyqyx6 & G5j7z6[23]));
assign G97iy6 = (~(B2ryx6 & M6j7z6[55]));
assign K77iy6 = (W97iy6 & Ea7iy6);
assign Ea7iy6 = (Ma7iy6 & Ua7iy6);
assign Ua7iy6 = (~(J2ryx6 & M6j7z6[23]));
assign Ma7iy6 = (~(D1ryx6 & Ohj7z6[55]));
assign W97iy6 = (Cb7iy6 & Kb7iy6);
assign Kb7iy6 = (~(X3ryx6 & Ohj7z6[23]));
assign Cb7iy6 = (~(STCALIB[23] & F4ryx6));
assign Kr6iy6 = (~(Klo7z6[2] & Sb7iy6));
assign Sb7iy6 = (~(Ac7iy6 & Ic7iy6));
assign Ic7iy6 = (Qc7iy6 & Yc7iy6);
assign Yc7iy6 = (Gd7iy6 & Od7iy6);
assign Od7iy6 = (~(Diset6 & S4kiw6));
assign Gd7iy6 = (Wd7iy6 & Ee7iy6);
assign Ee7iy6 = (~(Nqo7z6[21] & M8kiw6));
assign Wd7iy6 = (~(Fpo7z6[21] & H9kiw6));
assign Qc7iy6 = (Me7iy6 & Ue7iy6);
assign Ue7iy6 = (~(Ouo7z6[21] & K7kiw6));
assign Me7iy6 = (~(Hxo7z6[21] & W6kiw6));
assign Ac7iy6 = (Cf7iy6 & Kf7iy6);
assign Kf7iy6 = (Sf7iy6 & Ag7iy6);
assign Ag7iy6 = (~(Vro7z6[21] & Y7kiw6));
assign Sf7iy6 = (~(T2p7z6[23] & U5kiw6));
assign Cf7iy6 = (Ig7iy6 & Qg7iy6);
assign Qg7iy6 = (~(W3p7z6[23] & G5kiw6));
assign Ig7iy6 = (~(A0p7z6[21] & I6kiw6));
assign Wp6iy6 = (Yg7iy6 & Gh7iy6);
assign Gh7iy6 = (~(Ies7z6[23] & Tltyx6));
assign Qc6iy6 = (~(HRDATAS[23] & Ad47x6));
assign Ac6iy6 = (Oh7iy6 & Wh7iy6);
assign Wh7iy6 = (~(HRDATAD[23] & Mc47x6));
assign Oh7iy6 = (~(Zmoyx6 & A1g7x6));
assign A1g7x6 = (~(Ei7iy6 & Mi7iy6));
assign Mi7iy6 = (~(Aszhy6 & Q8a7z6));
assign Q8a7z6 = (~(Ui7iy6 & Cj7iy6));
assign Cj7iy6 = (~(HRDATAD[23] & Qln7z6[0]));
assign Ui7iy6 = (~(HRDATAS[23] & Qln7z6[1]));
assign Ei7iy6 = (~(Tim7z6[23] & Yszhy6));
assign Kb6iy6 = (~(Lpryx6 & Xzp7x6));
assign Eko7v6 = (~(Kj7iy6 & Sj7iy6));
assign Sj7iy6 = (~(Jexmz6[24] & K94iw6));
assign Kj7iy6 = (Ak7iy6 & Ik7iy6);
assign Ik7iy6 = (~(Lloyx6 & Fd9ov6));
assign Fd9ov6 = (~(Qk7iy6 & Yk7iy6));
assign Yk7iy6 = (Gl7iy6 & Ol7iy6);
assign Ol7iy6 = (Bqoyx6 | Ddg7x6);
assign Ddg7x6 = (Wl7iy6 & Em7iy6);
assign Em7iy6 = (Mm7iy6 & Um7iy6);
assign Um7iy6 = (Cn7iy6 & Kn7iy6);
assign Kn7iy6 = (~(Rmzyx6 & Sn7iy6));
assign Sn7iy6 = (~(Ao7iy6 & Io7iy6));
assign Io7iy6 = (Qo7iy6 & Yo7iy6);
assign Yo7iy6 = (Gp7iy6 & Op7iy6);
assign Op7iy6 = (~(Hyj7z6[7] & Xwciw6));
assign Gp7iy6 = (~(Hyj7z6[0] & Dfk7z6[24]));
assign Qo7iy6 = (Wp7iy6 & Eq7iy6);
assign Eq7iy6 = (~(Hyj7z6[1] & Lpk7z6[24]));
assign Wp7iy6 = (~(Hyj7z6[2] & Tzk7z6[24]));
assign Ao7iy6 = (Mq7iy6 & Uq7iy6);
assign Uq7iy6 = (Cr7iy6 & Kr7iy6);
assign Kr7iy6 = (~(Hyj7z6[3] & Bal7z6[24]));
assign Cr7iy6 = (~(Hyj7z6[4] & Jkl7z6[24]));
assign Mq7iy6 = (Sr7iy6 & As7iy6);
assign As7iy6 = (~(Hyj7z6[5] & Rul7z6[24]));
assign Sr7iy6 = (~(Hyj7z6[6] & Z4m7z6[24]));
assign Cn7iy6 = (~(Xbzyx6 & Is7iy6));
assign Is7iy6 = (~(Qs7iy6 & Ys7iy6));
assign Ys7iy6 = (Gt7iy6 & Ot7iy6);
assign Ot7iy6 = (Wt7iy6 & Eu7iy6);
assign Eu7iy6 = (~(Hyj7z6[0] & Rbk7z6[20]));
assign Wt7iy6 = (~(Hyj7z6[1] & Zlk7z6[20]));
assign Gt7iy6 = (Mu7iy6 & Uu7iy6);
assign Uu7iy6 = (~(Hyj7z6[2] & Hwk7z6[20]));
assign Mu7iy6 = (~(Hyj7z6[3] & P6l7z6[20]));
assign Qs7iy6 = (Cv7iy6 & Kv7iy6);
assign Kv7iy6 = (Sv7iy6 & Aw7iy6);
assign Aw7iy6 = (~(Hyj7z6[4] & Xgl7z6[20]));
assign Sv7iy6 = (~(Hyj7z6[5] & Frl7z6[20]));
assign Cv7iy6 = (Iw7iy6 & Qw7iy6);
assign Qw7iy6 = (~(Hyj7z6[6] & N1m7z6[20]));
assign Iw7iy6 = (~(Hyj7z6[7] & Vbm7z6[20]));
assign Mm7iy6 = (Yw7iy6 & Gx7iy6);
assign Gx7iy6 = (~(Ox7iy6 & Ngqyx6));
assign Ox7iy6 = (~(Wx7iy6 & Ey7iy6));
assign Ey7iy6 = (My7iy6 & Uy7iy6);
assign Uy7iy6 = (Cz7iy6 & Kz7iy6);
assign Kz7iy6 = (Sz7iy6 & Bqyyx6);
assign Bqyyx6 = (~(A8yhy6 & A08iy6));
assign A08iy6 = (~(Hzuyx6 & I08iy6));
assign Sz7iy6 = (~(Q08iy6 & Fs0zx6));
assign Fs0zx6 = (Y08iy6 & G18iy6);
assign G18iy6 = (E32nv6 & D2k7x6);
assign Q08iy6 = (Koaiw6 & Jmqyx6);
assign Cz7iy6 = (O18iy6 & W18iy6);
assign W18iy6 = (~(Ttqyx6 & HTMDHBURST[0]));
assign Ttqyx6 = (~(E28iy6 | I08iy6));
assign O18iy6 = (~(Dheet6 & Buqyx6));
assign My7iy6 = (M28iy6 & U28iy6);
assign U28iy6 = (C38iy6 & K38iy6);
assign K38iy6 = (~(Bzi7z6[24] & Vsqyx6));
assign C38iy6 = (~(Wui7z6[24] & Lxqyx6));
assign M28iy6 = (S38iy6 & A48iy6);
assign A48iy6 = (~(Dri7z6[24] & Fwqyx6));
assign S38iy6 = (~(Bwi7z6[24] & Hzqyx6));
assign Wx7iy6 = (I48iy6 & Q48iy6);
assign Q48iy6 = (Y48iy6 & G58iy6);
assign G58iy6 = (O58iy6 & W58iy6);
assign W58iy6 = (~(Svkhy6 & Pnb7z6[24]));
assign O58iy6 = (~(Pzqyx6 & G5j7z6[56]));
assign Y48iy6 = (E68iy6 & M68iy6);
assign M68iy6 = (~(Jyqyx6 & G5j7z6[24]));
assign E68iy6 = (~(B2ryx6 & M6j7z6[56]));
assign I48iy6 = (U68iy6 & C78iy6);
assign C78iy6 = (K78iy6 & S78iy6);
assign S78iy6 = (~(J2ryx6 & M6j7z6[24]));
assign K78iy6 = (~(D1ryx6 & Ohj7z6[56]));
assign U68iy6 = (Pr0zx6 & A88iy6);
assign A88iy6 = (~(X3ryx6 & Ohj7z6[24]));
assign Pr0zx6 = (Z2ryx6 & Dhsyx6);
assign Dhsyx6 = (~(I88iy6 & Koaiw6));
assign I88iy6 = (Voqyx6 & Q88iy6);
assign Z2ryx6 = (U2vhy6 & Ykthy6);
assign Yw7iy6 = (~(Klo7z6[1] & Y88iy6));
assign Y88iy6 = (~(G98iy6 & O98iy6));
assign O98iy6 = (W98iy6 & Ea8iy6);
assign Ea8iy6 = (Ma8iy6 & Ua8iy6);
assign Ua8iy6 = (~(Bqp7z6[24] & D5qyx6));
assign Ma8iy6 = (Cb8iy6 & Ravyx6);
assign Cb8iy6 = (~(T9tyx6 & Yo77z6));
assign W98iy6 = (Kb8iy6 & Sb8iy6);
assign Sb8iy6 = (~(E6p7z6[24] & L9qyx6));
assign Kb8iy6 = (Ac8iy6 & Ic8iy6);
assign Ic8iy6 = (~(Fk2ft6 & P3a8x6));
assign Ac8iy6 = (~(Gg2ft6 & Ua9ov6));
assign G98iy6 = (Qc8iy6 & Yc8iy6);
assign Yc8iy6 = (Gd8iy6 & Od8iy6);
assign Od8iy6 = (~(Eo2ft6 & Q0a8x6));
assign Gd8iy6 = (Wd8iy6 & Ee8iy6);
assign Ee8iy6 = (~(B2q7z6[24] & Fcqyx6));
assign Wd8iy6 = (~(W94ft6 & Nao7x6));
assign Qc8iy6 = (Me8iy6 & Ue8iy6);
assign Ue8iy6 = (~(Mkp7z6[24] & Tdqyx6));
assign Me8iy6 = (~(Hfqyx6 & U9p7z6[24]));
assign Wl7iy6 = (Cf8iy6 & Kf8iy6);
assign Kf8iy6 = (Sf8iy6 & Ag8iy6);
assign Ag8iy6 = (~(Klo7z6[2] & Ig8iy6));
assign Ig8iy6 = (~(Qg8iy6 & Yg8iy6));
assign Yg8iy6 = (Gh8iy6 & Oh8iy6);
assign Oh8iy6 = (Wh8iy6 & Ei8iy6);
assign Ei8iy6 = (~(Cgset6 & S4kiw6));
assign Wh8iy6 = (Mi8iy6 & Ui8iy6);
assign Ui8iy6 = (~(Nqo7z6[22] & M8kiw6));
assign Mi8iy6 = (~(Fpo7z6[22] & H9kiw6));
assign Gh8iy6 = (Cj8iy6 & Kj8iy6);
assign Kj8iy6 = (~(Ouo7z6[22] & K7kiw6));
assign Cj8iy6 = (~(Hxo7z6[22] & W6kiw6));
assign Qg8iy6 = (Sj8iy6 & Ak8iy6);
assign Ak8iy6 = (Ik8iy6 & Qk8iy6);
assign Qk8iy6 = (~(Vro7z6[22] & Y7kiw6));
assign Ik8iy6 = (~(T2p7z6[24] & U5kiw6));
assign Sj8iy6 = (Yk8iy6 & Gl8iy6);
assign Gl8iy6 = (~(W3p7z6[24] & G5kiw6));
assign Yk8iy6 = (~(A0p7z6[22] & I6kiw6));
assign Sf8iy6 = (~(Bv1nz6[0] & Ol8iy6));
assign Cf8iy6 = (O53iy6 & Wl8iy6);
assign Wl8iy6 = (~(Ies7z6[24] & Tltyx6));
assign Gl7iy6 = (~(Zmoyx6 & Kdg7x6));
assign Kdg7x6 = (~(Em8iy6 & Mm8iy6));
assign Mm8iy6 = (~(Um8iy6 & I8a7z6));
assign I8a7z6 = (~(Cn8iy6 & Kn8iy6));
assign Kn8iy6 = (~(HRDATAD[24] & Qln7z6[0]));
assign Cn8iy6 = (~(HRDATAS[24] & Qln7z6[1]));
assign Em8iy6 = (Sn8iy6 & Ao8iy6);
assign Ao8iy6 = (~(Munhy6 & S7n7z6[1]));
assign Munhy6 = (Lpoyx6 & Evadt6);
assign Lpoyx6 = (Io8iy6 & Qxxet6);
assign Io8iy6 = (Qo8iy6 & A9gxx6);
assign Sn8iy6 = (~(Tim7z6[24] & Yo8iy6));
assign Qk7iy6 = (Gp8iy6 & Op8iy6);
assign Op8iy6 = (~(HRDATAS[24] & Ad47x6));
assign Gp8iy6 = (~(HRDATAD[24] & Mc47x6));
assign Ak7iy6 = (~(Lpryx6 & Yqonv6));
assign Xjo7v6 = (~(Wp8iy6 & Eq8iy6));
assign Eq8iy6 = (~(Jexmz6[25] & K94iw6));
assign Wp8iy6 = (Mq8iy6 & Uq8iy6);
assign Uq8iy6 = (~(Lloyx6 & Vv77x6));
assign Vv77x6 = (~(Cr8iy6 & Kr8iy6));
assign Kr8iy6 = (Sr8iy6 & As8iy6);
assign As8iy6 = (Bqoyx6 | Q9g7x6);
assign Q9g7x6 = (Is8iy6 & Qs8iy6);
assign Qs8iy6 = (Ys8iy6 & Gt8iy6);
assign Gt8iy6 = (Ot8iy6 & Wt8iy6);
assign Wt8iy6 = (~(Rmzyx6 & Eu8iy6));
assign Eu8iy6 = (~(Mu8iy6 & Uu8iy6));
assign Uu8iy6 = (Cv8iy6 & Kv8iy6);
assign Kv8iy6 = (Sv8iy6 & Aw8iy6);
assign Aw8iy6 = (~(Hyj7z6[3] & Sxciw6));
assign Sv8iy6 = (~(Hyj7z6[2] & Lxciw6));
assign Cv8iy6 = (Iw8iy6 & Qw8iy6);
assign Qw8iy6 = (~(Hyj7z6[1] & Exciw6));
assign Iw8iy6 = (~(Hyj7z6[5] & Zxciw6));
assign Mu8iy6 = (Yw8iy6 & Gx8iy6);
assign Gx8iy6 = (Ox8iy6 & Wx8iy6);
assign Wx8iy6 = (~(Hyj7z6[6] & Gyciw6));
assign Ox8iy6 = (~(Hyj7z6[0] & Dfk7z6[25]));
assign Yw8iy6 = (Ey8iy6 & My8iy6);
assign My8iy6 = (~(Hyj7z6[4] & Jkl7z6[25]));
assign Ey8iy6 = (~(Hyj7z6[7] & Hfm7z6[25]));
assign Ot8iy6 = (Uy8iy6 & Cz8iy6);
assign Cz8iy6 = (~(Kz8iy6 & Sz8iy6));
assign Kz8iy6 = (Ok77v6 & D1pyx6);
assign Uy8iy6 = (~(Klo7z6[1] & A09iy6));
assign A09iy6 = (~(I09iy6 & Q09iy6));
assign Q09iy6 = (Y09iy6 & G19iy6);
assign G19iy6 = (~(B2q7z6[25] & Fcqyx6));
assign Y09iy6 = (O19iy6 & W19iy6);
assign W19iy6 = (~(Bqp7z6[25] & D5qyx6));
assign O19iy6 = (~(E6p7z6[25] & L9qyx6));
assign I09iy6 = (E29iy6 & M29iy6);
assign M29iy6 = (~(Mkp7z6[25] & Tdqyx6));
assign E29iy6 = (~(Hfqyx6 & U9p7z6[25]));
assign Ys8iy6 = (U29iy6 & C39iy6);
assign C39iy6 = (~(Xbzyx6 & K39iy6));
assign K39iy6 = (~(S39iy6 & A49iy6));
assign A49iy6 = (I49iy6 & Q49iy6);
assign Q49iy6 = (Y49iy6 & G59iy6);
assign G59iy6 = (~(Hyj7z6[0] & Rbk7z6[21]));
assign Y49iy6 = (~(Hyj7z6[1] & Zlk7z6[21]));
assign I49iy6 = (O59iy6 & W59iy6);
assign W59iy6 = (~(Hyj7z6[2] & Hwk7z6[21]));
assign O59iy6 = (~(Hyj7z6[3] & P6l7z6[21]));
assign S39iy6 = (E69iy6 & M69iy6);
assign M69iy6 = (U69iy6 & C79iy6);
assign C79iy6 = (~(Hyj7z6[4] & Xgl7z6[21]));
assign U69iy6 = (~(Hyj7z6[5] & Frl7z6[21]));
assign E69iy6 = (K79iy6 & S79iy6);
assign S79iy6 = (~(Hyj7z6[6] & N1m7z6[21]));
assign K79iy6 = (~(Hyj7z6[7] & Vbm7z6[21]));
assign U29iy6 = (~(A89iy6 & Ngqyx6));
assign A89iy6 = (~(I89iy6 & Q89iy6));
assign Q89iy6 = (Y89iy6 & G99iy6);
assign G99iy6 = (O99iy6 & W99iy6);
assign W99iy6 = (Ea9iy6 & Ma9iy6);
assign Ma9iy6 = (~(Ijeet6 & Buqyx6));
assign Buqyx6 = (Ua9iy6 & Voqyx6);
assign Ua9iy6 = (!E28iy6);
assign Ea9iy6 = (~(Bzi7z6[25] & Vsqyx6));
assign Vsqyx6 = (~(Ua0iy6 | Zyuyx6));
assign O99iy6 = (Cb9iy6 & Kb9iy6);
assign Kb9iy6 = (~(Wui7z6[25] & Lxqyx6));
assign Cb9iy6 = (~(Dri7z6[25] & Fwqyx6));
assign Y89iy6 = (Sb9iy6 & Ac9iy6);
assign Ac9iy6 = (~(Pzqyx6 & G5j7z6[57]));
assign Sb9iy6 = (Ic9iy6 & Qc9iy6);
assign Qc9iy6 = (~(Bwi7z6[25] & Hzqyx6));
assign Ic9iy6 = (~(Svkhy6 & Pnb7z6[25]));
assign I89iy6 = (Yc9iy6 & Gd9iy6);
assign Gd9iy6 = (Od9iy6 & Wd9iy6);
assign Wd9iy6 = (~(J2ryx6 & M6j7z6[25]));
assign Od9iy6 = (Ee9iy6 & Me9iy6);
assign Me9iy6 = (~(Jyqyx6 & G5j7z6[25]));
assign Ee9iy6 = (~(B2ryx6 & M6j7z6[57]));
assign Yc9iy6 = (Ue9iy6 & Meyhy6);
assign Meyhy6 = (Ywwhy6 & K33iy6);
assign K33iy6 = (~(Lpyyx6 & A8yhy6));
assign Ue9iy6 = (Cf9iy6 & Kf9iy6);
assign Kf9iy6 = (~(D1ryx6 & Ohj7z6[57]));
assign Cf9iy6 = (~(X3ryx6 & Ohj7z6[25]));
assign Is8iy6 = (Sf9iy6 & Ag9iy6);
assign Ag9iy6 = (Ig9iy6 & Qg9iy6);
assign Qg9iy6 = (~(Cr6iy6 & Qo77z6));
assign Ig9iy6 = (Yg9iy6 & Gh9iy6);
assign Gh9iy6 = (~(Klo7z6[2] & Oh9iy6));
assign Oh9iy6 = (~(Wh9iy6 & Ei9iy6));
assign Ei9iy6 = (Mi9iy6 & Ui9iy6);
assign Ui9iy6 = (Cj9iy6 & Kj9iy6);
assign Kj9iy6 = (~(Beset6 & S4kiw6));
assign Cj9iy6 = (Sj9iy6 & Ak9iy6);
assign Ak9iy6 = (~(Nqo7z6[23] & M8kiw6));
assign Sj9iy6 = (~(Fpo7z6[23] & H9kiw6));
assign Mi9iy6 = (Ik9iy6 & Qk9iy6);
assign Qk9iy6 = (~(Ouo7z6[23] & K7kiw6));
assign Ik9iy6 = (~(Hxo7z6[23] & W6kiw6));
assign Wh9iy6 = (Yk9iy6 & Gl9iy6);
assign Gl9iy6 = (Ol9iy6 & Wl9iy6);
assign Wl9iy6 = (~(Vro7z6[23] & Y7kiw6));
assign Ol9iy6 = (~(T2p7z6[25] & U5kiw6));
assign Yk9iy6 = (Em9iy6 & Mm9iy6);
assign Mm9iy6 = (~(W3p7z6[25] & G5kiw6));
assign Em9iy6 = (~(A0p7z6[23] & I6kiw6));
assign Yg9iy6 = (~(Bv1nz6[1] & Ol8iy6));
assign Sf9iy6 = (Um9iy6 & Cn9iy6);
assign Cn9iy6 = (~(Ies7z6[25] & Tltyx6));
assign Sr8iy6 = (~(Zmoyx6 & X9g7x6));
assign X9g7x6 = (~(Kn9iy6 & Sn9iy6));
assign Sn9iy6 = (~(Um8iy6 & A8a7z6));
assign A8a7z6 = (~(Ao9iy6 & Io9iy6));
assign Io9iy6 = (~(HRDATAD[25] & Qln7z6[0]));
assign Ao9iy6 = (~(HRDATAS[25] & Qln7z6[1]));
assign Kn9iy6 = (~(Tim7z6[25] & Yo8iy6));
assign Cr8iy6 = (Qo9iy6 & Yo9iy6);
assign Yo9iy6 = (~(HRDATAS[25] & Ad47x6));
assign Qo9iy6 = (~(HRDATAD[25] & Mc47x6));
assign Mq8iy6 = (~(Lpryx6 & C6q7x6));
assign Qjo7v6 = (~(Gp9iy6 & Op9iy6));
assign Op9iy6 = (~(Jexmz6[26] & K94iw6));
assign Gp9iy6 = (Wp9iy6 & Eq9iy6);
assign Eq9iy6 = (~(Lloyx6 & Bcfov6));
assign Bcfov6 = (~(Mq9iy6 & Uq9iy6));
assign Uq9iy6 = (Cr9iy6 & Kr9iy6);
assign Kr9iy6 = (Bqoyx6 | Ww98x6);
assign Ww98x6 = (Sr9iy6 & As9iy6);
assign As9iy6 = (Is9iy6 & Qs9iy6);
assign Qs9iy6 = (Ys9iy6 & Gt9iy6);
assign Gt9iy6 = (~(Xbzyx6 & Ot9iy6));
assign Ot9iy6 = (~(Wt9iy6 & Eu9iy6));
assign Eu9iy6 = (Mu9iy6 & Uu9iy6);
assign Uu9iy6 = (Cv9iy6 & Kv9iy6);
assign Kv9iy6 = (~(Hyj7z6[0] & Rbk7z6[22]));
assign Cv9iy6 = (~(Hyj7z6[1] & Zlk7z6[22]));
assign Mu9iy6 = (Sv9iy6 & Aw9iy6);
assign Aw9iy6 = (~(Hyj7z6[2] & Hwk7z6[22]));
assign Sv9iy6 = (~(Hyj7z6[3] & P6l7z6[22]));
assign Wt9iy6 = (Iw9iy6 & Qw9iy6);
assign Qw9iy6 = (Yw9iy6 & Gx9iy6);
assign Gx9iy6 = (~(Hyj7z6[4] & Xgl7z6[22]));
assign Yw9iy6 = (~(Hyj7z6[5] & Frl7z6[22]));
assign Iw9iy6 = (Ox9iy6 & Wx9iy6);
assign Wx9iy6 = (~(Hyj7z6[6] & N1m7z6[22]));
assign Ox9iy6 = (~(Hyj7z6[7] & Vbm7z6[22]));
assign Ys9iy6 = (Ey9iy6 & My9iy6);
assign My9iy6 = (~(Klo7z6[1] & Uy9iy6));
assign Uy9iy6 = (~(Cz9iy6 & Kz9iy6));
assign Kz9iy6 = (Sz9iy6 & A0aiy6);
assign A0aiy6 = (~(B2q7z6[26] & Fcqyx6));
assign Sz9iy6 = (I0aiy6 & Q0aiy6);
assign Q0aiy6 = (~(Bqp7z6[26] & D5qyx6));
assign I0aiy6 = (~(E6p7z6[26] & L9qyx6));
assign Cz9iy6 = (Y0aiy6 & G1aiy6);
assign G1aiy6 = (~(Mkp7z6[26] & Tdqyx6));
assign Y0aiy6 = (~(Hfqyx6 & U9p7z6[26]));
assign Ey9iy6 = (~(Rmzyx6 & O1aiy6));
assign O1aiy6 = (~(W1aiy6 & E2aiy6));
assign E2aiy6 = (M2aiy6 & U2aiy6);
assign U2aiy6 = (C3aiy6 & K3aiy6);
assign K3aiy6 = (~(Hyj7z6[3] & Bzciw6));
assign C3aiy6 = (~(Hyj7z6[2] & Uyciw6));
assign M2aiy6 = (S3aiy6 & A4aiy6);
assign A4aiy6 = (~(Hyj7z6[1] & Nyciw6));
assign S3aiy6 = (~(Hyj7z6[5] & Izciw6));
assign W1aiy6 = (I4aiy6 & Q4aiy6);
assign Q4aiy6 = (Y4aiy6 & G5aiy6);
assign G5aiy6 = (~(Hyj7z6[6] & Pzciw6));
assign Y4aiy6 = (~(Hyj7z6[7] & Wzciw6));
assign I4aiy6 = (O5aiy6 & W5aiy6);
assign W5aiy6 = (~(Hyj7z6[0] & Dfk7z6[26]));
assign O5aiy6 = (~(Hyj7z6[4] & Jkl7z6[26]));
assign Is9iy6 = (E6aiy6 & M6aiy6);
assign M6aiy6 = (~(U6aiy6 & Ngqyx6));
assign U6aiy6 = (~(C7aiy6 & K7aiy6));
assign K7aiy6 = (S7aiy6 & A8aiy6);
assign A8aiy6 = (I8aiy6 & Q8aiy6);
assign Q8aiy6 = (~(Dri7z6[26] & Fwqyx6));
assign I8aiy6 = (Y8aiy6 & G9aiy6);
assign G9aiy6 = (~(Dxqyx6 & Zfcet6));
assign Y8aiy6 = (~(Wui7z6[26] & Lxqyx6));
assign S7aiy6 = (O9aiy6 & W9aiy6);
assign W9aiy6 = (~(Pzqyx6 & G5j7z6[58]));
assign O9aiy6 = (Eaaiy6 & Maaiy6);
assign Maaiy6 = (~(Bwi7z6[26] & Hzqyx6));
assign Eaaiy6 = (~(Svkhy6 & Pnb7z6[26]));
assign C7aiy6 = (Uaaiy6 & Cbaiy6);
assign Cbaiy6 = (Kbaiy6 & Sbaiy6);
assign Sbaiy6 = (~(J2ryx6 & M6j7z6[26]));
assign Kbaiy6 = (Acaiy6 & Icaiy6);
assign Icaiy6 = (~(Jyqyx6 & G5j7z6[26]));
assign Acaiy6 = (~(B2ryx6 & M6j7z6[58]));
assign Uaaiy6 = (Qcaiy6 & Ycaiy6);
assign Ycaiy6 = (~(D1ryx6 & Ohj7z6[58]));
assign Qcaiy6 = (~(X3ryx6 & Ohj7z6[26]));
assign E6aiy6 = (~(Klo7z6[2] & Gdaiy6));
assign Gdaiy6 = (~(Odaiy6 & Wdaiy6));
assign Wdaiy6 = (Eeaiy6 & Meaiy6);
assign Meaiy6 = (Ueaiy6 & Cfaiy6);
assign Cfaiy6 = (~(Acset6 & S4kiw6));
assign Ueaiy6 = (Kfaiy6 & Sfaiy6);
assign Sfaiy6 = (~(Nqo7z6[24] & M8kiw6));
assign Kfaiy6 = (~(Fpo7z6[24] & H9kiw6));
assign Eeaiy6 = (Agaiy6 & Igaiy6);
assign Igaiy6 = (~(Ouo7z6[24] & K7kiw6));
assign Agaiy6 = (~(Hxo7z6[24] & W6kiw6));
assign Odaiy6 = (Qgaiy6 & Ygaiy6);
assign Ygaiy6 = (Ghaiy6 & Ohaiy6);
assign Ohaiy6 = (~(Vro7z6[24] & Y7kiw6));
assign Ghaiy6 = (~(T2p7z6[26] & U5kiw6));
assign Qgaiy6 = (Whaiy6 & Eiaiy6);
assign Eiaiy6 = (~(W3p7z6[26] & G5kiw6));
assign Whaiy6 = (~(A0p7z6[24] & I6kiw6));
assign Sr9iy6 = (Miaiy6 & Uiaiy6);
assign Uiaiy6 = (Cjaiy6 & Kjaiy6);
assign Kjaiy6 = (~(W197z6 & Ol8iy6));
assign Cjaiy6 = (~(Cr6iy6 & Io77z6));
assign Miaiy6 = (Yg7iy6 & Sjaiy6);
assign Sjaiy6 = (~(Ies7z6[26] & Tltyx6));
assign Cr9iy6 = (~(HRDATAS[26] & Ad47x6));
assign Mq9iy6 = (Akaiy6 & Ikaiy6);
assign Ikaiy6 = (~(HRDATAD[26] & Mc47x6));
assign Akaiy6 = (~(Zmoyx6 & Dx98x6));
assign Dx98x6 = (~(Qkaiy6 & Ykaiy6));
assign Ykaiy6 = (~(Um8iy6 & S7a7z6));
assign S7a7z6 = (~(Glaiy6 & Olaiy6));
assign Olaiy6 = (~(HRDATAD[26] & Qln7z6[0]));
assign Glaiy6 = (~(HRDATAS[26] & Qln7z6[1]));
assign Qkaiy6 = (~(Tim7z6[26] & Yo8iy6));
assign Wp9iy6 = (~(Lpryx6 & Mbq7x6));
assign Jjo7v6 = (~(Wlaiy6 & Emaiy6));
assign Emaiy6 = (~(Jexmz6[27] & K94iw6));
assign Wlaiy6 = (Mmaiy6 & Umaiy6);
assign Umaiy6 = (~(Lloyx6 & Fmlov6));
assign Fmlov6 = (~(Cnaiy6 & Knaiy6));
assign Knaiy6 = (Snaiy6 & Aoaiy6);
assign Aoaiy6 = (Bqoyx6 | Voyxx6);
assign Voyxx6 = (Ioaiy6 & Qoaiy6);
assign Qoaiy6 = (Yoaiy6 & Gpaiy6);
assign Gpaiy6 = (Opaiy6 & Wpaiy6);
assign Wpaiy6 = (~(Klo7z6[1] & Eqaiy6));
assign Eqaiy6 = (~(Mqaiy6 & Uqaiy6));
assign Uqaiy6 = (Craiy6 & Kraiy6);
assign Kraiy6 = (~(B2q7z6[27] & Fcqyx6));
assign Craiy6 = (Sraiy6 & Asaiy6);
assign Asaiy6 = (~(Bqp7z6[27] & D5qyx6));
assign Sraiy6 = (~(E6p7z6[27] & L9qyx6));
assign Mqaiy6 = (Isaiy6 & Qsaiy6);
assign Qsaiy6 = (~(Mkp7z6[27] & Tdqyx6));
assign Isaiy6 = (~(Hfqyx6 & U9p7z6[27]));
assign Opaiy6 = (Ysaiy6 & Gd2iy6);
assign Ysaiy6 = (~(Gtaiy6 & U2jhy6));
assign Gtaiy6 = (Otaiy6 & K3jhy6);
assign Otaiy6 = (~(Wtaiy6 & Euaiy6));
assign Euaiy6 = (Muaiy6 & Uuaiy6);
assign Uuaiy6 = (Cvaiy6 & Kvaiy6);
assign Kvaiy6 = (~(Hyj7z6[3] & R0diw6));
assign Cvaiy6 = (~(Hyj7z6[2] & K0diw6));
assign Muaiy6 = (Svaiy6 & Awaiy6);
assign Awaiy6 = (~(Hyj7z6[1] & D0diw6));
assign Svaiy6 = (~(Hyj7z6[5] & Y0diw6));
assign Wtaiy6 = (Iwaiy6 & Qwaiy6);
assign Qwaiy6 = (Ywaiy6 & Gxaiy6);
assign Gxaiy6 = (~(Hyj7z6[6] & F1diw6));
assign Ywaiy6 = (~(Hyj7z6[7] & M1diw6));
assign Iwaiy6 = (Oxaiy6 & Wxaiy6);
assign Wxaiy6 = (~(Hyj7z6[0] & Dfk7z6[27]));
assign Oxaiy6 = (~(Hyj7z6[4] & Jkl7z6[27]));
assign Yoaiy6 = (Eyaiy6 & Myaiy6);
assign Myaiy6 = (~(Uyaiy6 & Ngqyx6));
assign Uyaiy6 = (~(Czaiy6 & Kzaiy6));
assign Kzaiy6 = (Szaiy6 & A0biy6);
assign A0biy6 = (I0biy6 & Q0biy6);
assign Q0biy6 = (~(Dri7z6[27] & Fwqyx6));
assign I0biy6 = (Y0biy6 & Ywwhy6);
assign Y0biy6 = (~(Wui7z6[27] & Lxqyx6));
assign Szaiy6 = (G1biy6 & O1biy6);
assign O1biy6 = (~(Pzqyx6 & G5j7z6[59]));
assign G1biy6 = (W1biy6 & E2biy6);
assign E2biy6 = (~(Bwi7z6[27] & Hzqyx6));
assign W1biy6 = (~(Svkhy6 & Pnb7z6[27]));
assign Czaiy6 = (M2biy6 & U2biy6);
assign U2biy6 = (C3biy6 & K3biy6);
assign K3biy6 = (~(J2ryx6 & M6j7z6[27]));
assign C3biy6 = (S3biy6 & A4biy6);
assign A4biy6 = (~(Jyqyx6 & G5j7z6[27]));
assign S3biy6 = (~(B2ryx6 & M6j7z6[59]));
assign M2biy6 = (I4biy6 & Q4biy6);
assign Q4biy6 = (~(D1ryx6 & Ohj7z6[59]));
assign I4biy6 = (~(X3ryx6 & Ohj7z6[27]));
assign Eyaiy6 = (~(Klo7z6[2] & Y4biy6));
assign Y4biy6 = (~(G5biy6 & O5biy6));
assign O5biy6 = (W5biy6 & E6biy6);
assign E6biy6 = (M6biy6 & U6biy6);
assign U6biy6 = (~(Z9set6 & S4kiw6));
assign M6biy6 = (C7biy6 & K7biy6);
assign K7biy6 = (~(Nqo7z6[25] & M8kiw6));
assign C7biy6 = (~(Fpo7z6[25] & H9kiw6));
assign W5biy6 = (S7biy6 & A8biy6);
assign A8biy6 = (~(Ouo7z6[25] & K7kiw6));
assign S7biy6 = (~(Hxo7z6[25] & W6kiw6));
assign G5biy6 = (I8biy6 & Q8biy6);
assign Q8biy6 = (Y8biy6 & G9biy6);
assign G9biy6 = (~(Vro7z6[25] & Y7kiw6));
assign Y8biy6 = (~(T2p7z6[27] & U5kiw6));
assign I8biy6 = (O9biy6 & W9biy6);
assign W9biy6 = (~(W3p7z6[27] & G5kiw6));
assign O9biy6 = (~(A0p7z6[25] & I6kiw6));
assign Ioaiy6 = (Eabiy6 & Mabiy6);
assign Mabiy6 = (Uabiy6 & Cbbiy6);
assign Cbbiy6 = (~(Pp1nz6[0] & Ol8iy6));
assign Uabiy6 = (~(Cr6iy6 & Ao77z6));
assign Eabiy6 = (Yg7iy6 & Kbbiy6);
assign Kbbiy6 = (~(Ies7z6[27] & Tltyx6));
assign Snaiy6 = (~(Zmoyx6 & Dpyxx6));
assign Dpyxx6 = (~(Sbbiy6 & Acbiy6));
assign Acbiy6 = (~(Um8iy6 & K7a7z6));
assign K7a7z6 = (~(Icbiy6 & Qcbiy6));
assign Qcbiy6 = (~(HRDATAD[27] & Qln7z6[0]));
assign Icbiy6 = (~(HRDATAS[27] & Qln7z6[1]));
assign Sbbiy6 = (~(Tim7z6[27] & Yo8iy6));
assign Cnaiy6 = (Ycbiy6 & Gdbiy6);
assign Gdbiy6 = (~(HRDATAS[27] & Ad47x6));
assign Ycbiy6 = (~(HRDATAD[27] & Mc47x6));
assign Mmaiy6 = (~(Lpryx6 & Wgq7x6));
assign Cjo7v6 = (~(Odbiy6 & Wdbiy6));
assign Wdbiy6 = (~(Jexmz6[28] & K94iw6));
assign Odbiy6 = (Eebiy6 & Mebiy6);
assign Mebiy6 = (~(Lloyx6 & T977x6));
assign T977x6 = (~(Uebiy6 & Cfbiy6));
assign Cfbiy6 = (Kfbiy6 & Sfbiy6);
assign Sfbiy6 = (Bqoyx6 | Vsyxx6);
assign Vsyxx6 = (Agbiy6 & Igbiy6);
assign Igbiy6 = (Qgbiy6 & Ygbiy6);
assign Ygbiy6 = (Ghbiy6 & Ohbiy6);
assign Ohbiy6 = (~(Klo7z6[1] & Whbiy6));
assign Whbiy6 = (~(Eibiy6 & Mibiy6));
assign Mibiy6 = (Uibiy6 & Cjbiy6);
assign Cjbiy6 = (~(B2q7z6[28] & Fcqyx6));
assign Uibiy6 = (Kjbiy6 & Sjbiy6);
assign Sjbiy6 = (~(Bqp7z6[28] & D5qyx6));
assign Kjbiy6 = (~(E6p7z6[28] & L9qyx6));
assign Eibiy6 = (Akbiy6 & Ikbiy6);
assign Ikbiy6 = (~(Mkp7z6[28] & Tdqyx6));
assign Akbiy6 = (~(Hfqyx6 & U9p7z6[28]));
assign Ghbiy6 = (Qkbiy6 & Gd2iy6);
assign Gd2iy6 = (~(Ykbiy6 & D1pyx6));
assign Ykbiy6 = (Ied8x6 & W5qhy6);
assign Qkbiy6 = (~(Yg3iy6 & Xz67v6));
assign Yg3iy6 = (Iknhy6 & Klo7z6[3]);
assign Iknhy6 = (Fgpyx6 & Mphiw6);
assign Qgbiy6 = (Glbiy6 & Olbiy6);
assign Olbiy6 = (~(Xbzyx6 & Wlbiy6));
assign Wlbiy6 = (~(Embiy6 & Mmbiy6));
assign Mmbiy6 = (Umbiy6 & Cnbiy6);
assign Cnbiy6 = (Knbiy6 & Snbiy6);
assign Snbiy6 = (~(Rbk7z6[23] & Hyj7z6[0]));
assign Knbiy6 = (~(Zlk7z6[23] & Hyj7z6[1]));
assign Umbiy6 = (Aobiy6 & Iobiy6);
assign Iobiy6 = (~(Hwk7z6[23] & Hyj7z6[2]));
assign Aobiy6 = (~(P6l7z6[23] & Hyj7z6[3]));
assign Embiy6 = (Qobiy6 & Yobiy6);
assign Yobiy6 = (Gpbiy6 & Opbiy6);
assign Opbiy6 = (~(Xgl7z6[23] & Hyj7z6[4]));
assign Gpbiy6 = (~(Frl7z6[23] & Hyj7z6[5]));
assign Qobiy6 = (Wpbiy6 & Eqbiy6);
assign Eqbiy6 = (~(N1m7z6[23] & Hyj7z6[6]));
assign Wpbiy6 = (~(Vbm7z6[23] & Hyj7z6[7]));
assign Xbzyx6 = (Mqbiy6 & Klo7z6[5]);
assign Mqbiy6 = (K3jhy6 & Rediw6);
assign Glbiy6 = (Uqbiy6 & Crbiy6);
assign Crbiy6 = (~(Krbiy6 & Ngqyx6));
assign Krbiy6 = (~(Srbiy6 & Asbiy6));
assign Asbiy6 = (Isbiy6 & Qsbiy6);
assign Qsbiy6 = (Ysbiy6 & Gtbiy6);
assign Gtbiy6 = (~(Wui7z6[28] & Lxqyx6));
assign Ysbiy6 = (Otbiy6 & Ywwhy6);
assign Otbiy6 = (~(Dxqyx6 & Fhcet6));
assign Isbiy6 = (Wtbiy6 & Eubiy6);
assign Eubiy6 = (~(Svkhy6 & Pnb7z6[28]));
assign Wtbiy6 = (Mubiy6 & Uubiy6);
assign Uubiy6 = (~(Dri7z6[28] & Fwqyx6));
assign Mubiy6 = (~(Bwi7z6[28] & Hzqyx6));
assign Srbiy6 = (Cvbiy6 & Kvbiy6);
assign Kvbiy6 = (Svbiy6 & Awbiy6);
assign Awbiy6 = (~(B2ryx6 & M6j7z6[60]));
assign Svbiy6 = (Iwbiy6 & Qwbiy6);
assign Qwbiy6 = (~(Pzqyx6 & G5j7z6[60]));
assign Iwbiy6 = (~(Jyqyx6 & G5j7z6[28]));
assign Cvbiy6 = (Ywbiy6 & Gxbiy6);
assign Gxbiy6 = (~(X3ryx6 & Ohj7z6[28]));
assign Ywbiy6 = (Oxbiy6 & Wxbiy6);
assign Wxbiy6 = (~(J2ryx6 & M6j7z6[28]));
assign Oxbiy6 = (~(D1ryx6 & Ohj7z6[60]));
assign Uqbiy6 = (~(Rmzyx6 & Eybiy6));
assign Eybiy6 = (~(Mybiy6 & Uybiy6));
assign Uybiy6 = (Czbiy6 & Kzbiy6);
assign Kzbiy6 = (Szbiy6 & A0ciy6);
assign A0ciy6 = (~(Hyj7z6[3] & O2diw6));
assign Szbiy6 = (~(Hyj7z6[2] & H2diw6));
assign Czbiy6 = (I0ciy6 & Q0ciy6);
assign Q0ciy6 = (~(Hyj7z6[1] & A2diw6));
assign I0ciy6 = (~(Hyj7z6[5] & V2diw6));
assign Mybiy6 = (Y0ciy6 & G1ciy6);
assign G1ciy6 = (O1ciy6 & W1ciy6);
assign W1ciy6 = (~(Hyj7z6[6] & J3diw6));
assign O1ciy6 = (~(Hyj7z6[7] & Q3diw6));
assign Y0ciy6 = (E2ciy6 & M2ciy6);
assign M2ciy6 = (~(Hyj7z6[0] & Dfk7z6[28]));
assign E2ciy6 = (~(Hyj7z6[4] & Jkl7z6[28]));
assign Rmzyx6 = (U2jhy6 & K3jhy6);
assign Agbiy6 = (U2ciy6 & C3ciy6);
assign C3ciy6 = (K3ciy6 & S3ciy6);
assign S3ciy6 = (~(Cr6iy6 & Sn77z6));
assign K3ciy6 = (A4ciy6 & I4ciy6);
assign I4ciy6 = (~(Klo7z6[2] & Q4ciy6));
assign Q4ciy6 = (~(Y4ciy6 & G5ciy6));
assign G5ciy6 = (O5ciy6 & W5ciy6);
assign W5ciy6 = (E6ciy6 & M6ciy6);
assign M6ciy6 = (~(Y7set6 & S4kiw6));
assign E6ciy6 = (U6ciy6 & C7ciy6);
assign C7ciy6 = (~(Nqo7z6[26] & M8kiw6));
assign M8kiw6 = (~(K7ciy6 | Z4p7z6[0]));
assign U6ciy6 = (~(Fpo7z6[26] & H9kiw6));
assign H9kiw6 = (S7ciy6 & Z4p7z6[0]);
assign S7ciy6 = (!K7ciy6);
assign K7ciy6 = (~(A8ciy6 & I8ciy6));
assign I8ciy6 = (Q8ciy6 & Uamhy6);
assign Q8ciy6 = (~(Z4p7z6[2] | Z4p7z6[5]));
assign A8ciy6 = (Z4p7z6[4] & Z4p7z6[3]);
assign O5ciy6 = (Y8ciy6 & G9ciy6);
assign G9ciy6 = (~(Ouo7z6[26] & K7kiw6));
assign Y8ciy6 = (~(Hxo7z6[26] & W6kiw6));
assign Y4ciy6 = (O9ciy6 & W9ciy6);
assign W9ciy6 = (Eaciy6 & Maciy6);
assign Maciy6 = (~(Vro7z6[26] & Y7kiw6));
assign Eaciy6 = (~(T2p7z6[28] & U5kiw6));
assign O9ciy6 = (Uaciy6 & Cbciy6);
assign Cbciy6 = (~(W3p7z6[28] & G5kiw6));
assign Uaciy6 = (~(A0p7z6[26] & I6kiw6));
assign A4ciy6 = (~(Pp1nz6[1] & Ol8iy6));
assign U2ciy6 = (Um9iy6 & Kbciy6);
assign Kbciy6 = (~(Ies7z6[28] & Tltyx6));
assign Kfbiy6 = (~(Zmoyx6 & Dtyxx6));
assign Dtyxx6 = (~(Sbciy6 & Acciy6));
assign Acciy6 = (~(Um8iy6 & C7a7z6));
assign C7a7z6 = (~(Icciy6 & Qcciy6));
assign Qcciy6 = (~(HRDATAD[28] & Qln7z6[0]));
assign Icciy6 = (~(HRDATAS[28] & Qln7z6[1]));
assign Sbciy6 = (~(Tim7z6[28] & Yo8iy6));
assign Uebiy6 = (Ycciy6 & Gdciy6);
assign Gdciy6 = (~(HRDATAS[28] & Ad47x6));
assign Ycciy6 = (~(HRDATAD[28] & Mc47x6));
assign Eebiy6 = (~(Lpryx6 & Gmq7x6));
assign Vio7v6 = (~(Odciy6 & Wdciy6));
assign Wdciy6 = (~(Jexmz6[29] & K94iw6));
assign Odciy6 = (Eeciy6 & Meciy6);
assign Meciy6 = (~(Lloyx6 & T277x6));
assign T277x6 = (~(Ueciy6 & Cfciy6));
assign Cfciy6 = (Kfciy6 & Sfciy6);
assign Sfciy6 = (Bqoyx6 | Xvjyx6);
assign Xvjyx6 = (Agciy6 & Igciy6);
assign Igciy6 = (Qgciy6 & Ygciy6);
assign Ygciy6 = (Ghciy6 & Ohciy6);
assign Ohciy6 = (~(Whciy6 & U2jhy6));
assign Whciy6 = (Eiciy6 & K3jhy6);
assign Eiciy6 = (~(Miciy6 & Uiciy6));
assign Uiciy6 = (Cjciy6 & Kjciy6);
assign Kjciy6 = (Sjciy6 & Akciy6);
assign Akciy6 = (~(Hyj7z6[3] & L4diw6));
assign Sjciy6 = (~(Hyj7z6[2] & E4diw6));
assign Cjciy6 = (Ikciy6 & Qkciy6);
assign Qkciy6 = (~(Hyj7z6[1] & X3diw6));
assign Ikciy6 = (~(Hyj7z6[5] & S4diw6));
assign Miciy6 = (Ykciy6 & Glciy6);
assign Glciy6 = (Olciy6 & Wlciy6);
assign Wlciy6 = (~(Hyj7z6[6] & Z4diw6));
assign Olciy6 = (~(Hyj7z6[7] & G5diw6));
assign Ykciy6 = (Emciy6 & Mmciy6);
assign Mmciy6 = (~(Hyj7z6[0] & Dfk7z6[29]));
assign Emciy6 = (~(Hyj7z6[4] & Jkl7z6[29]));
assign Ghciy6 = (~(Klo7z6[1] & Umciy6));
assign Umciy6 = (~(Cnciy6 & Knciy6));
assign Knciy6 = (Snciy6 & Aociy6);
assign Aociy6 = (~(B2q7z6[29] & Fcqyx6));
assign Snciy6 = (Iociy6 & Qociy6);
assign Qociy6 = (~(Bqp7z6[29] & D5qyx6));
assign Iociy6 = (~(E6p7z6[29] & L9qyx6));
assign Cnciy6 = (Yociy6 & Gpciy6);
assign Gpciy6 = (~(Mkp7z6[29] & Tdqyx6));
assign Yociy6 = (~(Hfqyx6 & U9p7z6[29]));
assign Qgciy6 = (Opciy6 & Wpciy6);
assign Wpciy6 = (~(Txhyx6 & Ol8iy6));
assign Ol8iy6 = (Xjtyx6 | Pjtyx6);
assign Pjtyx6 = (U2mhy6 & Klo7z6[3]);
assign U2mhy6 = (~(Gl5ov6 | Qgnhy6));
assign Gl5ov6 = (!Ri3yx6);
assign Ri3yx6 = (~(Eqciy6 | Puhiw6));
assign Xjtyx6 = (S3mhy6 & Klo7z6[3]);
assign S3mhy6 = (~(P72yx6 | Qgnhy6));
assign Txhyx6 = (Ig27v6 ? Ln6ft6 : La6ft6);
assign Opciy6 = (~(Mqciy6 & Ngqyx6));
assign Mqciy6 = (~(Uqciy6 & Crciy6));
assign Crciy6 = (Krciy6 & Srciy6);
assign Srciy6 = (Asciy6 & Isciy6);
assign Isciy6 = (Qsciy6 & Ysciy6);
assign Ysciy6 = (Ykthy6 & Ywwhy6);
assign Ykthy6 = (~(A8yhy6 & Jmqyx6));
assign A8yhy6 = (Q88iy6 & Tpyyx6);
assign Q88iy6 = (Gtciy6 & Otciy6);
assign Otciy6 = (Toi7z6[6] & D2k7x6);
assign D2k7x6 = (!Toi7z6[7]);
assign Gtciy6 = (Wtciy6 & Toi7z6[5]);
assign Qsciy6 = (Euciy6 & Muciy6);
assign Muciy6 = (~(Uuciy6 & Nksyx6));
assign Uuciy6 = (Hjsyx6 & Gaj7z6[0]);
assign Euciy6 = (~(Wui7z6[29] & Lxqyx6));
assign Asciy6 = (Cvciy6 & Kvciy6);
assign Kvciy6 = (Svciy6 & Awciy6);
assign Awciy6 = (~(Dri7z6[29] & Fwqyx6));
assign Svciy6 = (~(Bwi7z6[29] & Hzqyx6));
assign Cvciy6 = (Iwciy6 & Qwciy6);
assign Qwciy6 = (~(Ba0zx6 & T7j7z6[0]));
assign Iwciy6 = (~(Svkhy6 & Pnb7z6[29]));
assign Krciy6 = (Ywciy6 & Gxciy6);
assign Gxciy6 = (Oxciy6 & Wxciy6);
assign Wxciy6 = (Eyciy6 & Myciy6);
assign Myciy6 = (~(D90zx6 & Lgj7z6[189]));
assign Eyciy6 = (~(Za0zx6 & Lgj7z6[177]));
assign Oxciy6 = (Uyciy6 & Czciy6);
assign Czciy6 = (~(Hb0zx6 & Lgj7z6[165]));
assign Uyciy6 = (~(Vc0zx6 & Lgj7z6[153]));
assign Ywciy6 = (Kzciy6 & Szciy6);
assign Szciy6 = (~(Je0zx6 & Lgj7z6[117]));
assign Kzciy6 = (A0diy6 & I0diy6);
assign I0diy6 = (~(Dd0zx6 & Lgj7z6[141]));
assign A0diy6 = (~(Be0zx6 & Lgj7z6[129]));
assign Uqciy6 = (Q0diy6 & Y0diy6);
assign Y0diy6 = (G1diy6 & O1diy6);
assign O1diy6 = (W1diy6 & E2diy6);
assign E2diy6 = (M2diy6 & U2diy6);
assign U2diy6 = (~(Bi0zx6 & Lgj7z6[105]));
assign M2diy6 = (~(Ji0zx6 & Lgj7z6[93]));
assign W1diy6 = (C3diy6 & K3diy6);
assign K3diy6 = (~(Dh0zx6 & Lgj7z6[81]));
assign C3diy6 = (~(Hj0zx6 & Lgj7z6[69]));
assign G1diy6 = (S3diy6 & A4diy6);
assign A4diy6 = (I4diy6 & Q4diy6);
assign Q4diy6 = (~(Pj0zx6 & Lgj7z6[57]));
assign I4diy6 = (~(Dl0zx6 & Lgj7z6[45]));
assign S3diy6 = (Y4diy6 & G5diy6);
assign G5diy6 = (~(Ll0zx6 & Lgj7z6[33]));
assign Y4diy6 = (~(Jm0zx6 & Lgj7z6[21]));
assign Q0diy6 = (O5diy6 & W5diy6);
assign W5diy6 = (E6diy6 & M6diy6);
assign M6diy6 = (U6diy6 & C7diy6);
assign C7diy6 = (~(Rm0zx6 & Lgj7z6[9]));
assign U6diy6 = (~(Pzqyx6 & G5j7z6[61]));
assign E6diy6 = (K7diy6 & S7diy6);
assign S7diy6 = (~(Jyqyx6 & G5j7z6[29]));
assign K7diy6 = (~(B2ryx6 & M6j7z6[61]));
assign O5diy6 = (A8diy6 & I8diy6);
assign I8diy6 = (~(X3ryx6 & Ohj7z6[29]));
assign A8diy6 = (Q8diy6 & Y8diy6);
assign Y8diy6 = (~(J2ryx6 & M6j7z6[29]));
assign Q8diy6 = (~(D1ryx6 & Ohj7z6[61]));
assign Agciy6 = (G9diy6 & O9diy6);
assign O9diy6 = (W9diy6 & Eadiy6);
assign Eadiy6 = (~(S4kiw6 & Klo7z6[2]));
assign S4kiw6 = (Madiy6 & A0phy6);
assign Madiy6 = (Z4p7z6[0] & Uamhy6);
assign Uamhy6 = (!Z4p7z6[1]);
assign W9diy6 = (~(Cr6iy6 & Kn77z6));
assign G9diy6 = (Um9iy6 & Uadiy6);
assign Uadiy6 = (~(Ies7z6[29] & Tltyx6));
assign Kfciy6 = (~(Zmoyx6 & Fwjyx6));
assign Fwjyx6 = (~(Cbdiy6 & Kbdiy6));
assign Kbdiy6 = (~(Um8iy6 & U6a7z6));
assign U6a7z6 = (~(Sbdiy6 & Acdiy6));
assign Acdiy6 = (~(HRDATAD[29] & Qln7z6[0]));
assign Sbdiy6 = (~(HRDATAS[29] & Qln7z6[1]));
assign Cbdiy6 = (~(Tim7z6[29] & Yo8iy6));
assign Ueciy6 = (Icdiy6 & Qcdiy6);
assign Qcdiy6 = (~(HRDATAS[29] & Ad47x6));
assign Icdiy6 = (~(HRDATAD[29] & Mc47x6));
assign Eeciy6 = (~(Lpryx6 & Qrq7x6));
assign Oio7v6 = (~(Ycdiy6 & Gddiy6));
assign Gddiy6 = (~(Jexmz6[30] & K94iw6));
assign Ycdiy6 = (Oddiy6 & Wddiy6);
assign Wddiy6 = (~(Lloyx6 & Tv67x6));
assign Tv67x6 = (~(Eediy6 & Mediy6));
assign Mediy6 = (Uediy6 & Cfdiy6);
assign Cfdiy6 = (~(Kfdiy6 & Sfdiy6));
assign Uediy6 = (~(Zmoyx6 & Agdiy6));
assign Eediy6 = (Igdiy6 & Qgdiy6);
assign Qgdiy6 = (~(HRDATAS[30] & Ad47x6));
assign Igdiy6 = (~(HRDATAD[30] & Mc47x6));
assign Oddiy6 = (~(Lpryx6 & Vxq7x6));
assign Hio7v6 = (~(Ygdiy6 & Ghdiy6));
assign Ghdiy6 = (~(Jexmz6[31] & K94iw6));
assign Ygdiy6 = (Ohdiy6 & Whdiy6);
assign Whdiy6 = (~(Lpryx6 & Ht1ov6));
assign Lpryx6 = (~(K94iw6 | Cjh7v6));
assign Ohdiy6 = (~(Lloyx6 & Kn67x6));
assign Kn67x6 = (~(Eidiy6 & Midiy6));
assign Midiy6 = (Uidiy6 & Cjdiy6);
assign Cjdiy6 = (Bqoyx6 | Dbwnv6);
assign Dbwnv6 = (Kjdiy6 & Sjdiy6);
assign Sjdiy6 = (Akdiy6 & Ikdiy6);
assign Ikdiy6 = (Qkdiy6 & Ykdiy6);
assign Ykdiy6 = (~(Gldiy6 & U2jhy6));
assign Gldiy6 = (Oldiy6 & K3jhy6);
assign Oldiy6 = (~(Wldiy6 & Emdiy6));
assign Emdiy6 = (Mmdiy6 & Umdiy6);
assign Umdiy6 = (Cndiy6 & Kndiy6);
assign Kndiy6 = (~(Hyj7z6[3] & Jadiw6));
assign Cndiy6 = (Ldsyx6 | Sr87z6);
assign Ldsyx6 = (!Hyj7z6[2]);
assign Mmdiy6 = (Sndiy6 & Aodiy6);
assign Aodiy6 = (Tlpyx6 | Yk87z6);
assign Tlpyx6 = (!Hyj7z6[1]);
assign Sndiy6 = (Llpyx6 | Ee87z6);
assign Llpyx6 = (!Hyj7z6[5]);
assign Wldiy6 = (Iodiy6 & Qodiy6);
assign Qodiy6 = (Yodiy6 & Gpdiy6);
assign Gpdiy6 = (Ddsyx6 | K787z6);
assign Ddsyx6 = (!Hyj7z6[6]);
assign Yodiy6 = (C09iw6 | Iw77z6);
assign C09iw6 = (!Hyj7z6[7]);
assign Iodiy6 = (Opdiy6 & Wpdiy6);
assign Wpdiy6 = (~(Hyj7z6[0] & Dfk7z6[31]));
assign Opdiy6 = (~(Hyj7z6[4] & Jkl7z6[31]));
assign Qkdiy6 = (~(Klo7z6[1] & Eqdiy6));
assign Eqdiy6 = (~(Mqdiy6 & Uqdiy6));
assign Uqdiy6 = (Crdiy6 & Krdiy6);
assign Krdiy6 = (~(B2q7z6[31] & Fcqyx6));
assign Crdiy6 = (Srdiy6 & Asdiy6);
assign Asdiy6 = (~(Bqp7z6[31] & D5qyx6));
assign Srdiy6 = (~(E6p7z6[31] & L9qyx6));
assign Mqdiy6 = (Isdiy6 & Qsdiy6);
assign Qsdiy6 = (~(Mkp7z6[31] & Tdqyx6));
assign Isdiy6 = (~(Hfqyx6 & U9p7z6[31]));
assign Akdiy6 = (Ysdiy6 & Gtdiy6);
assign Gtdiy6 = (~(Klo7z6[2] & Otdiy6));
assign Otdiy6 = (~(Wtdiy6 & Eudiy6));
assign Eudiy6 = (Mudiy6 & Uudiy6);
assign Uudiy6 = (~(Dto7z6[1] & Y7kiw6));
assign Mudiy6 = (Cvdiy6 & Kvdiy6);
assign Kvdiy6 = (~(Wvo7z6[1] & K7kiw6));
assign Cvdiy6 = (~(Pyo7z6[1] & W6kiw6));
assign Wtdiy6 = (Svdiy6 & Awdiy6);
assign Awdiy6 = (~(I1p7z6[1] & I6kiw6));
assign Svdiy6 = (Iwdiy6 & Qwdiy6);
assign Qwdiy6 = (~(Cu1ft6 & U5kiw6));
assign Iwdiy6 = (~(Tx1ft6 & G5kiw6));
assign Ysdiy6 = (~(Cr6iy6 & Um77z6));
assign Kjdiy6 = (Ywdiy6 & Yg7iy6);
assign Yg7iy6 = (Um9iy6 & Gxdiy6);
assign Gxdiy6 = (~(Ys0iy6 & D1pyx6));
assign Ys0iy6 = (P3xyx6 & J2xyx6);
assign Um9iy6 = (Oxdiy6 & Qg3iy6);
assign Oxdiy6 = (~(Cr6iy6 & A9i8v6));
assign Cr6iy6 = (Klo7z6[1] & T9tyx6);
assign Ywdiy6 = (Wxdiy6 & Eydiy6);
assign Eydiy6 = (~(Mydiy6 & Ngqyx6));
assign Mydiy6 = (~(Uydiy6 & Czdiy6));
assign Czdiy6 = (Kzdiy6 & Szdiy6);
assign Szdiy6 = (A0eiy6 & I0eiy6);
assign I0eiy6 = (Q0eiy6 & Y0eiy6);
assign Y0eiy6 = (G1eiy6 & Ywwhy6);
assign G1eiy6 = (~(Hjsyx6 & O1eiy6));
assign O1eiy6 = (~(W1eiy6 & E2eiy6));
assign E2eiy6 = (~(Nksyx6 & Gaj7z6[2]));
assign W1eiy6 = (~(Byi7z6[31] & Zisyx6));
assign Q0eiy6 = (M2eiy6 & U2eiy6);
assign U2eiy6 = (~(Hdcet6 & Dxqyx6));
assign Dxqyx6 = (C3eiy6 & Lpyyx6);
assign M2eiy6 = (~(Wui7z6[31] & Lxqyx6));
assign A0eiy6 = (K3eiy6 & S3eiy6);
assign S3eiy6 = (A4eiy6 & I4eiy6);
assign I4eiy6 = (~(Dri7z6[31] & Fwqyx6));
assign A4eiy6 = (~(Bwi7z6[31] & Hzqyx6));
assign K3eiy6 = (Q4eiy6 & Y4eiy6);
assign Y4eiy6 = (~(Ba0zx6 & T7j7z6[2]));
assign Q4eiy6 = (~(Svkhy6 & Pnb7z6[31]));
assign Kzdiy6 = (G5eiy6 & O5eiy6);
assign O5eiy6 = (W5eiy6 & E6eiy6);
assign E6eiy6 = (M6eiy6 & U6eiy6);
assign U6eiy6 = (~(D90zx6 & Lgj7z6[191]));
assign M6eiy6 = (~(Za0zx6 & Lgj7z6[179]));
assign W5eiy6 = (C7eiy6 & K7eiy6);
assign K7eiy6 = (~(Hb0zx6 & Lgj7z6[167]));
assign C7eiy6 = (~(Vc0zx6 & Lgj7z6[155]));
assign G5eiy6 = (S7eiy6 & A8eiy6);
assign A8eiy6 = (I8eiy6 & Q8eiy6);
assign Q8eiy6 = (~(Dd0zx6 & Lgj7z6[143]));
assign I8eiy6 = (~(Be0zx6 & Lgj7z6[131]));
assign S7eiy6 = (Y8eiy6 & G9eiy6);
assign G9eiy6 = (~(Je0zx6 & Lgj7z6[119]));
assign Y8eiy6 = (~(Bi0zx6 & Lgj7z6[107]));
assign Uydiy6 = (O9eiy6 & W9eiy6);
assign W9eiy6 = (Eaeiy6 & Maeiy6);
assign Maeiy6 = (Uaeiy6 & Cbeiy6);
assign Cbeiy6 = (Kbeiy6 & Sbeiy6);
assign Sbeiy6 = (~(Ji0zx6 & Lgj7z6[95]));
assign Kbeiy6 = (~(Dh0zx6 & Lgj7z6[83]));
assign Uaeiy6 = (Aceiy6 & Iceiy6);
assign Iceiy6 = (~(Hj0zx6 & Lgj7z6[71]));
assign Aceiy6 = (~(Pj0zx6 & Lgj7z6[59]));
assign Eaeiy6 = (Qceiy6 & Yceiy6);
assign Yceiy6 = (Gdeiy6 & Odeiy6);
assign Odeiy6 = (~(Dl0zx6 & Lgj7z6[47]));
assign Gdeiy6 = (~(Ll0zx6 & Lgj7z6[35]));
assign Qceiy6 = (Wdeiy6 & Eeeiy6);
assign Eeeiy6 = (~(Jm0zx6 & Lgj7z6[23]));
assign Wdeiy6 = (~(Rm0zx6 & Lgj7z6[11]));
assign O9eiy6 = (Meeiy6 & Ueeiy6);
assign Ueeiy6 = (Cfeiy6 & Kfeiy6);
assign Kfeiy6 = (Sfeiy6 & Ageiy6);
assign Ageiy6 = (~(Pzqyx6 & G5j7z6[63]));
assign Sfeiy6 = (~(Jyqyx6 & G5j7z6[31]));
assign Cfeiy6 = (Igeiy6 & Qgeiy6);
assign Qgeiy6 = (~(B2ryx6 & M6j7z6[63]));
assign Igeiy6 = (~(J2ryx6 & M6j7z6[31]));
assign Meeiy6 = (Ygeiy6 & Gheiy6);
assign Gheiy6 = (~(STCALIB[25] & F4ryx6));
assign Ygeiy6 = (Oheiy6 & Wheiy6);
assign Wheiy6 = (~(D1ryx6 & Ohj7z6[63]));
assign Oheiy6 = (~(X3ryx6 & Ohj7z6[31]));
assign Wxdiy6 = (~(Ies7z6[31] & Tltyx6));
assign Bqoyx6 = (!Kfdiy6);
assign Uidiy6 = (~(Zmoyx6 & Kbwnv6));
assign Eidiy6 = (Eieiy6 & Mieiy6);
assign Mieiy6 = (~(HRDATAS[31] & Ad47x6));
assign Eieiy6 = (~(HRDATAD[31] & Mc47x6));
assign Lloyx6 = (Cjh7v6 & Ob4iw6);
assign Aio7v6 = (~(Uieiy6 & Cjeiy6));
assign Cjeiy6 = (~(Fcwnv6 & Zqyhw6));
assign Zqyhw6 = (JTAGNSW ? Aixmz6[30] : Ulxmz6[30]);
assign Fcwnv6 = (Dbymz6[0] & Fvd7x6);
assign Uieiy6 = (Kjeiy6 & Sjeiy6);
assign Sjeiy6 = (~(G9wnv6 & Akeiy6));
assign Akeiy6 = (~(Ikeiy6 & Qkeiy6));
assign Qkeiy6 = (Ykeiy6 & Gleiy6);
assign Gleiy6 = (~(Dtm7z6[2] & Sfdiy6));
assign Sfdiy6 = (~(Oleiy6 & Wleiy6));
assign Wleiy6 = (Emeiy6 & Mmeiy6);
assign Mmeiy6 = (~(Klo7z6[1] & Umeiy6));
assign Umeiy6 = (~(Cneiy6 & Kneiy6));
assign Kneiy6 = (Sneiy6 & Aoeiy6);
assign Aoeiy6 = (Ravyx6 & Ioeiy6);
assign Ioeiy6 = (!B6qyx6);
assign Ravyx6 = (~(A9i8v6 & T9tyx6));
assign Sneiy6 = (Qoeiy6 & Yoeiy6);
assign Yoeiy6 = (~(T9tyx6 & Cn77z6));
assign T9tyx6 = (~(Cflhy6 | Kflhy6));
assign Cflhy6 = (~(Gpeiy6 & Hbvyx6));
assign Qoeiy6 = (~(Bqp7z6[30] & D5qyx6));
assign Cneiy6 = (Opeiy6 & Wpeiy6);
assign Wpeiy6 = (Eqeiy6 & Mqeiy6);
assign Mqeiy6 = (~(E6p7z6[30] & L9qyx6));
assign Eqeiy6 = (~(B2q7z6[30] & Fcqyx6));
assign Opeiy6 = (Uqeiy6 & Creiy6);
assign Creiy6 = (~(Mkp7z6[30] & Tdqyx6));
assign Uqeiy6 = (~(Hfqyx6 & U9p7z6[30]));
assign Emeiy6 = (Kreiy6 & Sreiy6);
assign Sreiy6 = (~(Aseiy6 & U2jhy6));
assign U2jhy6 = (Ptbiw6 & Klo7z6[5]);
assign Aseiy6 = (Iseiy6 & K3jhy6);
assign K3jhy6 = (T9uyx6 | Nsoyx6);
assign Nsoyx6 = (~(Vociw6 | Qseiy6));
assign Qseiy6 = (!Rmget6);
assign Vociw6 = (T59iw6 | Dtj7z6[2]);
assign T9uyx6 = (Ptbiw6 & Rmget6);
assign Ptbiw6 = (!Rediw6);
assign Rediw6 = (~(Dtj7z6[2] & Yseiy6));
assign Yseiy6 = (~(T59iw6 ^ Q9eiw6));
assign Q9eiw6 = (Dtj7z6[4] & Dtj7z6[3]);
assign T59iw6 = (!Dtj7z6[5]);
assign Iseiy6 = (~(Gteiy6 & Oteiy6));
assign Oteiy6 = (Wteiy6 & Eueiy6);
assign Eueiy6 = (Mueiy6 & Uueiy6);
assign Uueiy6 = (~(Hyj7z6[3] & B6diw6));
assign Mueiy6 = (~(Hyj7z6[2] & U5diw6));
assign Wteiy6 = (Cveiy6 & Kveiy6);
assign Kveiy6 = (~(Hyj7z6[1] & N5diw6));
assign Cveiy6 = (~(Hyj7z6[5] & I6diw6));
assign Gteiy6 = (Sveiy6 & Aweiy6);
assign Aweiy6 = (Iweiy6 & Qweiy6);
assign Qweiy6 = (~(Hyj7z6[6] & P6diw6));
assign Iweiy6 = (~(Hyj7z6[7] & W6diw6));
assign Sveiy6 = (Yweiy6 & Gxeiy6);
assign Gxeiy6 = (~(Hyj7z6[0] & Dfk7z6[30]));
assign Yweiy6 = (~(Hyj7z6[4] & Jkl7z6[30]));
assign Kreiy6 = (~(Klo7z6[2] & Oxeiy6));
assign Oxeiy6 = (~(Wxeiy6 & Eyeiy6));
assign Eyeiy6 = (Myeiy6 & Uyeiy6);
assign Uyeiy6 = (~(Dto7z6[0] & Y7kiw6));
assign Y7kiw6 = (Czeiy6 & Z4p7z6[0]);
assign Czeiy6 = (!Kzeiy6);
assign Myeiy6 = (Szeiy6 & A0fiy6);
assign A0fiy6 = (~(Wvo7z6[0] & K7kiw6));
assign K7kiw6 = (~(Kzeiy6 | Z4p7z6[0]));
assign Kzeiy6 = (~(I0fiy6 & Q0fiy6));
assign I0fiy6 = (Z4p7z6[2] & Z4p7z6[1]);
assign Szeiy6 = (~(Pyo7z6[0] & W6kiw6));
assign W6kiw6 = (Y0fiy6 & Pfuyx6);
assign Y0fiy6 = (Q0fiy6 & Z4p7z6[0]);
assign Wxeiy6 = (G1fiy6 & O1fiy6);
assign O1fiy6 = (~(I1p7z6[0] & I6kiw6));
assign I6kiw6 = (W1fiy6 & Pfuyx6);
assign Pfuyx6 = (~(R2syx6 | Z4p7z6[1]));
assign W1fiy6 = (Q0fiy6 & Hfuyx6);
assign G1fiy6 = (E2fiy6 & M2fiy6);
assign M2fiy6 = (~(Ws1ft6 & U5kiw6));
assign U5kiw6 = (U2fiy6 & A0phy6);
assign U2fiy6 = (Z4p7z6[1] & Z4p7z6[0]);
assign E2fiy6 = (~(Nw1ft6 & G5kiw6));
assign G5kiw6 = (C3fiy6 & A0phy6);
assign A0phy6 = (Q0fiy6 & R2syx6);
assign R2syx6 = (!Z4p7z6[2]);
assign Q0fiy6 = (K3fiy6 & Z4p7z6[4]);
assign K3fiy6 = (~(Z4p7z6[3] | Z4p7z6[5]));
assign C3fiy6 = (Z4p7z6[1] & Hfuyx6);
assign Hfuyx6 = (!Z4p7z6[0]);
assign Oleiy6 = (S3fiy6 & O53iy6);
assign O53iy6 = (Qg3iy6 & A4fiy6);
assign A4fiy6 = (~(C7xhy6 & D1pyx6));
assign D1pyx6 = (~(Otshy6 | I4fiy6));
assign C7xhy6 = (W5qhy6 & J2xyx6);
assign Qg3iy6 = (~(F0pyx6 & Q4fiy6));
assign Q4fiy6 = (~(Pntyx6 & Xntyx6));
assign Xntyx6 = (Kr0iy6 & Y4fiy6);
assign Y4fiy6 = (~(G5fiy6 & Ti2nz6[1]));
assign G5fiy6 = (~(O5fiy6 | Ti2nz6[2]));
assign Kr0iy6 = (S7xhy6 | Z6wyx6);
assign Pntyx6 = (W5fiy6 & E6fiy6);
assign E6fiy6 = (Q0mhy6 | O5fiy6);
assign Q0mhy6 = (!O1mhy6);
assign O1mhy6 = (R2uyx6 & Bmvyx6);
assign Bmvyx6 = (!Ti2nz6[2]);
assign W5fiy6 = (Gtshy6 & Cr0iy6);
assign Cr0iy6 = (O5fiy6 | Z6wyx6);
assign Z6wyx6 = (~(Ti2nz6[2] & R2uyx6));
assign R2uyx6 = (!Ti2nz6[1]);
assign O5fiy6 = (~(M6fiy6 & U6fiy6));
assign M6fiy6 = (Ti2nz6[4] & Ti2nz6[0]);
assign Gtshy6 = (S7xhy6 | Ti2nz6[2]);
assign S7xhy6 = (~(C7fiy6 & U6fiy6));
assign U6fiy6 = (~(Ti2nz6[3] | Ti2nz6[5]));
assign C7fiy6 = (Ti2nz6[4] & B2uyx6);
assign B2uyx6 = (!Ti2nz6[0]);
assign F0pyx6 = (~(Oduhy6 | I4fiy6));
assign S3fiy6 = (K7fiy6 & S7fiy6);
assign S7fiy6 = (~(A8fiy6 & Ngqyx6));
assign A8fiy6 = (~(I8fiy6 & Q8fiy6));
assign Q8fiy6 = (Y8fiy6 & G9fiy6);
assign G9fiy6 = (O9fiy6 & W9fiy6);
assign W9fiy6 = (Eafiy6 & Ea0iy6);
assign Ea0iy6 = (U2vhy6 & Ywwhy6);
assign Ywwhy6 = (~(C3eiy6 & Hjsyx6));
assign U2vhy6 = (~(C3eiy6 & Voqyx6));
assign C3eiy6 = (Dlqyx6 & Wtciy6);
assign Eafiy6 = (Mafiy6 & Uafiy6);
assign Uafiy6 = (~(Hjsyx6 & Cbfiy6));
assign Cbfiy6 = (~(Kbfiy6 & Sbfiy6));
assign Sbfiy6 = (~(Nksyx6 & Gaj7z6[1]));
assign Nksyx6 = (!Knohy6);
assign Knohy6 = (~(Acfiy6 & Wtciy6));
assign Kbfiy6 = (~(Byi7z6[30] & Zisyx6));
assign Mafiy6 = (~(Wui7z6[30] & Lxqyx6));
assign Lxqyx6 = (Xryyx6 & Icfiy6);
assign Icfiy6 = (~(Tlqyx6 & Zyuyx6));
assign O9fiy6 = (Qcfiy6 & Ycfiy6);
assign Ycfiy6 = (Gdfiy6 & Odfiy6);
assign Odfiy6 = (~(Dri7z6[30] & Fwqyx6));
assign Fwqyx6 = (~(E28iy6 | Zyuyx6));
assign E28iy6 = (~(Wdfiy6 & Qw2iy6));
assign Qw2iy6 = (Y08iy6 & Koaiw6);
assign Y08iy6 = (Wtciy6 & Toi7z6[6]);
assign Wdfiy6 = (Toi7z6[5] & Toi7z6[7]);
assign Gdfiy6 = (~(Bwi7z6[30] & Hzqyx6));
assign Hzqyx6 = (Xryyx6 & Hjsyx6);
assign Xryyx6 = (Eefiy6 & Mefiy6);
assign Eefiy6 = (Koaiw6 & Wtciy6);
assign Qcfiy6 = (Uefiy6 & Cffiy6);
assign Cffiy6 = (~(Ba0zx6 & T7j7z6[1]));
assign Ba0zx6 = (~(Ua0iy6 | Hzuyx6));
assign Ua0iy6 = (!Zisyx6);
assign Zisyx6 = (Kffiy6 & Wtciy6);
assign Uefiy6 = (~(Svkhy6 & Pnb7z6[30]));
assign Svkhy6 = (Sffiy6 & Dlqyx6);
assign Sffiy6 = (Wtciy6 & Jmqyx6);
assign Wtciy6 = (Agfiy6 & Igfiy6);
assign Agfiy6 = (Qgfiy6 & Ygfiy6);
assign Y8fiy6 = (Ghfiy6 & Ohfiy6);
assign Ohfiy6 = (Whfiy6 & Eifiy6);
assign Eifiy6 = (Mifiy6 & Uifiy6);
assign Uifiy6 = (~(D90zx6 & Lgj7z6[190]));
assign D90zx6 = (~(Cjfiy6 | I08iy6));
assign Mifiy6 = (~(Za0zx6 & Lgj7z6[178]));
assign Za0zx6 = (Kjfiy6 & Jmqyx6);
assign Kjfiy6 = (!Cjfiy6);
assign Whfiy6 = (Sjfiy6 & Akfiy6);
assign Akfiy6 = (~(Hb0zx6 & Lgj7z6[166]));
assign Hb0zx6 = (~(Cjfiy6 | Tlqyx6));
assign Sjfiy6 = (~(Vc0zx6 & Lgj7z6[154]));
assign Vc0zx6 = (~(Cjfiy6 | Hzuyx6));
assign Cjfiy6 = (~(Ikfiy6 & Mefiy6));
assign Mefiy6 = (Qkfiy6 & Toi7z6[5]);
assign Ikfiy6 = (Ykfiy6 & Koaiw6);
assign Ghfiy6 = (Glfiy6 & Olfiy6);
assign Olfiy6 = (Wlfiy6 & Emfiy6);
assign Emfiy6 = (~(Dd0zx6 & Lgj7z6[142]));
assign Dd0zx6 = (~(Mmfiy6 | I08iy6));
assign Wlfiy6 = (~(Be0zx6 & Lgj7z6[130]));
assign Be0zx6 = (~(Mmfiy6 | Zyuyx6));
assign Zyuyx6 = (!Jmqyx6);
assign Glfiy6 = (Umfiy6 & Cnfiy6);
assign Cnfiy6 = (~(Je0zx6 & Lgj7z6[118]));
assign Je0zx6 = (~(Mmfiy6 | Tlqyx6));
assign Umfiy6 = (~(Bi0zx6 & Lgj7z6[106]));
assign Bi0zx6 = (~(Mmfiy6 | Hzuyx6));
assign Mmfiy6 = (~(Ykfiy6 & Kffiy6));
assign Kffiy6 = (Knfiy6 & Qkfiy6);
assign Knfiy6 = (Toi7z6[5] & Tpyyx6);
assign I8fiy6 = (Snfiy6 & Aofiy6);
assign Aofiy6 = (Iofiy6 & Qofiy6);
assign Qofiy6 = (Yofiy6 & Gpfiy6);
assign Gpfiy6 = (Opfiy6 & Wpfiy6);
assign Wpfiy6 = (~(Ji0zx6 & Lgj7z6[94]));
assign Ji0zx6 = (~(Eqfiy6 | I08iy6));
assign Opfiy6 = (~(Dh0zx6 & Lgj7z6[82]));
assign Dh0zx6 = (Mqfiy6 & Jmqyx6);
assign Yofiy6 = (Uqfiy6 & Crfiy6);
assign Crfiy6 = (~(Hj0zx6 & Lgj7z6[70]));
assign Hj0zx6 = (~(Eqfiy6 | Tlqyx6));
assign Uqfiy6 = (~(Pj0zx6 & Lgj7z6[58]));
assign Pj0zx6 = (~(Eqfiy6 | Hzuyx6));
assign Hzuyx6 = (!Voqyx6);
assign Eqfiy6 = (!Mqfiy6);
assign Mqfiy6 = (Ykfiy6 & Acfiy6);
assign Iofiy6 = (Krfiy6 & Srfiy6);
assign Srfiy6 = (Asfiy6 & Isfiy6);
assign Isfiy6 = (~(Dl0zx6 & Lgj7z6[46]));
assign Dl0zx6 = (Qsfiy6 & Ykfiy6);
assign Qsfiy6 = (Hjsyx6 & Dlqyx6);
assign Asfiy6 = (~(Ll0zx6 & Lgj7z6[34]));
assign Ll0zx6 = (Xzuyx6 & Ykfiy6);
assign Xzuyx6 = (Dlqyx6 & Jmqyx6);
assign Jmqyx6 = (Ysfiy6 & Pb8iw6);
assign Krfiy6 = (Gtfiy6 & Otfiy6);
assign Otfiy6 = (~(Jm0zx6 & Lgj7z6[22]));
assign Jm0zx6 = (Wtfiy6 & Ykfiy6);
assign Wtfiy6 = (Lpyyx6 & Dlqyx6);
assign Lpyyx6 = (!Tlqyx6);
assign Gtfiy6 = (~(Rm0zx6 & Lgj7z6[10]));
assign Rm0zx6 = (Eufiy6 & Ykfiy6);
assign Ykfiy6 = (~(Mufiy6 | Uufiy6));
assign Mufiy6 = (Je2iw6 | Cvfiy6);
assign Je2iw6 = (!Lxbet6);
assign Eufiy6 = (Voqyx6 & Dlqyx6);
assign Snfiy6 = (Kvfiy6 & Svfiy6);
assign Svfiy6 = (Awfiy6 & Iwfiy6);
assign Iwfiy6 = (Qwfiy6 & Ywfiy6);
assign Ywfiy6 = (~(Pzqyx6 & G5j7z6[62]));
assign Pzqyx6 = (~(Gxfiy6 | Tlqyx6));
assign Qwfiy6 = (~(Jyqyx6 & G5j7z6[30]));
assign Jyqyx6 = (Oxfiy6 & Voqyx6);
assign Oxfiy6 = (!Gxfiy6);
assign Gxfiy6 = (~(Wxfiy6 & Eyfiy6));
assign Eyfiy6 = (Myfiy6 & Igfiy6);
assign Wxfiy6 = (Dlqyx6 & Ealhy6);
assign Dlqyx6 = (Uyfiy6 & Qkfiy6);
assign Uyfiy6 = (Tpyyx6 & E32nv6);
assign Awfiy6 = (Czfiy6 & Kzfiy6);
assign Kzfiy6 = (~(B2ryx6 & M6j7z6[62]));
assign B2ryx6 = (~(Szfiy6 | Tlqyx6));
assign Czfiy6 = (~(J2ryx6 & M6j7z6[30]));
assign J2ryx6 = (A0giy6 & Voqyx6);
assign A0giy6 = (!Szfiy6);
assign Szfiy6 = (~(I0giy6 & Q0giy6));
assign Q0giy6 = (Tpyyx6 & Malhy6);
assign I0giy6 = (~(Pdm7x6 | Ygfiy6));
assign Kvfiy6 = (Y0giy6 & G1giy6);
assign G1giy6 = (~(STCALIB[24] & F4ryx6));
assign F4ryx6 = (~(Lxuyx6 | I08iy6));
assign I08iy6 = (!Hjsyx6);
assign Hjsyx6 = (Ysfiy6 & Toi7z6[2]);
assign Lxuyx6 = (!Noqyx6);
assign Noqyx6 = (Acfiy6 & Vkqyx6);
assign Vkqyx6 = (~(Uufiy6 | Toi7z6[10]));
assign Uufiy6 = (~(O1giy6 & Malhy6));
assign O1giy6 = (~(Ealhy6 | Toi7z6[11]));
assign Acfiy6 = (W1giy6 & Koaiw6);
assign W1giy6 = (Qkfiy6 & E32nv6);
assign Y0giy6 = (E2giy6 & M2giy6);
assign M2giy6 = (~(D1ryx6 & Ohj7z6[62]));
assign D1ryx6 = (~(U2giy6 | Tlqyx6));
assign Tlqyx6 = (~(C3giy6 & Lxbet6));
assign C3giy6 = (Toi7z6[2] & K3giy6);
assign E2giy6 = (~(X3ryx6 & Ohj7z6[30]));
assign X3ryx6 = (S3giy6 & Voqyx6);
assign Voqyx6 = (K3giy6 & Pb8iw6);
assign K3giy6 = (!Ysfiy6);
assign Ysfiy6 = (Lxbet6 & Toi7z6[3]);
assign S3giy6 = (!U2giy6);
assign U2giy6 = (~(A4giy6 & I4giy6));
assign I4giy6 = (Tpyyx6 & Ygfiy6);
assign Ygfiy6 = (!Ealhy6);
assign Ealhy6 = (Lxbet6 & Toi7z6[9]);
assign Tpyyx6 = (!Koaiw6);
assign Koaiw6 = (Lxbet6 & Toi7z6[4]);
assign A4giy6 = (~(Pdm7x6 | Malhy6));
assign Malhy6 = (!Igfiy6);
assign Igfiy6 = (Lxbet6 & Toi7z6[8]);
assign Pdm7x6 = (~(Myfiy6 & Q4giy6));
assign Q4giy6 = (~(Toi7z6[5] | Toi7z6[6]));
assign Myfiy6 = (~(Toi7z6[10] | Toi7z6[11]));
assign K7fiy6 = (~(Ies7z6[30] & Tltyx6));
assign Tltyx6 = (Y4giy6 & Klo7z6[0]);
assign Y4giy6 = (Hfryx6 & Pfryx6);
assign Ykeiy6 = (~(Dtm7z6[3] & Agdiy6));
assign Ikeiy6 = (G5giy6 & O5giy6);
assign O5giy6 = (~(Dtm7z6[0] & HRDATAD[30]));
assign G5giy6 = (~(Dtm7z6[1] & HRDATAS[30]));
assign Kjeiy6 = (~(L8wnv6 & Itb7z6[30]));
assign L8wnv6 = (~(Fvd7x6 | G9wnv6));
assign G9wnv6 = (Ahe7x6 & W5giy6);
assign W5giy6 = (~(Ohe7x6 & E6giy6));
assign E6giy6 = (~(Ugo7z6[1] & Ncf7x6));
assign Ncf7x6 = (M6giy6 ? Ugo7z6[0] : Jie7x6);
assign Ahe7x6 = (~(Aglov6 | L3bdt6));
assign Fvd7x6 = (U6giy6 & L3bdt6);
assign U6giy6 = (~(T5wnv6 | A6wnv6));
assign T5wnv6 = (~(C7giy6 & Q7wnv6));
assign C7giy6 = (Dx1iw6 | K7giy6);
assign Dx1iw6 = (~(S7giy6 & A8giy6));
assign A8giy6 = (~(HREADYD & Vm1ov6));
assign S7giy6 = (I8giy6 & Q8giy6);
assign Q8giy6 = (~(Y8giy6 & Ee3iw6));
assign Y8giy6 = (M52iw6 & Vd2iw6);
assign I8giy6 = (~(Fk9ov6 & HREADYS));
assign Mho7v6 = (!Yp5xx6);
assign Yp5xx6 = (G9giy6 & O9giy6);
assign O9giy6 = (~(J5exx6 & Bgt8v6));
assign J5exx6 = (W9giy6 & W26xx6);
assign W26xx6 = (!T51nz6[2]);
assign G9giy6 = (T51nz6[2] ? Magiy6 : Eagiy6);
assign Magiy6 = (~(Bgt8v6 ^ W9giy6));
assign Eagiy6 = (Bgt8v6 | W9giy6);
assign W9giy6 = (!T3exx6);
assign T3exx6 = (~(Uagiy6 & Cbgiy6));
assign Cbgiy6 = (~(Ei9xx6 & Kbgiy6));
assign Kbgiy6 = (~(Zi9xx6 & P26xx6));
assign P26xx6 = (!T51nz6[1]);
assign Zi9xx6 = (!Let8v6);
assign Ei9xx6 = (T51nz6[0] & Wsc7v6);
assign Wsc7v6 = (~(Sbgiy6 & Acgiy6));
assign Acgiy6 = (Icgiy6 & Kkaxx6);
assign Kkaxx6 = (~(Mt9xx6 & Ztb7v6));
assign Mt9xx6 = (!Zp9xx6);
assign Icgiy6 = (~(Qcgiy6 & Ycgiy6));
assign Ycgiy6 = (~(Gdgiy6 & Oiexx6));
assign Oiexx6 = (!Gnzmz6[39]);
assign Gdgiy6 = (Odgiy6 | Wdgiy6);
assign Wdgiy6 = (Eegiy6 & Lrexx6);
assign Sbgiy6 = (Megiy6 & Uegiy6);
assign Uegiy6 = (~(Cfgiy6 & Dl9xx6));
assign Cfgiy6 = (~(Kfgiy6 | Sfgiy6));
assign Kfgiy6 = (Pssnv6 & Aggiy6);
assign Pssnv6 = (!B0snv6);
assign Megiy6 = (B0snv6 ? Zp9xx6 : Cuaxx6);
assign Uagiy6 = (~(T51nz6[1] & Let8v6));
assign Let8v6 = (~(Iggiy6 & Qggiy6));
assign Qggiy6 = (Yggiy6 & Ghgiy6);
assign Ghgiy6 = (~(Ohgiy6 & Whgiy6));
assign Whgiy6 = (Eigiy6 | Sfgiy6);
assign Yggiy6 = (~(Fsaxx6 & B0snv6));
assign Fsaxx6 = (!Cuaxx6);
assign Cuaxx6 = (J4snv6 | Migiy6);
assign Iggiy6 = (Uigiy6 & Cjgiy6);
assign Cjgiy6 = (~(Qcgiy6 & Kjgiy6));
assign Kjgiy6 = (~(Sjgiy6 ^ Odgiy6));
assign Bgt8v6 = (Akgiy6 | Ikgiy6);
assign Ikgiy6 = (C5exx6 ? Ohgiy6 : V4exx6);
assign C5exx6 = (~(Qkgiy6 & Ykgiy6));
assign Ykgiy6 = (~(Glgiy6 & Yodxx6));
assign Qkgiy6 = (Olgiy6 & Wlgiy6);
assign Ohgiy6 = (Dl9xx6 & Emgiy6);
assign Emgiy6 = (~(Sfgiy6 & Eigiy6));
assign V4exx6 = (Mmgiy6 & Dl9xx6);
assign Dl9xx6 = (~(Migiy6 | H2tnv6));
assign H2tnv6 = (!J4snv6);
assign J4snv6 = (~(Ztb7v6 & Fgzmz6[0]));
assign Migiy6 = (~(Umgiy6 & Cngiy6));
assign Cngiy6 = (Kngiy6 & Uzrnv6);
assign Uzrnv6 = (!Fgzmz6[1]);
assign Umgiy6 = (~(Lp9xx6 | Hbb7v6));
assign Lp9xx6 = (!I0snv6);
assign Mmgiy6 = (Sfgiy6 & Eigiy6);
assign Eigiy6 = (~(Sngiy6 & Aogiy6));
assign Aogiy6 = (~(Iogiy6 & Y6axx6));
assign Iogiy6 = (Taexx6 & Wlgiy6);
assign Sngiy6 = (Qogiy6 & Jqexx6);
assign Jqexx6 = (!Nfdxx6);
assign Nfdxx6 = (~(Toexx6 | Yodxx6));
assign Qogiy6 = (~(Yogiy6 & Ynexx6));
assign Yogiy6 = (Yodxx6 & Gpgiy6);
assign Gpgiy6 = (~(Wlgiy6 & Lmcxx6));
assign Wlgiy6 = (!Mhexx6);
assign Sfgiy6 = (Opgiy6 & B0snv6);
assign B0snv6 = (~(Wpgiy6 & Eqgiy6));
assign Eqgiy6 = (~(Mqgiy6 & Uqgiy6));
assign Uqgiy6 = (~(Crgiy6 & Uctnv6));
assign Crgiy6 = (Sgbxx6 & Idtnv6);
assign Mqgiy6 = (~(Krgiy6 & Srgiy6));
assign Srgiy6 = (Asgiy6 & Isgiy6);
assign Isgiy6 = (Qsgiy6 & Izsnv6);
assign Izsnv6 = (!Bba7v6);
assign Qsgiy6 = (~(Mbc7v6 | I9b7v6));
assign Asgiy6 = (Jjrnv6 & A04xx6);
assign Jjrnv6 = (~(A377v6 & Wnqnv6));
assign Wnqnv6 = (Ipymz6[0] & Fpqnv6);
assign Fpqnv6 = (!Ipymz6[1]);
assign Krgiy6 = (Ysgiy6 & Gtgiy6);
assign Gtgiy6 = (Otgiy6 & Fgzmz6[0]);
assign Otgiy6 = (Wtgiy6 & Eugiy6);
assign Eugiy6 = (~(Mugiy6 & Uugiy6));
assign Uugiy6 = (Lczmz6[1] & Cvgiy6);
assign Cvgiy6 = (~(Idtnv6 & Detnv6));
assign Mugiy6 = (Lczmz6[3] & Lczmz6[2]);
assign Wtgiy6 = (~(W9c7v6 & H8c7v6));
assign Ysgiy6 = (Kvgiy6 & Tz3xx6);
assign Kvgiy6 = (Qxb7v6 ? Awgiy6 : Svgiy6);
assign Awgiy6 = (~(Iwgiy6 & Qwgiy6));
assign Iwgiy6 = (Zvaxx6 & Kngiy6);
assign Zvaxx6 = (!Ro87v6);
assign Svgiy6 = (~(Tf87v6 & K1snv6));
assign K1snv6 = (!De87v6);
assign Wpgiy6 = (~(Pdtnv6 | Ifb7v6));
assign Pdtnv6 = (Tkb7v6 & Bdtnv6);
assign Bdtnv6 = (!Bhb7v6);
assign Opgiy6 = (!Aggiy6);
assign Aggiy6 = (Ywgiy6 ^ Gxgiy6);
assign Gxgiy6 = (Lmcxx6 ^ Glexx6);
assign Glexx6 = (!Maexx6);
assign Maexx6 = (~(Hpexx6 | Mhexx6));
assign Mhexx6 = (Yodxx6 & Y9exx6);
assign Y9exx6 = (~(Oxgiy6 & Wxgiy6));
assign Wxgiy6 = (Eygiy6 & Ibbxx6);
assign Ibbxx6 = (!Pazmz6[6]);
assign Eygiy6 = (~(Pazmz6[7] | Pazmz6[8]));
assign Oxgiy6 = (~(Pazmz6[4] | Pazmz6[5]));
assign Hpexx6 = (!Yodxx6);
assign Yodxx6 = (Cdb7v6 & Rmb7v6);
assign Lmcxx6 = (!Dz9xx6);
assign Dz9xx6 = (Jezmz6[31] & Ro87v6);
assign Ywgiy6 = (Mygiy6 ^ Y6axx6);
assign Y6axx6 = (Jezmz6[7] & Ro87v6);
assign Mygiy6 = (~(Uygiy6 & Toexx6));
assign Toexx6 = (!Skexx6);
assign Skexx6 = (~(Taexx6 | Ynexx6));
assign Uygiy6 = (~(Czgiy6 & Taexx6));
assign Taexx6 = (!Glgiy6);
assign Glgiy6 = (Jezmz6[15] & Ro87v6);
assign Czgiy6 = (~(Ro87v6 & Olgiy6));
assign Olgiy6 = (!Ynexx6);
assign Ynexx6 = (Jezmz6[23] & Ro87v6);
assign Akgiy6 = (~(Uigiy6 & Kzgiy6));
assign Kzgiy6 = (~(Qcgiy6 & Szgiy6));
assign Szgiy6 = (Sjgiy6 | Odgiy6);
assign Odgiy6 = (~(Lrexx6 | Eegiy6));
assign Eegiy6 = (A0hiy6 ^ Ueexx6);
assign Ueexx6 = (!Gnzmz6[23]);
assign Lrexx6 = (!Gnzmz6[31]);
assign Sjgiy6 = (~(I0hiy6 & Q0hiy6));
assign Q0hiy6 = (~(Gnzmz6[23] & A0hiy6));
assign A0hiy6 = (B987v6 ^ Gnzmz6[15]);
assign I0hiy6 = (~(B987v6 & Gnzmz6[15]));
assign Uigiy6 = (Y0hiy6 & Zp9xx6);
assign Zp9xx6 = (~(G1hiy6 & Z24xx6));
assign Z24xx6 = (~(Hbb7v6 | Fgzmz6[1]));
assign G1hiy6 = (Oob7v6 & I0snv6);
assign Y0hiy6 = (~(Gnzmz6[39] & Qcgiy6));
assign Qcgiy6 = (~(I0snv6 | Ka87v6));
assign I0snv6 = (~(O1hiy6 & W1hiy6));
assign W1hiy6 = (E2hiy6 & Uctnv6);
assign E2hiy6 = (X3tnv6 & Qch7v6);
assign X3tnv6 = (Bke8x6 & O04xx6);
assign O04xx6 = (!Tftnv6);
assign Tftnv6 = (M2hiy6 & Fgzmz6[0]);
assign M2hiy6 = (Qxb7v6 & Kngiy6);
assign Kngiy6 = (!Oob7v6);
assign Bke8x6 = (!Mftnv6);
assign Mftnv6 = (Kkd7v6 & N6dov6);
assign N6dov6 = (C4dov6 & Jrqnv6);
assign C4dov6 = (~(Y9rnv6 & U2hiy6));
assign U2hiy6 = (~(C3hiy6 & K3hiy6));
assign K3hiy6 = (S3hiy6 & A4hiy6);
assign A4hiy6 = (~(I4hiy6 | H71nz6[6]));
assign I4hiy6 = (H71nz6[7] | H71nz6[8]);
assign S3hiy6 = (~(H71nz6[4] | H71nz6[5]));
assign C3hiy6 = (Q4hiy6 & Y4hiy6);
assign Y4hiy6 = (~(H71nz6[2] | H71nz6[3]));
assign Q4hiy6 = (~(H71nz6[0] | H71nz6[1]));
assign Y9rnv6 = (!Gernv6);
assign Gernv6 = (Qc77v6 & Jrqnv6);
assign Jrqnv6 = (!C477v6);
assign O1hiy6 = (De87v6 & Tf87v6);
assign Kgo7v6 = (~(Aiadt6 | Gonov6));
assign Pfo7v6 = (!Cpsnv6);
assign Ueo7v6 = (!Eqlnv6);
assign Eqlnv6 = (G5hiy6 & O5hiy6);
assign O5hiy6 = (W5hiy6 & E6hiy6);
assign E6hiy6 = (Jsaov6 & Kb9iw6);
assign Kb9iw6 = (!Dysiw6);
assign Dysiw6 = (Lyknv6 & Gvvnv6);
assign Jsaov6 = (M6hiy6 | Dwb7z6[5]);
assign W5hiy6 = (Zyxxx6 & L0bov6);
assign Zyxxx6 = (~(U6hiy6 & Aqihw6));
assign G5hiy6 = (C7hiy6 & K7hiy6);
assign K7hiy6 = (S7hiy6 & Gpmov6);
assign Gpmov6 = (~(Lna7x6 & Ywaov6));
assign S7hiy6 = (~(A8hiy6 & Bhoov6));
assign A8hiy6 = (Xfa7x6 & Fxaov6);
assign C7hiy6 = (I8hiy6 & Q8hiy6);
assign Q8hiy6 = (~(G6xiw6 & Y8hiy6));
assign G6xiw6 = (~(T4jnv6 | Ecc7z6[11]));
assign I8hiy6 = (Ecc7z6[11] ? O9hiy6 : G9hiy6);
assign O9hiy6 = (Y8hiy6 | T4jnv6);
assign Y8hiy6 = (~(Yioov6 & Zayxx6));
assign Zayxx6 = (!Mwphw6);
assign G9hiy6 = (W9hiy6 & Eahiy6);
assign Eahiy6 = (~(Mahiy6 & Fxaov6));
assign W9hiy6 = (~(Wnihw6 | Pi9ov6));
assign Wnihw6 = (Uahiy6 & Ywaov6);
assign Uahiy6 = (Fulnv6 & Uvvnv6);
assign Neo7v6 = (Dte7z6[9] & Fhc7z6[31]);
assign Geo7v6 = (~(Cbhiy6 | Fre7z6[1]));
assign Cbhiy6 = (~(Kbhiy6 | Fre7z6[0]));
assign Kbhiy6 = (~(Onf7z6[31] ^ Elgdt6));
assign Zdo7v6 = (Sbhiy6 & Fflov6);
assign Fflov6 = (Achiy6 & Opd7x6);
assign Opd7x6 = (!Dkeiw6);
assign Dkeiw6 = (~(Ichiy6 & Qchiy6));
assign Qchiy6 = (~(Fvb7z6[13] & M52iw6));
assign Ichiy6 = (~(Se3iw6 & Cmm7z6[13]));
assign Achiy6 = (Oteiw6 & Jrhiw6);
assign Jrhiw6 = (~(Ychiy6 & Gdhiy6));
assign Gdhiy6 = (~(Fvb7z6[12] & M52iw6));
assign Ychiy6 = (~(Se3iw6 & Cmm7z6[12]));
assign Oteiw6 = (Odhiy6 & Kkeiw6);
assign Kkeiw6 = (Wdhiy6 & Vqhiw6);
assign Vqhiw6 = (Eehiy6 & Mehiy6);
assign Mehiy6 = (~(Fvb7z6[16] & M52iw6));
assign Eehiy6 = (~(Se3iw6 & Cmm7z6[16]));
assign Wdhiy6 = (~(Hqhiw6 | Jneiw6));
assign Hqhiw6 = (~(Uehiy6 & Cfhiy6));
assign Cfhiy6 = (~(Fvb7z6[17] & M52iw6));
assign Uehiy6 = (~(Se3iw6 & Cmm7z6[17]));
assign Odhiy6 = (~(Wjeiw6 | Pjeiw6));
assign Pjeiw6 = (~(Kfhiy6 & Sfhiy6));
assign Sfhiy6 = (~(Fvb7z6[14] & M52iw6));
assign Kfhiy6 = (~(Se3iw6 & Cmm7z6[14]));
assign Wjeiw6 = (~(Aghiy6 & Ighiy6));
assign Ighiy6 = (~(Fvb7z6[15] & M52iw6));
assign Aghiy6 = (~(Se3iw6 & Cmm7z6[15]));
assign Sbhiy6 = (~(Da3iw6 | Kygnv6));
assign Sdo7v6 = (~(Da3iw6 | Relov6));
assign Relov6 = (!Jneiw6);
assign Jneiw6 = (P5fov6 | Aqhiw6);
assign Aqhiw6 = (~(Qghiy6 & Yghiy6));
assign Yghiy6 = (~(Fvb7z6[18] & M52iw6));
assign Qghiy6 = (~(Se3iw6 & Cmm7z6[18]));
assign P5fov6 = (~(Ghhiy6 & Ohhiy6));
assign Ohhiy6 = (~(Fvb7z6[19] & M52iw6));
assign Ghhiy6 = (~(Se3iw6 & Cmm7z6[19]));
assign Da3iw6 = (C63iw6 | B23iw6);
assign B23iw6 = (!Iu4ov6);
assign Iu4ov6 = (~(Whhiy6 & Eihiy6));
assign Eihiy6 = (~(Se3iw6 & Hjqnv6));
assign Whhiy6 = (~(K2bdt6 & M52iw6));
assign C63iw6 = (U13iw6 | Pdlov6);
assign Pdlov6 = (!Vd2iw6);
assign U13iw6 = (Mihiy6 & Uihiy6);
assign Uihiy6 = (~(Veonv6 & B2jnv6));
assign Veonv6 = (Ee3iw6 & Se3iw6);
assign Mihiy6 = (~(Ee3iw6 & M52iw6));
assign Edo7v6 = (Fgzmz6[0] & Cjhiy6);
assign Cjhiy6 = (~(Z2vnv6 & A04xx6));
assign A04xx6 = (!Q4c7v6);
assign Z2vnv6 = (!Zz97v6);
assign Zz97v6 = (~(Kjhiy6 & Lqsnv6));
assign Lqsnv6 = (Thh7v6 & Sjhiy6);
assign Sjhiy6 = (~(I9b7v6 & F02nv6));
assign Kjhiy6 = (Akhiy6 & Ikhiy6);
assign Ikhiy6 = (~(Mbc7v6 & Qkhiy6));
assign Qkhiy6 = (~(Ykhiy6 & Glhiy6));
assign Glhiy6 = (Olhiy6 & Idtnv6);
assign Idtnv6 = (!Lczmz6[0]);
assign Olhiy6 = (~(Ztb7v6 | Cdb7v6));
assign Ykhiy6 = (Uctnv6 & Sgbxx6);
assign Sgbxx6 = (!Uib7v6);
assign Uctnv6 = (Wlhiy6 & Tusnv6);
assign Tusnv6 = (!Lczmz6[1]);
assign Wlhiy6 = (Z8cxx6 & Wvcxx6);
assign Wvcxx6 = (!Lczmz6[3]);
assign Z8cxx6 = (!Lczmz6[2]);
assign Akhiy6 = (Sqsnv6 | Tz3xx6);
assign Tz3xx6 = (Emhiy6 & Yc77z6);
assign Sqsnv6 = (~(Qwgiy6 & Mmhiy6));
assign Mmhiy6 = (Ursnv6 | O777v6);
assign Ursnv6 = (!Fs3xx6);
assign Fs3xx6 = (~(Cpsnv6 | W9c7v6));
assign Qwgiy6 = (Gdc7v6 | O777v6);
assign Xco7v6 = (~(Umhiy6 & Cnhiy6));
assign Cnhiy6 = (~(Knhiy6 & Soa7v6));
assign Knhiy6 = (~(Pxunv6 | W1a7v6));
assign Pxunv6 = (I1c7v6 ? Z2c7v6 : Snhiy6);
assign Snhiy6 = (~(Aohiy6 & F8tnv6));
assign Aohiy6 = (~(G197z6 | Gdc7v6));
assign Umhiy6 = (~(Mya7v6 | J2b7v6));
assign J2b7v6 = (!F8tnv6);
assign F8tnv6 = (~(Iohiy6 & A9tnv6));
assign A9tnv6 = (Wfo7v6 & Ldo7v6);
assign Iohiy6 = (I9b7v6 & Kwl8v6);
assign Mya7v6 = (~(Qohiy6 | Emhiy6));
assign Emhiy6 = (!D4b7v6);
assign Qohiy6 = (O9tnv6 | W1a7v6);
assign O9tnv6 = (!Kwl8v6);
assign Kwl8v6 = (~(Yohiy6 | Glh7v6));
assign Qco7v6 = (~(Gphiy6 & Ophiy6));
assign Ophiy6 = (~(HRDATAD[4] & Qln7z6[0]));
assign Gphiy6 = (~(HRDATAS[4] & Qln7z6[1]));
assign Jco7v6 = (~(Wphiy6 & Eqhiy6));
assign Eqhiy6 = (~(HRDATAD[12] & Qln7z6[0]));
assign Wphiy6 = (~(HRDATAS[12] & Qln7z6[1]));
assign Cco7v6 = (~(Mqhiy6 & Uqhiy6));
assign Uqhiy6 = (~(HRDATAD[20] & Qln7z6[0]));
assign Mqhiy6 = (~(HRDATAS[20] & Qln7z6[1]));
assign Obo7v6 = (Crhiy6 & Gjdiw6);
assign Crhiy6 = (Krhiy6 & Lgonv6);
assign Krhiy6 = (~(Srhiy6 & Ashiy6));
assign Ashiy6 = (~(Ishiy6 & Wbhnv6));
assign Ishiy6 = (Cmm7z6[1] & Cmm7z6[0]);
assign Abo7v6 = (!Vstiw6);
assign Vstiw6 = (~(S9tiw6 & Qshiy6));
assign Qshiy6 = (~(Yshiy6 & Gthiy6));
assign Gthiy6 = (Othiy6 & Wthiy6);
assign Wthiy6 = (Kxtiw6 & Z6jhw6);
assign Kxtiw6 = (~(Euhiy6 & Bdf7z6[2]));
assign Euhiy6 = (Muhiy6 & R4aov6);
assign Othiy6 = (Uuhiy6 & Cvhiy6);
assign Cvhiy6 = (~(Hetiw6 & Kvhiy6));
assign Kvhiy6 = (~(Ghtiw6 & Svhiy6));
assign Svhiy6 = (~(Awhiy6 & Go37x6));
assign Awhiy6 = (Iwhiy6 & Xftiw6);
assign Xftiw6 = (~(Qwhiy6 & Mrbdt6));
assign Qwhiy6 = (Ywhiy6 & Cu27x6);
assign Ywhiy6 = (~(Nh2ov6 & Zn37x6));
assign Zn37x6 = (!Kxb7z6[31]);
assign Nh2ov6 = (!Fhc7z6[31]);
assign Ghtiw6 = (Gxhiy6 & Fnfxx6);
assign Fnfxx6 = (!Tk8iw6);
assign Gxhiy6 = (~(Mnfxx6 & Lgtiw6));
assign Lgtiw6 = (~(Entiw6 & Lntiw6));
assign Uuhiy6 = (~(Frtiw6 & Trtiw6));
assign Trtiw6 = (~(Oxhiy6 & Wxhiy6));
assign Wxhiy6 = (~(Eyhiy6 & Myhiy6));
assign Eyhiy6 = (!Qftiw6);
assign Qftiw6 = (Iwhiy6 | Mnfxx6);
assign Oxhiy6 = (~(Xjxxx6 & Go37x6));
assign Go37x6 = (!Entiw6);
assign Entiw6 = (~(Uyhiy6 & Czhiy6));
assign Czhiy6 = (Kzhiy6 & Szhiy6);
assign Szhiy6 = (A0iiy6 & I0iiy6);
assign I0iiy6 = (~(Kxb7z6[8] | Kxb7z6[9]));
assign A0iiy6 = (~(Kxb7z6[6] | Kxb7z6[7]));
assign Kzhiy6 = (Q0iiy6 & Y0iiy6);
assign Y0iiy6 = (~(Kxb7z6[4] | Kxb7z6[5]));
assign Q0iiy6 = (~(Kxb7z6[2] | Kxb7z6[3]));
assign Uyhiy6 = (G1iiy6 & O1iiy6);
assign O1iiy6 = (W1iiy6 & E2iiy6);
assign E2iiy6 = (~(Kxb7z6[15] | Kxb7z6[1]));
assign W1iiy6 = (~(Kxb7z6[13] | Kxb7z6[14]));
assign G1iiy6 = (M2iiy6 & U2iiy6);
assign U2iiy6 = (~(Kxb7z6[11] | Kxb7z6[12]));
assign M2iiy6 = (~(Kxb7z6[0] | Kxb7z6[10]));
assign Xjxxx6 = (~(Mnfxx6 | Myhiy6));
assign Mnfxx6 = (C3iiy6 & K3iiy6);
assign K3iiy6 = (S3iiy6 & A4iiy6);
assign A4iiy6 = (I4iiy6 & Q4iiy6);
assign Q4iiy6 = (~(Kxb7z6[30] | Kxb7z6[31]));
assign I4iiy6 = (~(Kxb7z6[28] | Kxb7z6[29]));
assign S3iiy6 = (Vl37x6 & Tk37x6);
assign Tk37x6 = (~(Kxb7z6[26] | Kxb7z6[27]));
assign Vl37x6 = (~(Kxb7z6[24] | Kxb7z6[25]));
assign C3iiy6 = (Y4iiy6 & G5iiy6);
assign G5iiy6 = (O5iiy6 & Ol37x6);
assign Ol37x6 = (~(Kxb7z6[22] | Kxb7z6[23]));
assign O5iiy6 = (~(Kxb7z6[20] | Kxb7z6[21]));
assign Y4iiy6 = (W5iiy6 & E6iiy6);
assign E6iiy6 = (~(Kxb7z6[18] | Kxb7z6[19]));
assign W5iiy6 = (~(Kxb7z6[16] | Kxb7z6[17]));
assign Frtiw6 = (!A127x6);
assign A127x6 = (~(M6iiy6 & Ngxxx6));
assign M6iiy6 = (Bdf7z6[1] & Ju27x6);
assign Yshiy6 = (U6iiy6 & Dfkov6);
assign Dfkov6 = (~(Y3bov6 | Qf2ov6));
assign Qf2ov6 = (C7iiy6 & Bdf7z6[2]);
assign C7iiy6 = (Bdf7z6[0] & Muhiy6);
assign Y3bov6 = (!Wi2ov6);
assign Wi2ov6 = (~(K7iiy6 & S7iiy6));
assign S7iiy6 = (Bdf7z6[3] & R4aov6);
assign K7iiy6 = (Bdf7z6[2] & Bdf7z6[1]);
assign U6iiy6 = (Bitiw6 & Ts27x6);
assign Ts27x6 = (!Gcmnv6);
assign Gcmnv6 = (~(X927x6 & A8iiy6));
assign A8iiy6 = (~(Notiw6 & R4aov6));
assign X927x6 = (~(I8iiy6 & G427x6));
assign Bitiw6 = (Aofxx6 & Cmtiw6);
assign Cmtiw6 = (Q8iiy6 | K4aov6);
assign Aofxx6 = (~(Uotiw6 & Dqtiw6));
assign Dqtiw6 = (Notiw6 & Bdf7z6[0]);
assign Uotiw6 = (!Zgtiw6);
assign S9tiw6 = (Ozvnv6 & Y8iiy6);
assign Y8iiy6 = (~(Ketnv6 & G9iiy6));
assign G9iiy6 = (~(X3lhw6 & Z6jhw6));
assign Z6jhw6 = (~(O9iiy6 & G427x6));
assign O9iiy6 = (Bdf7z6[3] & D4aov6);
assign X3lhw6 = (~(Yxtiw6 | Hetiw6));
assign Hetiw6 = (!Ilfxx6);
assign Ilfxx6 = (~(W9iiy6 & I8iiy6));
assign I8iiy6 = (D4aov6 & Ju27x6);
assign W9iiy6 = (Bdf7z6[0] & K4aov6);
assign Yxtiw6 = (Ngxxx6 & Muhiy6);
assign Ozvnv6 = (!Dj9ov6);
assign Dj9ov6 = (Tnzdt6 & Ga3nv6);
assign Tao7v6 = (!A4a7z6);
assign A4a7z6 = (~(Eaiiy6 & G4mov6));
assign G4mov6 = (~(Maiiy6 & Uaiiy6));
assign Uaiiy6 = (Cbiiy6 & Kbiiy6);
assign Kbiiy6 = (Sbiiy6 & Aciiy6);
assign Sbiiy6 = (~(L9onv6 | Dpadt6));
assign L9onv6 = (Iciiy6 & Qciiy6);
assign Qciiy6 = (Yciiy6 & Gdiiy6);
assign Gdiiy6 = (Odiiy6 & B5siw6);
assign Odiiy6 = (Zplhw6 & Hcviw6);
assign Yciiy6 = (Wdiiy6 & Rlriw6);
assign Wdiiy6 = (!Mtehw6);
assign Iciiy6 = (Eeiiy6 & Meiiy6);
assign Meiiy6 = (Ueiiy6 & Anriw6);
assign Ueiiy6 = (Cfiiy6 & Kfiiy6);
assign Kfiiy6 = (Q9fhw6 | Sfiiy6);
assign Eeiiy6 = (Siriw6 & K4uiw6);
assign Cbiiy6 = (Chm7x6 & Agiiy6);
assign Agiiy6 = (~(Igiiy6 & Qgiiy6));
assign Qgiiy6 = (~(Ygiiy6 & Ghiiy6));
assign Ygiiy6 = (Ohiiy6 & Fjaov6);
assign Chm7x6 = (~(Fe2nv6 & Ayeet6));
assign Maiiy6 = (Whiiy6 & Eiiiy6);
assign Eiiiy6 = (Miiiy6 & Uiiiy6);
assign Miiiy6 = (Cjiiy6 & Kjiiy6);
assign Kjiiy6 = (~(Sjiiy6 & Vzbet6));
assign Sjiiy6 = (E1cet6 & Amg7x6);
assign Cjiiy6 = (~(Akiiy6 & Ikiiy6));
assign Ikiiy6 = (~(Z147x6 | My37x6));
assign My37x6 = (Qkiiy6 & Ykiiy6);
assign Ykiiy6 = (Gliiy6 & Oliiy6);
assign Oliiy6 = (~(Zec7z6[2] & Wliiy6));
assign Wliiy6 = (~(Siriw6 & Emiiy6));
assign Gliiy6 = (Mmiiy6 & Umiiy6);
assign Umiiy6 = (~(Zec7z6[2] & Cniiy6));
assign Mmiiy6 = (Painv6 | Cfiiy6);
assign Qkiiy6 = (Kniiy6 & Sniiy6);
assign Kniiy6 = (Wcsiw6 & Aoiiy6);
assign Aoiiy6 = (~(Zec7z6[10] & Ioiiy6));
assign Z147x6 = (M547x6 & Qoiiy6);
assign Qoiiy6 = (Yoiiy6 & Gpiiy6);
assign Gpiiy6 = (~(Zec7z6[8] & Opiiy6));
assign Yoiiy6 = (~(Zec7z6[0] & Wpiiy6));
assign Wpiiy6 = (~(Eqiiy6 & Siriw6));
assign Eqiiy6 = (Emiiy6 & I4ghw6);
assign M547x6 = (Sniiy6 & Wcsiw6);
assign Sniiy6 = (~(G5sov6 | Mqiiy6));
assign Akiiy6 = (C047x6 & Uqiiy6);
assign Uqiiy6 = (~(Wcsiw6 & R447x6));
assign C047x6 = (Criiy6 & Kriiy6);
assign Kriiy6 = (Sriiy6 & Amtov6);
assign Sriiy6 = (~(Zec7z6[9] & Opiiy6));
assign Opiiy6 = (~(Cfiiy6 & G3ghw6));
assign Criiy6 = (Asiiy6 & Isiiy6);
assign Isiiy6 = (~(Zec7z6[1] & Qsiiy6));
assign Qsiiy6 = (~(Siriw6 & I4ghw6));
assign Siriw6 = (~(Nxlhw6 | Ysiiy6));
assign Ysiiy6 = (!C3riw6);
assign Whiiy6 = (N3onv6 & Gtiiy6);
assign N3onv6 = (!Vs9ov6);
assign Eaiiy6 = (~(W6u6x6 & Otiiy6));
assign Mao7v6 = (!H2mnv6);
assign H2mnv6 = (~(Wtiiy6 & Euiiy6));
assign Euiiy6 = (Muiiy6 & Pj1ov6);
assign Muiiy6 = (~(Fetov6 & Rdtov6));
assign Rdtov6 = (~(Uuiiy6 & Jamnv6));
assign Uuiiy6 = (Vs9ov6 & A9mnv6);
assign A9mnv6 = (~(Grfxx6 & Cviiy6));
assign Cviiy6 = (~(B8cdt6 & Kviiy6));
assign Kviiy6 = (Sviiy6 | Vmnnv6);
assign Sviiy6 = (Amnnv6 | Awiiy6);
assign Grfxx6 = (Ihaov6 | Ktfxx6);
assign Vs9ov6 = (~(L2o7x6 & X1o7x6));
assign X1o7x6 = (Osa7x6 & Iwiiy6);
assign Iwiiy6 = (Qwiiy6 & S2onv6);
assign Qwiiy6 = (~(Kslov6 & Ywiiy6));
assign Ywiiy6 = (~(Rihov6 & Qg2nv6));
assign Kslov6 = (Vsgov6 & Ga3nv6);
assign Vsgov6 = (Gxiiy6 & Oxiiy6);
assign Oxiiy6 = (~(Wxiiy6 & Eyiiy6));
assign Eyiiy6 = (Kioov6 & Qg2nv6);
assign Wxiiy6 = (Hbo7v6 & Ggoov6);
assign Gxiiy6 = (~(Myiiy6 & Tqinv6));
assign Tqinv6 = (Uyiiy6 & Hbo7v6);
assign Uyiiy6 = (Cziiy6 & Lxydt6);
assign Myiiy6 = (Wxsiw6 & O5a7z6);
assign Wxsiw6 = (!Fiihw6);
assign Osa7x6 = (G3onv6 & W6u6x6);
assign G3onv6 = (Kziiy6 & Sziiy6);
assign Sziiy6 = (A0jiy6 & I0jiy6);
assign I0jiy6 = (~(Tuddt6 | Nneet6));
assign A0jiy6 = (Jnsiw6 & Vzvnv6);
assign Kziiy6 = (Q0jiy6 & Y0jiy6);
assign Y0jiy6 = (Ldo7v6 & D7u6x6);
assign Q0jiy6 = (E1wnv6 & Y7u6x6);
assign Y7u6x6 = (G1jiy6 & O1jiy6);
assign O1jiy6 = (Nneet6 ? E2jiy6 : W1jiy6);
assign E2jiy6 = (~(Ypinv6 | M2jiy6));
assign W1jiy6 = (~(U2jiy6 & W6u6x6));
assign U2jiy6 = (C3jiy6 & Vzvnv6);
assign C3jiy6 = (~(K3jiy6 & S3jiy6));
assign S3jiy6 = (~(A4jiy6 & I4jiy6));
assign I4jiy6 = (Q4jiy6 & Y4jiy6);
assign Y4jiy6 = (~(G5jiy6 & O5jiy6));
assign Q4jiy6 = (W5jiy6 & Qg2nv6);
assign W5jiy6 = (~(E6jiy6 & M6jiy6));
assign A4jiy6 = (S6cdt6 & Rihov6);
assign K3jiy6 = (~(U6jiy6 & I5cdt6));
assign U6jiy6 = (C7jiy6 & K7jiy6);
assign K7jiy6 = (~(H2sov6 & T1sov6));
assign H2sov6 = (!Wpnhw6);
assign C7jiy6 = (~(S6cdt6 & Tnzdt6));
assign G1jiy6 = (I5fov6 ? O5a7z6 : S7jiy6);
assign I5fov6 = (~(Whhov6 | Qg2nv6));
assign S7jiy6 = (~(Zgadt6 & C0wnv6));
assign L2o7x6 = (Jta7x6 & A8jiy6);
assign Jta7x6 = (I8jiy6 & Q8jiy6);
assign Q8jiy6 = (~(Y8jiy6 & G9jiy6));
assign G9jiy6 = (~(O9jiy6 | W9jiy6));
assign Y8jiy6 = (Eajiy6 & Majiy6);
assign Majiy6 = (~(Uajiy6 & Cbjiy6));
assign Uajiy6 = (Kbjiy6 ? Pxfhw6 : Dyfhw6);
assign Eajiy6 = (~(Sbjiy6 & Ixfhw6));
assign Ixfhw6 = (Zofhw6 & Z9nhw6);
assign I8jiy6 = (~(Acjiy6 & Icjiy6));
assign Icjiy6 = (~(Qcjiy6 & W9jiy6));
assign Qcjiy6 = (O9jiy6 & Sbjiy6);
assign Acjiy6 = (W9jiy6 ? Gdjiy6 : Ycjiy6);
assign W9jiy6 = (Odjiy6 & Wdjiy6);
assign Wdjiy6 = (~(Eejiy6 & Xlaov6));
assign Odjiy6 = (~(Mejiy6 & Mzmov6));
assign Gdjiy6 = (Uejiy6 & Cfjiy6);
assign Cfjiy6 = (~(Sbjiy6 & Lcqiw6));
assign Uejiy6 = (Kbjiy6 ? Sfjiy6 : Kfjiy6);
assign Sfjiy6 = (Qgjiy6 ? Igjiy6 : Agjiy6);
assign Igjiy6 = (O9jiy6 ? I6riw6 : P0qiw6);
assign I6riw6 = (!Otfhw6);
assign P0qiw6 = (!Svfhw6);
assign Agjiy6 = (O9jiy6 ? Dmqiw6 : Dnpiw6);
assign Dmqiw6 = (!Vtfhw6);
assign Dnpiw6 = (!Zvfhw6);
assign Kfjiy6 = (Ygjiy6 | Qgjiy6);
assign Qgjiy6 = (!Cbjiy6);
assign Ygjiy6 = (O9jiy6 ? Msfhw6 : Qufhw6);
assign Ycjiy6 = (Ghjiy6 & O9jiy6);
assign O9jiy6 = (Ohjiy6 & Whjiy6);
assign Whjiy6 = (~(Eejiy6 & Kpaov6));
assign Ohjiy6 = (~(Mejiy6 & L2nov6));
assign Ghjiy6 = (Eijiy6 & Mijiy6);
assign Mijiy6 = (~(Uijiy6 & Bqfhw6));
assign Uijiy6 = (Cjjiy6 & Cbjiy6);
assign Eijiy6 = (~(Zofhw6 & Kjjiy6));
assign Kjjiy6 = (~(Sjjiy6 & Akjiy6));
assign Akjiy6 = (~(Ikjiy6 & Kbjiy6));
assign Ikjiy6 = (Cbjiy6 ? Zec7z6[27] : Zec7z6[25]);
assign Sjjiy6 = (~(Sbjiy6 & Zec7z6[24]));
assign Sbjiy6 = (~(Cbjiy6 | Kbjiy6));
assign Kbjiy6 = (!Cjjiy6);
assign Cjjiy6 = (Qkjiy6 & Ykjiy6);
assign Ykjiy6 = (~(Eejiy6 & Pxmov6));
assign Qkjiy6 = (~(Mejiy6 & Gwmov6));
assign Cbjiy6 = (~(Gljiy6 & Oljiy6));
assign Oljiy6 = (~(Eejiy6 & Xumov6));
assign Eejiy6 = (Yl2et6 & Wljiy6);
assign Wljiy6 = (~(Emjiy6 & Mmjiy6));
assign Mmjiy6 = (~(Ltvxx6 & Fulnv6));
assign Gljiy6 = (~(Mejiy6 & Y5nov6));
assign Mejiy6 = (Otsiw6 & Umjiy6);
assign Umjiy6 = (~(Emjiy6 & Tq9iw6));
assign Tq9iw6 = (!Qusiw6);
assign Qusiw6 = (~(Ruvxx6 | Luvnv6));
assign Emjiy6 = (Fiihw6 & Cnjiy6);
assign Cnjiy6 = (~(Ggoov6 & Kioov6));
assign Fiihw6 = (Ayaov6 | Dwb7z6[5]);
assign Wtiiy6 = (O4piw6 & Rihov6);
assign Rihov6 = (Ihaov6 & Qv0ov6);
assign Qv0ov6 = (~(Knjiy6 & Snjiy6));
assign Snjiy6 = (Aojiy6 & Gfihw6);
assign Aojiy6 = (Qdihw6 & Vcihw6);
assign Knjiy6 = (M637x6 & Seihw6);
assign M637x6 = (Iojiy6 & Qojiy6);
assign Qojiy6 = (~(Ypinv6 & Yojiy6));
assign Yojiy6 = (~(Gpjiy6 & Opjiy6));
assign Opjiy6 = (Wpjiy6 & Eqjiy6);
assign Eqjiy6 = (Mqjiy6 & Ajihw6);
assign Mqjiy6 = (Uqjiy6 & Tulnv6);
assign Uqjiy6 = (!Ztaov6);
assign Wpjiy6 = (X1a7x6 & N3a7x6);
assign Gpjiy6 = (Crjiy6 & Krjiy6);
assign Krjiy6 = (Srjiy6 & Asjiy6);
assign Asjiy6 = (~(S2a7x6 & Isjiy6));
assign Srjiy6 = (Qsjiy6 & Qxknv6);
assign Qsjiy6 = (~(Ysjiy6 & Fulnv6));
assign Ysjiy6 = (Dwb7z6[5] & Uvvnv6);
assign Crjiy6 = (At97x6 & Tpxxx6);
assign Tpxxx6 = (~(Ytlnv6 & Gvvnv6));
assign Iojiy6 = (Gtjiy6 & Otjiy6);
assign Otjiy6 = (~(Wtjiy6 & Eujiy6));
assign Eujiy6 = (Mujiy6 & Uujiy6);
assign Uujiy6 = (Cvjiy6 & Kvjiy6);
assign Kvjiy6 = (Svjiy6 & Vcyxx6);
assign Svjiy6 = (Awjiy6 & X1a7x6);
assign Awjiy6 = (!Vpknv6);
assign Vpknv6 = (S2a7x6 & Nvvnv6);
assign Cvjiy6 = (Z2a7x6 & Iwjiy6);
assign Z2a7x6 = (Qwjiy6 | Buvxx6);
assign Qwjiy6 = (!Riuxx6);
assign Mujiy6 = (Ywjiy6 & Gxjiy6);
assign Gxjiy6 = (Oxjiy6 & Wxjiy6);
assign Wxjiy6 = (~(Eyjiy6 & Myjiy6));
assign Myjiy6 = (Uyjiy6 & Czjiy6);
assign Uyjiy6 = (~(Kzjiy6 & Szjiy6));
assign Szjiy6 = (U3a7x6 & A0kiy6);
assign Kzjiy6 = (~(I0kiy6 | Qg2nv6));
assign Eyjiy6 = (Aulov6 & Q0kiy6);
assign Q0kiy6 = (~(Y0kiy6 & G1kiy6));
assign G1kiy6 = (~(Bh2et6 & O1kiy6));
assign O1kiy6 = (~(W1kiy6 & Zdxdt6));
assign W1kiy6 = (~(I0kiy6 | A0kiy6));
assign A0kiy6 = (!O5h7z6[1]);
assign I0kiy6 = (~(E2kiy6 & O5h7z6[2]));
assign E2kiy6 = (O5h7z6[3] & O5h7z6[0]);
assign Y0kiy6 = (~(M2kiy6 & R3h7z6[0]));
assign Aulov6 = (M6a7x6 & Ijmov6);
assign Oxjiy6 = (~(U2kiy6 & X4eet6));
assign U2kiy6 = (Ldmyx6 & C3kiy6);
assign C3kiy6 = (~(K3kiy6 & Qij7z6[4]));
assign K3kiy6 = (~(Qij7z6[0] ^ Qij7z6[1]));
assign Ywjiy6 = (S3kiy6 & A4kiy6);
assign A4kiy6 = (~(I4kiy6 & Whxdt6));
assign I4kiy6 = (Uebdt6 & Czjiy6);
assign Czjiy6 = (Q4kiy6 | M2kiy6);
assign S3kiy6 = (~(Y4kiy6 & Xsinv6));
assign Y4kiy6 = (~(Ix97x6 & Uw97x6));
assign Uw97x6 = (~(Vqihw6 & G5kiy6));
assign Wtjiy6 = (O5kiy6 & W5kiy6);
assign W5kiy6 = (E6kiy6 & M6kiy6);
assign M6kiy6 = (U6kiy6 & C7kiy6);
assign C7kiy6 = (~(K7kiy6 & Lxydt6));
assign K7kiy6 = (~(S7kiy6 & A8kiy6));
assign A8kiy6 = (~(Noa7x6 & Fpphw6));
assign Fpphw6 = (Cwlnv6 & Xdphw6);
assign S7kiy6 = (~(Vxihw6 & I8kiy6));
assign I8kiy6 = (~(Tulnv6 & Q8kiy6));
assign Q8kiy6 = (~(Mwphw6 & Cwlnv6));
assign Mwphw6 = (X4xiw6 & Ecc7z6[10]);
assign X4xiw6 = (Y8kiy6 & G9kiy6);
assign G9kiy6 = (P4c7z6[0] & O9kiy6);
assign Y8kiy6 = (P4c7z6[3] & P4c7z6[2]);
assign U6kiy6 = (~(Remyx6 & W9kiy6));
assign W9kiy6 = (~(Eakiy6 & At97x6));
assign At97x6 = (Makiy6 & Ayaov6);
assign Makiy6 = (~(Uakiy6 & Aqihw6));
assign Aqihw6 = (!Fkyxx6);
assign Fkyxx6 = (Buvxx6 & Bqvxx6);
assign Eakiy6 = (Cbkiy6 & Srknv6);
assign Cbkiy6 = (~(Zzihw6 & Ot97x6));
assign Remyx6 = (Lxydt6 & M6a7x6);
assign E6kiy6 = (Kbkiy6 & Sbkiy6);
assign Sbkiy6 = (~(Ackiy6 & Bfo7v6));
assign Ackiy6 = (~(Ickiy6 & Qckiy6));
assign Qckiy6 = (~(Zzihw6 & Yckiy6));
assign Ickiy6 = (Gdkiy6 & Odkiy6);
assign Odkiy6 = (~(Wdkiy6 & Ef47x6));
assign Wdkiy6 = (Hbo7v6 & Tnzdt6);
assign Gdkiy6 = (~(R3h7z6[0] & Q4kiy6));
assign Q4kiy6 = (~(Iqmov6 & N3a7x6));
assign Kbkiy6 = (~(Eyknv6 & Rgo7v6));
assign Eyknv6 = (Eekiy6 & Dioov6);
assign O5kiy6 = (Mekiy6 & Uekiy6);
assign Uekiy6 = (Dhyxx6 & Cfkiy6);
assign Cfkiy6 = (~(Clhhw6 & Kfkiy6));
assign Kfkiy6 = (Sfkiy6 | Agkiy6);
assign Agkiy6 = (Qgkiy6 ? Igkiy6 : Noa7x6);
assign Qgkiy6 = (Ygkiy6 & Bfo7v6);
assign Ygkiy6 = (~(W4a7x6 & Tnzdt6));
assign W4a7x6 = (Ghkiy6 & Hjihw6);
assign Igkiy6 = (Ohkiy6 & Zzihw6);
assign Ohkiy6 = (Whkiy6 & M6a7x6);
assign Whkiy6 = (~(Q9xdt6 & Eikiy6));
assign Noa7x6 = (~(Hsa7x6 | Mikiy6));
assign Sfkiy6 = (~(Uikiy6 & Cjkiy6));
assign Cjkiy6 = (~(Kjkiy6 & E9nov6));
assign E9nov6 = (~(F6a7x6 & Sjkiy6));
assign Sjkiy6 = (~(Mikiy6 & Eikiy6));
assign Kjkiy6 = (~(Akkiy6 & Ikkiy6));
assign Ikkiy6 = (~(Qkkiy6 & Ykkiy6));
assign Ykkiy6 = (~(M6a7x6 & Glkiy6));
assign Qkkiy6 = (Aga7z6 & Hjihw6);
assign Akkiy6 = (~(Olkiy6 & M6a7x6));
assign Olkiy6 = (~(Vovxx6 & Pvhhw6));
assign Pvhhw6 = (!Emhhw6);
assign Uikiy6 = (~(Wlkiy6 & Iga7z6));
assign Wlkiy6 = (!F6a7x6);
assign Dhyxx6 = (~(U6hiy6 & Fulnv6));
assign Mekiy6 = (~(Emkiy6 | Ry97x6));
assign Ry97x6 = (~(Mmkiy6 & Umkiy6));
assign Umkiy6 = (~(Cnkiy6 & Ot97x6));
assign Emkiy6 = (Tnzdt6 ? Lyknv6 : Knkiy6);
assign Lyknv6 = (!Snkiy6);
assign Knkiy6 = (Px97x6 & Dwb7z6[5]);
assign Gtjiy6 = (~(Qsinv6 & Aokiy6));
assign Aokiy6 = (~(Iokiy6 & Qokiy6));
assign Qokiy6 = (Yokiy6 & T4jnv6);
assign Yokiy6 = (Tulnv6 & Xxknv6);
assign Iokiy6 = (~(Gpkiy6 | Lna7x6));
assign Lna7x6 = (Fulnv6 & Dioov6);
assign Gpkiy6 = (~(Qxknv6 & X1a7x6));
assign Qsinv6 = (!Aeonv6);
assign Ihaov6 = (!Jbd8x6);
assign Jbd8x6 = (Vuyiw6 & Opkiy6);
assign Vuyiw6 = (~(Wpkiy6 | Eqkiy6));
assign Eqkiy6 = (Xhlhw6 ? Uqkiy6 : Mqkiy6);
assign Xhlhw6 = (Crkiy6 & Krkiy6);
assign Krkiy6 = (~(Dte7z6[3] | Dte7z6[4]));
assign Crkiy6 = (Xu27x6 & J1gov6);
assign Xu27x6 = (Gsz6x6 & Sao6x6);
assign Sao6x6 = (!Dte7z6[15]);
assign Gsz6x6 = (~(Dte7z6[16] | Dte7z6[17]));
assign Mqkiy6 = (~(Srkiy6 & Askiy6));
assign Askiy6 = (~(Iskiy6 & Qskiy6));
assign Qskiy6 = (Yskiy6 & Aetiw6);
assign Iskiy6 = (~(Cu27x6 | Ixfov6));
assign Cu27x6 = (!Gtkiy6);
assign Srkiy6 = (Otkiy6 & Jm8iw6);
assign Otkiy6 = (~(Wtkiy6 & Eukiy6));
assign Eukiy6 = (Mukiy6 & Uukiy6);
assign Uukiy6 = (~(Cvkiy6 & Xariw6));
assign Xariw6 = (Kvkiy6 & Notiw6);
assign Kvkiy6 = (R4aov6 & Qg2nv6);
assign Cvkiy6 = (Svkiy6 & Oo07x6);
assign Svkiy6 = (!Opkiy6);
assign Opkiy6 = (~(Awkiy6 | Iwkiy6));
assign Iwkiy6 = (!B437x6);
assign Mukiy6 = (~(Qwkiy6 | A827x6));
assign Wtkiy6 = (Ywkiy6 & Gxkiy6);
assign Gxkiy6 = (~(Oxkiy6 & M5aov6));
assign Oxkiy6 = (Bdf7z6[1] & Qg2nv6);
assign Ywkiy6 = (~(Gtkiy6 & Yskiy6));
assign Yskiy6 = (!Uh2ov6);
assign Gtkiy6 = (Vo07x6 & Zgtiw6);
assign Zgtiw6 = (~(Zrz6x6 & Wxkiy6));
assign Zrz6x6 = (Dte7z6[13] & Nzz6x6);
assign Wpkiy6 = (~(Ubhdt6 & Pxfov6));
assign Fao7v6 = (Pkkiw6 ? P2xnv6 : Eykiy6);
assign Eykiy6 = (!Vbh7v6);
assign Y9o7v6 = (Pkkiw6 ? R9ynv6 : Mykiy6);
assign Pkkiw6 = (!Tqoov6);
assign Tqoov6 = (~(P6d7z6[0] & Cg1ov6));
assign Mykiy6 = (!Obh7v6);
assign R9o7v6 = (Klkiw6 ? Geynv6 : Uykiy6);
assign Geynv6 = (~(Czkiy6 & Kzkiy6));
assign Kzkiy6 = (~(G7piw6 & HRDATAS[14]));
assign Czkiy6 = (Szkiy6 & A0liy6);
assign A0liy6 = (~(K9piw6 & E4f7x6));
assign E4f7x6 = (~(I0liy6 & Q0liy6));
assign Q0liy6 = (~(Ysnhy6 & Cba7z6));
assign Cba7z6 = (~(Y0liy6 & G1liy6));
assign G1liy6 = (~(HRDATAD[14] & Qln7z6[0]));
assign Y0liy6 = (~(HRDATAS[14] & Qln7z6[1]));
assign I0liy6 = (~(Tim7z6[14] & Uunhy6));
assign Szkiy6 = (~(HRDATAI[14] & Xzjyx6));
assign Xzjyx6 = (~(O1liy6 & W1liy6));
assign W1liy6 = (~(R9piw6 & E2liy6));
assign Uykiy6 = (!Bfh7v6);
assign K9o7v6 = (Klkiw6 ? Zexnv6 : M2liy6);
assign Zexnv6 = (~(U2liy6 & C3liy6));
assign C3liy6 = (~(G7piw6 & HRDATAS[30]));
assign U2liy6 = (K3liy6 & S3liy6);
assign S3liy6 = (~(K9piw6 & Agdiy6));
assign Agdiy6 = (~(A4liy6 & I4liy6));
assign I4liy6 = (~(Um8iy6 & M6a7z6));
assign M6a7z6 = (~(Q4liy6 & Y4liy6));
assign Y4liy6 = (~(HRDATAD[30] & Qln7z6[0]));
assign Q4liy6 = (~(HRDATAS[30] & Qln7z6[1]));
assign A4liy6 = (~(Tim7z6[30] & Yo8iy6));
assign K3liy6 = (~(HRDATAI[30] & X3lyx6));
assign M2liy6 = (!Ueh7v6);
assign D9o7v6 = (Klkiw6 ? N6znv6 : G5liy6);
assign N6znv6 = (~(O5liy6 & W5liy6));
assign W5liy6 = (~(G7piw6 & HRDATAS[16]));
assign O5liy6 = (E6liy6 & M6liy6);
assign M6liy6 = (~(K9piw6 & N4g7x6));
assign N4g7x6 = (~(U6liy6 & C7liy6));
assign C7liy6 = (~(Maa7z6 & Aszhy6));
assign Aszhy6 = (~(K7liy6 & Wdmhy6));
assign K7liy6 = (~(Eemhy6 & S7liy6));
assign S7liy6 = (~(A8liy6 & Q8ixx6));
assign A8liy6 = (~(Ven7z6[0] & I8liy6));
assign Maa7z6 = (~(Q8liy6 & Y8liy6));
assign Y8liy6 = (~(HRDATAD[16] & Qln7z6[0]));
assign Q8liy6 = (~(HRDATAS[16] & Qln7z6[1]));
assign U6liy6 = (~(Tim7z6[16] & Yszhy6));
assign Yszhy6 = (~(G9liy6 & O9liy6));
assign O9liy6 = (Yxixx6 | Kfmhy6);
assign Yxixx6 = (~(Ven7z6[2] & Q8ixx6));
assign G9liy6 = (~(Uunhy6 & Q8ixx6));
assign Q8ixx6 = (!Ven7z6[1]);
assign E6liy6 = (~(HRDATAI[16] & X3lyx6));
assign X3lyx6 = (~(O1liy6 & W9liy6));
assign W9liy6 = (Ealiy6 | Fapiw6);
assign G5liy6 = (!Neh7v6);
assign W8o7v6 = (Klkiw6 ? R9ynv6 : Maliy6);
assign R9ynv6 = (~(Ualiy6 & Cbliy6));
assign Cbliy6 = (Kbliy6 & Bmkyx6);
assign Bmkyx6 = (E2liy6 | Ealiy6);
assign E2liy6 = (~(Hrb7z6[0] & Ryadt6));
assign Kbliy6 = (~(K9piw6 & R7f7x6));
assign R7f7x6 = (~(Sbliy6 & Acliy6));
assign Acliy6 = (~(Uaa7z6 & Ysnhy6));
assign Ysnhy6 = (~(Icliy6 & Wdmhy6));
assign Icliy6 = (~(Ven7z6[0] & Eemhy6));
assign Uaa7z6 = (~(Qcliy6 & Ycliy6));
assign Ycliy6 = (~(HRDATAD[15] & Qln7z6[0]));
assign Qcliy6 = (~(HRDATAS[15] & Qln7z6[1]));
assign Sbliy6 = (~(Tim7z6[15] & Uunhy6));
assign Uunhy6 = (~(Kfmhy6 | Ven7z6[0]));
assign Ualiy6 = (Gdliy6 & Odliy6);
assign Odliy6 = (~(HRDATAI[15] & D9piw6));
assign Gdliy6 = (~(G7piw6 & HRDATAS[15]));
assign Maliy6 = (!Hbh7v6);
assign P8o7v6 = (Klkiw6 ? P2xnv6 : Wdliy6);
assign Klkiw6 = (!As9ov6);
assign As9ov6 = (~(P6d7z6[1] & Cg1ov6));
assign Cg1ov6 = (H11ov6 & Wzcdt6);
assign P2xnv6 = (~(Eeliy6 & Meliy6));
assign Meliy6 = (Ueliy6 & Pnlyx6);
assign Pnlyx6 = (~(Fapiw6 & R9piw6));
assign Fapiw6 = (Hrb7z6[1] & Ryadt6);
assign Ueliy6 = (~(HRDATAI[31] & D9piw6));
assign D9piw6 = (~(O1liy6 & Ealiy6));
assign O1liy6 = (Cfliy6 & Kfliy6);
assign Eeliy6 = (Sfliy6 & Agliy6);
assign Agliy6 = (~(K9piw6 & Kbwnv6));
assign Kbwnv6 = (~(Igliy6 & Qgliy6));
assign Qgliy6 = (~(Vbo7v6 & Um8iy6));
assign Um8iy6 = (~(Ygliy6 & Wdmhy6));
assign Wdmhy6 = (~(Kfmhy6 & Ghliy6));
assign Ghliy6 = (~(Qo8iy6 & A9gxx6));
assign Ygliy6 = (~(Jkqnv6 & Eemhy6));
assign Vbo7v6 = (~(Ohliy6 & Whliy6));
assign Whliy6 = (~(HRDATAD[31] & Qln7z6[0]));
assign Ohliy6 = (~(HRDATAS[31] & Qln7z6[1]));
assign Igliy6 = (~(Tim7z6[31] & Yo8iy6));
assign Yo8iy6 = (~(Kfmhy6 | Jkqnv6));
assign Jkqnv6 = (Eiliy6 & Osixx6);
assign Osixx6 = (!Ven7z6[0]);
assign Kfmhy6 = (!Eemhy6);
assign Eemhy6 = (Ozixx6 & Benyx6);
assign Sfliy6 = (~(G7piw6 & HRDATAS[31]));
assign Wdliy6 = (!Abh7v6);
assign I8o7v6 = (Q52et6 ? Uah7z6[0] : Dwb7z6[0]);
assign B8o7v6 = (Q52et6 ? Uah7z6[1] : Dwb7z6[1]);
assign U7o7v6 = (Q52et6 ? Uah7z6[2] : Dwb7z6[2]);
assign N7o7v6 = (Q52et6 ? Uah7z6[3] : Dwb7z6[3]);
assign G7o7v6 = (Q52et6 ? Uah7z6[4] : Dwb7z6[4]);
assign Z6o7v6 = (Q52et6 ? Uah7z6[5] : Dwb7z6[5]);
assign S6o7v6 = (Cr97z6 ? BIGEND : Evadt6);
assign L6o7v6 = (!Miliy6);
assign Miliy6 = (Cjliy6 ? Uiliy6 : W1mhy6);
assign Uiliy6 = (~(Kjliy6 & Sjliy6));
assign Sjliy6 = (Akliy6 & Pjb7z6[9]);
assign Akliy6 = (Pjb7z6[10] & Pjb7z6[11]);
assign Kjliy6 = (Ikliy6 & Pjb7z6[6]);
assign Ikliy6 = (Pjb7z6[7] & Pjb7z6[8]);
assign W1mhy6 = (!Ti2nz6[5]);
assign E6o7v6 = (P9get6 ? S3a7z6 : Jqj7z6[0]);
assign S3a7z6 = (Uq97z6 | INTNMI);
assign X5o7v6 = (P9get6 ? Tib7z6[63] : Jqj7z6[72]);
assign Q5o7v6 = (P9get6 ? Tib7z6[62] : Jqj7z6[71]);
assign J5o7v6 = (P9get6 ? Tib7z6[61] : Jqj7z6[70]);
assign C5o7v6 = (P9get6 ? Tib7z6[60] : Jqj7z6[69]);
assign V4o7v6 = (P9get6 ? Tib7z6[59] : Jqj7z6[68]);
assign O4o7v6 = (P9get6 ? Tib7z6[58] : Jqj7z6[67]);
assign H4o7v6 = (P9get6 ? Tib7z6[57] : Jqj7z6[66]);
assign A4o7v6 = (P9get6 ? Tib7z6[56] : Jqj7z6[65]);
assign T3o7v6 = (P9get6 ? Tib7z6[55] : Jqj7z6[64]);
assign M3o7v6 = (P9get6 ? Tib7z6[54] : Jqj7z6[63]);
assign F3o7v6 = (P9get6 ? Tib7z6[53] : Jqj7z6[62]);
assign Y2o7v6 = (P9get6 ? Tib7z6[52] : Jqj7z6[61]);
assign R2o7v6 = (P9get6 ? Tib7z6[51] : Jqj7z6[60]);
assign K2o7v6 = (P9get6 ? Tib7z6[50] : Jqj7z6[59]);
assign D2o7v6 = (P9get6 ? Tib7z6[49] : Jqj7z6[58]);
assign W1o7v6 = (P9get6 ? Tib7z6[48] : Jqj7z6[57]);
assign P1o7v6 = (P9get6 ? Tib7z6[47] : Jqj7z6[56]);
assign I1o7v6 = (P9get6 ? Tib7z6[46] : Jqj7z6[55]);
assign B1o7v6 = (P9get6 ? Tib7z6[45] : Jqj7z6[54]);
assign U0o7v6 = (P9get6 ? Tib7z6[44] : Jqj7z6[53]);
assign N0o7v6 = (P9get6 ? Tib7z6[43] : Jqj7z6[52]);
assign G0o7v6 = (P9get6 ? Tib7z6[42] : Jqj7z6[51]);
assign Zzn7v6 = (P9get6 ? Tib7z6[41] : Jqj7z6[50]);
assign Szn7v6 = (P9get6 ? Tib7z6[40] : Jqj7z6[49]);
assign Lzn7v6 = (P9get6 ? Tib7z6[39] : Jqj7z6[48]);
assign Ezn7v6 = (P9get6 ? Tib7z6[38] : Jqj7z6[47]);
assign Xyn7v6 = (P9get6 ? Tib7z6[37] : Jqj7z6[46]);
assign Qyn7v6 = (P9get6 ? Tib7z6[36] : Jqj7z6[45]);
assign Jyn7v6 = (P9get6 ? Tib7z6[35] : Jqj7z6[44]);
assign Cyn7v6 = (P9get6 ? Tib7z6[34] : Jqj7z6[43]);
assign Vxn7v6 = (P9get6 ? Tib7z6[33] : Jqj7z6[42]);
assign Oxn7v6 = (P9get6 ? Tib7z6[32] : Jqj7z6[41]);
assign Hxn7v6 = (P9get6 ? Tib7z6[31] : Jqj7z6[40]);
assign Axn7v6 = (P9get6 ? Tib7z6[30] : Jqj7z6[39]);
assign Twn7v6 = (P9get6 ? Tib7z6[29] : Jqj7z6[38]);
assign Mwn7v6 = (P9get6 ? Tib7z6[28] : Jqj7z6[37]);
assign Fwn7v6 = (P9get6 ? Tib7z6[27] : Jqj7z6[36]);
assign Yvn7v6 = (P9get6 ? Tib7z6[26] : Jqj7z6[35]);
assign Rvn7v6 = (P9get6 ? Tib7z6[25] : Jqj7z6[34]);
assign Kvn7v6 = (P9get6 ? Tib7z6[24] : Jqj7z6[33]);
assign Dvn7v6 = (P9get6 ? Tib7z6[23] : Jqj7z6[32]);
assign Wun7v6 = (P9get6 ? Tib7z6[22] : Jqj7z6[31]);
assign Pun7v6 = (P9get6 ? Tib7z6[21] : Jqj7z6[30]);
assign Iun7v6 = (P9get6 ? Tib7z6[20] : Jqj7z6[29]);
assign Bun7v6 = (P9get6 ? Tib7z6[19] : Jqj7z6[28]);
assign Utn7v6 = (P9get6 ? Tib7z6[18] : Jqj7z6[27]);
assign Ntn7v6 = (P9get6 ? Tib7z6[17] : Jqj7z6[26]);
assign Gtn7v6 = (P9get6 ? Tib7z6[16] : Jqj7z6[25]);
assign Zsn7v6 = (P9get6 ? Tib7z6[15] : Jqj7z6[24]);
assign Ssn7v6 = (P9get6 ? Tib7z6[14] : Jqj7z6[23]);
assign Lsn7v6 = (P9get6 ? Tib7z6[13] : Jqj7z6[22]);
assign Esn7v6 = (P9get6 ? Tib7z6[12] : Jqj7z6[21]);
assign Xrn7v6 = (P9get6 ? Tib7z6[11] : Jqj7z6[20]);
assign Qrn7v6 = (P9get6 ? Tib7z6[10] : Jqj7z6[19]);
assign Jrn7v6 = (P9get6 ? Tib7z6[9] : Jqj7z6[18]);
assign Crn7v6 = (P9get6 ? Tib7z6[8] : Jqj7z6[17]);
assign Vqn7v6 = (P9get6 ? Tib7z6[7] : Jqj7z6[16]);
assign Oqn7v6 = (P9get6 ? Tib7z6[6] : Jqj7z6[15]);
assign Hqn7v6 = (P9get6 ? Tib7z6[5] : Jqj7z6[14]);
assign Aqn7v6 = (P9get6 ? Tib7z6[4] : Jqj7z6[13]);
assign Tpn7v6 = (P9get6 ? Tib7z6[3] : Jqj7z6[12]);
assign Mpn7v6 = (P9get6 ? Tib7z6[2] : Jqj7z6[11]);
assign Fpn7v6 = (P9get6 ? Tib7z6[1] : Jqj7z6[10]);
assign Yon7v6 = (P9get6 ? Tib7z6[0] : Jqj7z6[9]);
assign Ron7v6 = (P9get6 ? Qmj7z6[1] : Jqj7z6[1]);
assign Qmj7z6[1] = (!Mapiw6);
assign Mapiw6 = (Pmh7v6 & Qkliy6);
assign Qkliy6 = (Xsinv6 | F8m7x6);
assign F8m7x6 = (O9m7x6 & U5m7x6);
assign U5m7x6 = (!Ieadt6);
assign O9m7x6 = (Ykliy6 & Glliy6);
assign Glliy6 = (S8b7x6 | Sjcet6);
assign Kon7v6 = (Q0hhw6 ? Rphhw6 : Nzg7z6[0]);
assign Rphhw6 = (Olliy6 ^ Wlliy6);
assign Don7v6 = (Q0hhw6 ? Cehhw6 : Nzg7z6[1]);
assign Cehhw6 = (Emliy6 ^ Mmliy6);
assign Wnn7v6 = (Q0hhw6 ? Rbhhw6 : Nzg7z6[2]);
assign Rbhhw6 = (Umliy6 ^ Cnliy6);
assign Pnn7v6 = (Q0hhw6 ? A6hhw6 : Nzg7z6[3]);
assign A6hhw6 = (~(Knliy6 & Snliy6));
assign Snliy6 = (Aoliy6 & Ioliy6);
assign Ioliy6 = (Qoliy6 & Yoliy6);
assign Yoliy6 = (Gpliy6 | Opliy6);
assign Qoliy6 = (Wpliy6 & Eqliy6);
assign Eqliy6 = (Mqliy6 | Uqliy6);
assign Wpliy6 = (Crliy6 | Krliy6);
assign Aoliy6 = (Srliy6 & Asliy6);
assign Asliy6 = (Isliy6 | Qsliy6);
assign Srliy6 = (Ysliy6 | Gtliy6);
assign Knliy6 = (Otliy6 & Wtliy6);
assign Wtliy6 = (Euliy6 & Muliy6);
assign Muliy6 = (Uuliy6 | Cvliy6);
assign Euliy6 = (Kvliy6 | Svliy6);
assign Otliy6 = (Awliy6 & Iwliy6);
assign Iwliy6 = (Qwliy6 | Ywliy6);
assign Awliy6 = (~(Cnliy6 & Umliy6));
assign Umliy6 = (Ywliy6 ^ Qwliy6);
assign Qwliy6 = (Gxliy6 | Oxliy6);
assign Ywliy6 = (~(Svliy6 ^ Kvliy6));
assign Kvliy6 = (Wxliy6 | Eyliy6);
assign Svliy6 = (~(Cvliy6 ^ Uuliy6));
assign Uuliy6 = (Myliy6 | Uyliy6);
assign Cvliy6 = (~(Gtliy6 ^ Ysliy6));
assign Ysliy6 = (Czliy6 | Kzliy6);
assign Gtliy6 = (~(Qsliy6 ^ Isliy6));
assign Isliy6 = (Szliy6 | A0miy6);
assign Qsliy6 = (~(Opliy6 ^ Gpliy6));
assign Gpliy6 = (I0miy6 | Q0miy6);
assign Opliy6 = (~(Krliy6 ^ Crliy6));
assign Crliy6 = (Y0miy6 | G1miy6);
assign Krliy6 = (~(Uqliy6 ^ Mqliy6));
assign Mqliy6 = (O1miy6 | W1miy6);
assign Uqliy6 = (E2miy6 & M2miy6);
assign M2miy6 = (U2miy6 & C3miy6);
assign C3miy6 = (~(K3miy6 & S3miy6));
assign K3miy6 = (A4miy6 & I4miy6);
assign U2miy6 = (~(Q4miy6 & Y4miy6));
assign E2miy6 = (G5miy6 & O5miy6);
assign O5miy6 = (~(W5miy6 & E6miy6));
assign G5miy6 = (M6miy6 | U6miy6);
assign Cnliy6 = (Mmliy6 & Emliy6);
assign Emliy6 = (Oxliy6 ^ Gxliy6);
assign Gxliy6 = (C7miy6 | K7miy6);
assign Oxliy6 = (~(Eyliy6 ^ Wxliy6));
assign Wxliy6 = (~(S7miy6 & A8miy6));
assign Eyliy6 = (~(Uyliy6 ^ Myliy6));
assign Myliy6 = (I8miy6 | Q8miy6);
assign Uyliy6 = (~(Kzliy6 ^ Czliy6));
assign Czliy6 = (Y8miy6 | G9miy6);
assign Kzliy6 = (~(A0miy6 ^ Szliy6));
assign Szliy6 = (O9miy6 | W9miy6);
assign A0miy6 = (~(Q0miy6 ^ I0miy6));
assign I0miy6 = (~(Eamiy6 & Mamiy6));
assign Q0miy6 = (~(G1miy6 ^ Y0miy6));
assign Y0miy6 = (Uamiy6 | Cbmiy6);
assign G1miy6 = (~(W1miy6 ^ O1miy6));
assign O1miy6 = (Kbmiy6 | Sbmiy6);
assign W1miy6 = (~(U6miy6 ^ M6miy6));
assign M6miy6 = (Acmiy6 | Icmiy6);
assign U6miy6 = (~(Y4miy6 ^ Q4miy6));
assign Q4miy6 = (Qcmiy6 & Ycmiy6);
assign Y4miy6 = (E6miy6 ^ W5miy6);
assign W5miy6 = (~(Gdmiy6 | Odmiy6));
assign E6miy6 = (Wdmiy6 ^ Eemiy6);
assign Eemiy6 = (!A4miy6);
assign A4miy6 = (Memiy6 | Uemiy6);
assign Wdmiy6 = (~(S3miy6 & I4miy6));
assign Mmliy6 = (~(Olliy6 | Wlliy6));
assign Wlliy6 = (Cfmiy6 & Kfmiy6);
assign Kfmiy6 = (~(Sfmiy6 & Pxfhw6));
assign Pxfhw6 = (!L1ohw6);
assign L1ohw6 = (~(Agmiy6 | Igmiy6));
assign Cfmiy6 = (~(Qgmiy6 & R6xxx6));
assign Olliy6 = (~(C7miy6 ^ K7miy6));
assign K7miy6 = (Ygmiy6 & Ghmiy6);
assign Ghmiy6 = (~(Qgmiy6 & Vgwxx6));
assign Ygmiy6 = (Ohmiy6 & Whmiy6);
assign Whmiy6 = (~(Eimiy6 & Mimiy6));
assign Eimiy6 = (V1c7z6[14] & Pxmov6);
assign Ohmiy6 = (~(Sfmiy6 & Dyfhw6));
assign Dyfhw6 = (~(Uimiy6 & Cjmiy6));
assign Cjmiy6 = (Kjmiy6 | Zec7z6[11]);
assign Uimiy6 = (~(Zofhw6 & Zec7z6[30]));
assign C7miy6 = (~(A8miy6 ^ S7miy6));
assign S7miy6 = (Mimiy6 & V1c7z6[13]);
assign Mimiy6 = (Sjmiy6 & Akmiy6);
assign Sjmiy6 = (Q0hhw6 & Ikmiy6);
assign A8miy6 = (I8miy6 ^ Q8miy6);
assign Q8miy6 = (Qkmiy6 & Ykmiy6);
assign Ykmiy6 = (~(Lhwxx6 & Qgmiy6));
assign Qkmiy6 = (Glmiy6 & Olmiy6);
assign Olmiy6 = (~(Wlmiy6 & Q0hhw6));
assign Wlmiy6 = (V1c7z6[12] & Emmiy6);
assign Emmiy6 = (~(Rihhw6 & Mmmiy6));
assign Mmmiy6 = (Kihhw6 | Hir8v6);
assign Glmiy6 = (~(Ummiy6 & Z9nhw6));
assign I8miy6 = (~(Y8miy6 ^ G9miy6));
assign G9miy6 = (Cnmiy6 & Knmiy6);
assign Knmiy6 = (~(Qgmiy6 & L5xxx6));
assign Cnmiy6 = (Snmiy6 & Aomiy6);
assign Aomiy6 = (~(Iomiy6 & Q0hhw6));
assign Iomiy6 = (~(Ceohw6 | Kihhw6));
assign Ceohw6 = (!V1c7z6[11]);
assign Snmiy6 = (~(Ummiy6 & Zec7z6[27]));
assign Y8miy6 = (~(O9miy6 ^ W9miy6));
assign W9miy6 = (Qomiy6 & Yomiy6);
assign Yomiy6 = (~(Qgmiy6 & Pjwxx6));
assign Qomiy6 = (Gpmiy6 & Opmiy6);
assign Opmiy6 = (~(Wpmiy6 & Q0hhw6));
assign Wpmiy6 = (V1c7z6[10] & Eqmiy6);
assign Eqmiy6 = (~(Kihhw6 & Mqmiy6));
assign Mqmiy6 = (~(Uqmiy6 & Pxmov6));
assign Uqmiy6 = (Xumov6 & Xlaov6);
assign Gpmiy6 = (~(Sfmiy6 & Bqfhw6));
assign Bqfhw6 = (Zofhw6 & Zec7z6[26]);
assign O9miy6 = (~(Eamiy6 ^ Mamiy6));
assign Mamiy6 = (~(Crmiy6 & Krmiy6));
assign Krmiy6 = (~(Qgmiy6 & Dxwxx6));
assign Crmiy6 = (Srmiy6 & Asmiy6);
assign Asmiy6 = (~(Ismiy6 & Q0hhw6));
assign Ismiy6 = (V1c7z6[9] & Ikmiy6);
assign Srmiy6 = (~(Ummiy6 & Zec7z6[25]));
assign Eamiy6 = (Uamiy6 ^ Cbmiy6);
assign Cbmiy6 = (Qsmiy6 & Ysmiy6);
assign Ysmiy6 = (~(Gtmiy6 & Qgmiy6));
assign Qsmiy6 = (Otmiy6 & Wtmiy6);
assign Wtmiy6 = (~(Eumiy6 & Q0hhw6));
assign Eumiy6 = (~(E0phw6 | Mumiy6));
assign E0phw6 = (!V1c7z6[8]);
assign Otmiy6 = (~(Ummiy6 & Zec7z6[24]));
assign Ummiy6 = (~(Uumiy6 | Cvmiy6));
assign Uamiy6 = (~(Kbmiy6 ^ Sbmiy6));
assign Sbmiy6 = (Kvmiy6 & Svmiy6);
assign Svmiy6 = (Nwwxx6 | Awmiy6);
assign Kvmiy6 = (Iwmiy6 & Qwmiy6);
assign Qwmiy6 = (~(Ywmiy6 & Q0hhw6));
assign Ywmiy6 = (V1c7z6[7] & Xlaov6);
assign Iwmiy6 = (~(Sfmiy6 & Zvfhw6));
assign Zvfhw6 = (~(Gxmiy6 & Oxmiy6));
assign Oxmiy6 = (~(Zofhw6 & Oenhw6));
assign Gxmiy6 = (Xeinv6 | Bylhw6);
assign Kbmiy6 = (~(Acmiy6 ^ Icmiy6));
assign Icmiy6 = (Wxmiy6 & Eymiy6);
assign Eymiy6 = (Fwwxx6 | Awmiy6);
assign Wxmiy6 = (Mymiy6 & Uymiy6);
assign Uymiy6 = (~(Czmiy6 & Q0hhw6));
assign Czmiy6 = (V1c7z6[6] & Kzmiy6);
assign Kzmiy6 = (~(Dqr8v6 & Szmiy6));
assign Szmiy6 = (~(Akmiy6 & Pxmov6));
assign Akmiy6 = (Xumov6 & Kpaov6);
assign Mymiy6 = (Uumiy6 | Qufhw6);
assign Qufhw6 = (A0niy6 & I0niy6);
assign I0niy6 = (~(Zofhw6 & Uqd7z6[22]));
assign A0niy6 = (Fcinv6 | Bylhw6);
assign Acmiy6 = (~(Qcmiy6 ^ Ycmiy6));
assign Ycmiy6 = (~(Q0niy6 & Y0niy6));
assign Y0niy6 = (~(Qgmiy6 & G1niy6));
assign Q0niy6 = (O1niy6 & W1niy6);
assign W1niy6 = (~(E2niy6 & Q0hhw6));
assign E2niy6 = (~(S7phw6 | M2niy6));
assign S7phw6 = (!V1c7z6[5]);
assign O1niy6 = (~(Sfmiy6 & Svfhw6));
assign Svfhw6 = (~(U2niy6 & C3niy6));
assign C3niy6 = (~(Uqd7z6[21] & Zofhw6));
assign U2niy6 = (Zpehw6 | Bylhw6);
assign Qcmiy6 = (Gdmiy6 ^ Odmiy6);
assign Odmiy6 = (K3niy6 & S3niy6);
assign S3niy6 = (~(Sfmiy6 & Lcqiw6));
assign Lcqiw6 = (~(A4niy6 & I4niy6));
assign I4niy6 = (~(Uqd7z6[20] & Zofhw6));
assign A4niy6 = (Qtnov6 | Bylhw6);
assign K3niy6 = (Q4niy6 & Y4niy6);
assign Y4niy6 = (~(G5niy6 & Q0hhw6));
assign G5niy6 = (V1c7z6[4] & O5niy6);
assign O5niy6 = (~(M2niy6 & W5niy6));
assign W5niy6 = (~(Pxmov6 & Kpaov6));
assign M2niy6 = (Dqr8v6 & E6niy6);
assign E6niy6 = (~(Xumov6 & Kpaov6));
assign Q4niy6 = (~(Pzwxx6 & Qgmiy6));
assign Gdmiy6 = (S3miy6 ^ M6niy6);
assign M6niy6 = (!I4miy6);
assign I4miy6 = (~(U6niy6 & C7niy6));
assign C7niy6 = (~(Sfmiy6 & Vtfhw6));
assign Vtfhw6 = (~(K7niy6 & S7niy6));
assign S7niy6 = (~(Zofhw6 & Uqd7z6[19]));
assign K7niy6 = (U2ohw6 | Bylhw6);
assign U6niy6 = (A8niy6 & I8niy6);
assign I8niy6 = (~(Q8niy6 & Q0hhw6));
assign Q8niy6 = (V1c7z6[3] & Y8niy6);
assign A8niy6 = (Vkwxx6 | Awmiy6);
assign S3miy6 = (~(Memiy6 | G9niy6));
assign G9niy6 = (O9niy6 & W9niy6);
assign Memiy6 = (~(W9niy6 | O9niy6));
assign O9niy6 = (Eaniy6 & Maniy6);
assign Maniy6 = (Uumiy6 | Msfhw6);
assign Msfhw6 = (Uaniy6 & Cbniy6);
assign Cbniy6 = (~(Zofhw6 & Uqd7z6[18]));
assign Uaniy6 = (T5ohw6 | Bylhw6);
assign Uumiy6 = (!Sfmiy6);
assign Eaniy6 = (Kbniy6 & Sbniy6);
assign Sbniy6 = (~(Acniy6 & Icniy6));
assign Acniy6 = (V1c7z6[2] & Qcniy6);
assign Qcniy6 = (~(Hir8v6 & Ycniy6));
assign Kbniy6 = (N4wxx6 | Awmiy6);
assign Awmiy6 = (!Qgmiy6);
assign W9niy6 = (Uemiy6 | Gdniy6);
assign Gdniy6 = (Odniy6 & Wdniy6);
assign Uemiy6 = (~(Odniy6 | Wdniy6));
assign Wdniy6 = (Eeniy6 & Meniy6);
assign Meniy6 = (~(Sfmiy6 & Mhpiw6));
assign Mhpiw6 = (~(Ueniy6 & Cfniy6));
assign Cfniy6 = (~(Zofhw6 & Ovbdt6));
assign Ueniy6 = (Baohw6 | Bylhw6);
assign Eeniy6 = (Kfniy6 & Sfniy6);
assign Sfniy6 = (~(Agniy6 & Q0hhw6));
assign Agniy6 = (V1c7z6[0] & Igniy6);
assign Kfniy6 = (~(Qgniy6 & Qgmiy6));
assign Odniy6 = (Ygniy6 & Ghniy6);
assign Ghniy6 = (~(Ohniy6 & Qgmiy6));
assign Ygniy6 = (Whniy6 & Einiy6);
assign Einiy6 = (~(Icniy6 & V1c7z6[1]));
assign Icniy6 = (Q0hhw6 & Miniy6);
assign Miniy6 = (~(Xkr8v6 & Ycniy6));
assign Whniy6 = (~(Sfmiy6 & Otfhw6));
assign Otfhw6 = (~(Uiniy6 & Cjniy6));
assign Cjniy6 = (~(Zofhw6 & Uqd7z6[17]));
assign Uiniy6 = (S8ohw6 | Bylhw6);
assign Sfmiy6 = (~(Qgmiy6 | Q0hhw6));
assign Q0hhw6 = (Rmwxx6 & Doihw6);
assign Qgmiy6 = (Hjihw6 & Kjniy6);
assign Kjniy6 = (~(Tdxxx6 & Ajphw6));
assign Inn7v6 = (Zhg7x6 ? Sjniy6 : Oreet6);
assign Sjniy6 = (Akniy6 & Ikniy6);
assign Ikniy6 = (!Qkniy6);
assign Qkniy6 = (Shg7x6 ? Pohov6 : Ykniy6);
assign Shg7x6 = (Eofov6 & F02nv6);
assign Eofov6 = (A12nv6 & Glniy6);
assign Glniy6 = (~(Zhg7x6 & Olniy6));
assign Olniy6 = (!Ebdiw6);
assign Ebdiw6 = (U42nv6 & B52nv6);
assign A12nv6 = (~(Wlniy6 & Emniy6));
assign Emniy6 = (Mmniy6 & Umniy6);
assign Umniy6 = (~(X6eet6 & Cnniy6));
assign Cnniy6 = (Kdadt6 | Ldo7v6);
assign Mmniy6 = (~(Knniy6 | Ffeet6));
assign Wlniy6 = (Snniy6 & Opeet6);
assign Snniy6 = (Cbeet6 & Dgo7v6);
assign Ykniy6 = (~(Vveet6 & Cwadt6));
assign Akniy6 = (F52iw6 ? A0fet6 : U42nv6);
assign F52iw6 = (!Awbet6);
assign Bnn7v6 = (Iownv6 ? Khoet6 : Vm1ov6);
assign Umn7v6 = (Iownv6 ? Wmoet6 : Fk9ov6);
assign Nmn7v6 = (~(Ocd7v6 ^ Lkcov6));
assign Lkcov6 = (~(Wmcov6 & Hafxx6));
assign Hafxx6 = (~(Srcov6 | Ju1yx6));
assign Ju1yx6 = (~(Aoniy6 & E5d7v6));
assign Aoniy6 = (Rr0nz6[1] & Cxrnv6);
assign Cxrnv6 = (!Rr0nz6[0]);
assign Srcov6 = (Qqcov6 | Ercov6);
assign Ercov6 = (!Hw0nz6[2]);
assign Qqcov6 = (!Hw0nz6[1]);
assign Wmcov6 = (Ioniy6 & Uzcov6);
assign Uzcov6 = (Sr5ov6 & Nlcov6);
assign Nlcov6 = (!Fed7v6);
assign Sr5ov6 = (Gs5ov6 & Jysyx6);
assign Jysyx6 = (~(Ioniy6 & Fed7v6));
assign Gs5ov6 = (!Lr5ov6);
assign Lr5ov6 = (At67v6 ? Yoniy6 : Qoniy6);
assign Yoniy6 = (~(Bed8x6 & Pbpyx6));
assign Bed8x6 = (Xid8x6 & V4pyx6);
assign V4pyx6 = (Gpniy6 & Mulhy6);
assign Gpniy6 = (~(Opniy6 | Xfymz6[8]));
assign Qoniy6 = (N4pyx6 & W197z6);
assign N4pyx6 = (Byhyx6 ? Za2yx6 : Ziryx6);
assign Byhyx6 = (!Eee7v6);
assign Za2yx6 = (Hae7v6 ? Eqniy6 : Wpniy6);
assign Eqniy6 = (~(Mqniy6 & P72yx6));
assign P72yx6 = (!N82yx6);
assign N82yx6 = (Uqniy6 & Puhiw6);
assign Puhiw6 = (!J02nz6[4]);
assign Uqniy6 = (!Eqciy6);
assign Eqciy6 = (~(Crniy6 & Krniy6));
assign Krniy6 = (J02nz6[2] & Czlhy6);
assign Czlhy6 = (!J02nz6[8]);
assign Crniy6 = (Hae7v6 & Tppyx6);
assign Tppyx6 = (Srniy6 & J02nz6[5]);
assign Srniy6 = (J02nz6[3] & Xvxyx6);
assign Xvxyx6 = (Asniy6 & Isniy6);
assign Isniy6 = (J02nz6[6] & Thiiw6);
assign Thiiw6 = (Qsniy6 & J02nz6[9]);
assign Qsniy6 = (J02nz6[11] & J02nz6[10]);
assign Asniy6 = (Jke7v6 & J02nz6[7]);
assign Mqniy6 = (~(Bv1nz6[1] & Bv1nz6[0]));
assign Wpniy6 = (Ysniy6 & Gtniy6);
assign Gtniy6 = (~(L92yx6 ^ Ra3yx6));
assign Ra3yx6 = (~(Ja3yx6 ^ Lj1nz6[0]));
assign L92yx6 = (T92yx6 ^ Ja1nz6[0]);
assign Ysniy6 = (Otniy6 & Wtniy6);
assign Wtniy6 = (Ja1nz6[2] ^ Lj1nz6[2]);
assign Otniy6 = (T92yx6 ^ Ja3yx6);
assign Ja3yx6 = (Fah7v6 ^ Lj1nz6[2]);
assign T92yx6 = (Ja1nz6[1] ^ Ja1nz6[2]);
assign Ziryx6 = (!Hce7v6);
assign Ioniy6 = (Jazxx6 & D11yx6);
assign D11yx6 = (~(Euniy6 & Muniy6));
assign Muniy6 = (~(Uuniy6 | Ft0nz6[2]));
assign Uuniy6 = (Ft0nz6[3] | Ft0nz6[4]);
assign Euniy6 = (~(K1dov6 | Ft0nz6[1]));
assign K1dov6 = (!Ft0nz6[0]);
assign Jazxx6 = (!H3dov6);
assign H3dov6 = (~(E15xx6 | L15xx6));
assign L15xx6 = (!Az4xx6);
assign Az4xx6 = (Uu0nz6[2] | Uu0nz6[1]);
assign E15xx6 = (!S15xx6);
assign S15xx6 = (~(Uu0nz6[4] | Uu0nz6[3]));
assign Gmn7v6 = (P9get6 ? Qmj7z6[4] : Jqj7z6[4]);
assign Qmj7z6[4] = (Ykliy6 & Cvniy6);
assign Zln7v6 = (P9get6 ? Zrbet6 : Jqj7z6[6]);
assign Zrbet6 = (~(Kvniy6 & Svniy6));
assign Svniy6 = (~(Hyhov6 & Gr5iw6));
assign Kvniy6 = (Awniy6 & Iwniy6);
assign Iwniy6 = (~(Q7hov6 & Qwniy6));
assign Qwniy6 = (~(Kd2nv6 & Ywniy6));
assign Ywniy6 = (~(Zgadt6 & Gxniy6));
assign Gxniy6 = (~(Zamov6 & Oxniy6));
assign Oxniy6 = (~(Sa2nv6 & Iahov6));
assign Iahov6 = (!Lim7x6);
assign Lim7x6 = (C0i7x6 & Dc3nv6);
assign Dc3nv6 = (F4j7x6 & E7iov6);
assign E7iov6 = (!P2j7z6[4]);
assign F4j7x6 = (Owjov6 & Wfjov6);
assign Wfjov6 = (!P2j7z6[6]);
assign Owjov6 = (!P2j7z6[5]);
assign C0i7x6 = (Wxniy6 & Rc3nv6);
assign Rc3nv6 = (~(Z7iov6 | U1iov6));
assign U1iov6 = (!P2j7z6[2]);
assign Z7iov6 = (!P2j7z6[3]);
assign Wxniy6 = (Bgiov6 & Rgjov6);
assign Rgjov6 = (!P2j7z6[1]);
assign Bgiov6 = (!P2j7z6[0]);
assign Sa2nv6 = (!Ga3nv6);
assign Ga3nv6 = (~(Eyniy6 & Hbo7v6));
assign Eyniy6 = (Ggoov6 & Myniy6);
assign Myniy6 = (~(Xvxxx6 & Uyniy6));
assign Uyniy6 = (~(Czniy6 & Uuinv6));
assign Czniy6 = (O5a7z6 & Dwb7z6[1]);
assign Zamov6 = (Hwr7x6 & X0b7x6);
assign X0b7x6 = (~(Kzniy6 & E1wnv6));
assign E1wnv6 = (!J0b7x6);
assign J0b7x6 = (~(Szniy6 & A0oiy6));
assign A0oiy6 = (~(I0oiy6 | Jai8v6));
assign Jai8v6 = (Q0oiy6 & Qg2nv6);
assign I0oiy6 = (Loddt6 | Pqddt6);
assign Szniy6 = (Y0oiy6 & Drsiw6);
assign Drsiw6 = (G1oiy6 & O1oiy6);
assign O1oiy6 = (W1oiy6 & E2oiy6);
assign E2oiy6 = (~(M2oiy6 & Mrnov6));
assign Mrnov6 = (~(Ketnv6 | Tnzdt6));
assign M2oiy6 = (U2oiy6 & C0wnv6);
assign U2oiy6 = (M0edt6 | Qyddt6);
assign W1oiy6 = (Xfnov6 & C3oiy6);
assign C3oiy6 = (~(M3e7z6[1] & M2jiy6));
assign M2jiy6 = (~(Tnzdt6 | P6u6x6));
assign Xfnov6 = (~(Shfov6 & K3oiy6));
assign K3oiy6 = (~(Henov6 & S3oiy6));
assign Henov6 = (A4oiy6 & I4oiy6);
assign I4oiy6 = (~(Frgov6 & Ipgov6));
assign Ipgov6 = (Ibe7z6[2] | Ibe7z6[1]);
assign Frgov6 = (Q4oiy6 & Y4oiy6);
assign Y4oiy6 = (~(G5oiy6 & O5oiy6));
assign O5oiy6 = (~(Ppb7z6[7] & W5oiy6));
assign G5oiy6 = (E6oiy6 & J92nv6);
assign E6oiy6 = (~(M6oiy6 & U6oiy6));
assign U6oiy6 = (W5oiy6 | Ppb7z6[7]);
assign W5oiy6 = (!Fhc7z6[7]);
assign M6oiy6 = (C7oiy6 & K7oiy6);
assign K7oiy6 = (~(Fhc7z6[6] & S7oiy6));
assign S7oiy6 = (A8oiy6 | I8oiy6);
assign C7oiy6 = (~(A8oiy6 & I8oiy6));
assign A8oiy6 = (Q8oiy6 | Fhc7z6[5]);
assign A4oiy6 = (Y8oiy6 & G9oiy6);
assign G9oiy6 = (Jfnov6 | Nmadt6);
assign Jfnov6 = (O9oiy6 & W9oiy6);
assign W9oiy6 = (~(Ibe7z6[0] & E3c7z6[0]));
assign O9oiy6 = (~(I9e7z6[2] & I9e7z6[0]));
assign Y8oiy6 = (~(Etinv6 & Eaoiy6));
assign Eaoiy6 = (~(Flfov6 & Kkfov6));
assign Kkfov6 = (~(I9e7z6[1] & I9e7z6[0]));
assign Flfov6 = (~(Ibe7z6[3] & E3c7z6[0]));
assign Shfov6 = (~(Gbo6x6 | Z7edt6));
assign G1oiy6 = (Maoiy6 & Uaoiy6);
assign Uaoiy6 = (Tnzdt6 ? Kboiy6 : Cboiy6);
assign Kboiy6 = (~(Z7edt6 & S3oiy6));
assign S3oiy6 = (!Ibe7z6[4]);
assign Cboiy6 = (~(M3e7z6[0] & Bklhw6));
assign Bklhw6 = (~(Sboiy6 & Acoiy6));
assign Acoiy6 = (Fulnv6 & Spdiw6);
assign Sboiy6 = (P6u6x6 & Ltvxx6);
assign Maoiy6 = (M8lov6 & Ixfov6);
assign M8lov6 = (Icoiy6 & Qcoiy6);
assign Qcoiy6 = (Ycoiy6 & Gdoiy6);
assign Gdoiy6 = (Odoiy6 & Wdoiy6);
assign Wdoiy6 = (~(Dwb7z6[2] & Eeoiy6));
assign Eeoiy6 = (~(Meoiy6 & Ueoiy6));
assign Ueoiy6 = (~(Ypinv6 & Cfoiy6));
assign Cfoiy6 = (Htmov6 | Dwb7z6[0]);
assign Meoiy6 = (Buvxx6 & Sna7x6);
assign Buvxx6 = (!Fxaov6);
assign Odoiy6 = (Kfoiy6 & Sfoiy6);
assign Sfoiy6 = (!Eekiy6);
assign Ycoiy6 = (Agoiy6 & Igoiy6);
assign Igoiy6 = (~(Dwb7z6[3] & Ypinv6));
assign Ypinv6 = (!O5a7z6);
assign Agoiy6 = (Qgoiy6 & Ygoiy6);
assign Ygoiy6 = (~(Tka7x6 & Ghoiy6));
assign Ghoiy6 = (~(Ohoiy6 & Msmov6));
assign Msmov6 = (~(Vrinv6 | Aga7z6));
assign Vrinv6 = (!Gr2et6);
assign Ohoiy6 = (Whoiy6 & U1jnv6);
assign Whoiy6 = (~(Htmov6 & N1jnv6));
assign N1jnv6 = (~(Eioiy6 & Mioiy6));
assign Mioiy6 = (Ii9ov6 & Xodiw6);
assign Eioiy6 = (Qodiw6 & T3cdt6);
assign Htmov6 = (~(Cgsiw6 | Wp37x6));
assign Wp37x6 = (S0jnv6 & P2jnv6);
assign P2jnv6 = (~(Uioiy6 & T3cdt6));
assign Uioiy6 = (Kldiw6 & Ii9ov6);
assign Kldiw6 = (~(Hsa7x6 | Qodiw6));
assign Qodiw6 = (Cjoiy6 & Kjoiy6);
assign Kjoiy6 = (~(Sjoiy6 & Akoiy6));
assign Akoiy6 = (!Pgqnv6);
assign Sjoiy6 = (!Yhqnv6);
assign Cjoiy6 = (~(O7adt6 & Ikoiy6));
assign S0jnv6 = (Qkoiy6 & Ykoiy6);
assign Ykoiy6 = (Gloiy6 & Oloiy6);
assign Oloiy6 = (Dsriw6 & Tlyxx6);
assign Dsriw6 = (~(Wloiy6 & Axihw6));
assign Wloiy6 = (~(Hxihw6 | Lofhw6));
assign Gloiy6 = (Emoiy6 & O5jiy6);
assign O5jiy6 = (~(Mmoiy6 & Umoiy6));
assign Mmoiy6 = (Cnoiy6 & X7wxx6);
assign Cnoiy6 = (Knoiy6 | Ozbdt6);
assign Knoiy6 = (Pxfov6 & Snoiy6);
assign Snoiy6 = (~(Hsa7x6 & Xodiw6));
assign Xodiw6 = (!Bi9ov6);
assign Emoiy6 = (~(Aooiy6 & Bi9ov6));
assign Aooiy6 = (~(Ketnv6 | Iooiy6));
assign Qkoiy6 = (~(Qooiy6 | Yooiy6));
assign Yooiy6 = (Zzihw6 ? Gpoiy6 : Kvbov6);
assign Gpoiy6 = (~(Iooiy6 & Opoiy6));
assign Opoiy6 = (~(Wpoiy6 & Eqoiy6));
assign Eqoiy6 = (~(Ketnv6 & Mqoiy6));
assign Iooiy6 = (Uqoiy6 & Croiy6);
assign Croiy6 = (~(Kroiy6 & Sroiy6));
assign Sroiy6 = (Asoiy6 & Isoiy6);
assign Isoiy6 = (Z8c7z6[0] ^ Qsoiy6);
assign Asoiy6 = (Ysoiy6 & Gtoiy6);
assign Gtoiy6 = (Z8c7z6[2] ^ Otoiy6);
assign Ysoiy6 = (~(Wtoiy6 ^ Euoiy6));
assign Kroiy6 = (Xvehw6 & Muoiy6);
assign Muoiy6 = (~(Mqoiy6 ^ Uuoiy6));
assign Uqoiy6 = (~(Cvoiy6 & Kvoiy6));
assign Kvoiy6 = (Svoiy6 & Awoiy6);
assign Awoiy6 = (Mqoiy6 ^ Iwoiy6);
assign Svoiy6 = (Qwoiy6 ^ Ywoiy6);
assign Cvoiy6 = (Gxoiy6 & Oxoiy6);
assign Oxoiy6 = (Wtoiy6 ^ Wxoiy6);
assign Gxoiy6 = (Eyoiy6 ^ Myoiy6);
assign Qooiy6 = (~(Uyoiy6 & G5jiy6));
assign G5jiy6 = (~(Umoiy6 & Czoiy6));
assign Umoiy6 = (Qalhw6 & Kzoiy6);
assign Kzoiy6 = (~(Szoiy6 & A0piy6));
assign A0piy6 = (~(I0piy6 & Q0piy6));
assign Q0piy6 = (Y0piy6 & G1piy6);
assign G1piy6 = (O1piy6 ^ Ywoiy6);
assign Y0piy6 = (W1piy6 ^ Wxoiy6);
assign I0piy6 = (E2piy6 & M2piy6);
assign M2piy6 = (U2piy6 ^ Myoiy6);
assign E2piy6 = (C3piy6 ^ Iwoiy6);
assign Szoiy6 = (~(K3piy6 & S3piy6));
assign S3piy6 = (A4piy6 & I4piy6);
assign I4piy6 = (~(O1piy6 ^ Qsoiy6));
assign O1piy6 = (Q4piy6 & Y4piy6);
assign Y4piy6 = (~(Seihw6 & X7wxx6));
assign Seihw6 = (!P437x6);
assign P437x6 = (G5piy6 & O5piy6);
assign O5piy6 = (W5piy6 & E6piy6);
assign E6piy6 = (M6piy6 & U6piy6);
assign U6piy6 = (C7piy6 | K7piy6);
assign M6piy6 = (S7piy6 | A8piy6);
assign W5piy6 = (I8piy6 & Q8piy6);
assign Q8piy6 = (Hir8v6 | Y8piy6);
assign I8piy6 = (~(O5h7z6[0] & G9piy6));
assign G5piy6 = (O9piy6 & W9piy6);
assign W9piy6 = (Eapiy6 & Mapiy6);
assign Mapiy6 = (~(Qij7z6[0] & Ztaov6));
assign Eapiy6 = (~(Ts97x6 & Ntg7z6[0]));
assign O9piy6 = (Uapiy6 & Cbpiy6);
assign Cbpiy6 = (~(E8h7z6[0] & Kbpiy6));
assign Q4piy6 = (~(Oac7z6[0] & Czoiy6));
assign A4piy6 = (Sbpiy6 & Xvehw6);
assign Xvehw6 = (Acpiy6 & Icpiy6);
assign Icpiy6 = (Qcpiy6 & Ycpiy6);
assign Ycpiy6 = (~(Gdpiy6 | Odpiy6));
assign Qcpiy6 = (Fefhw6 & Wdpiy6);
assign Acpiy6 = (Eepiy6 & Mepiy6);
assign Mepiy6 = (C3riw6 & Cfiiy6);
assign Cfiiy6 = (Ddsiw6 & Aulhw6);
assign Eepiy6 = (Wcsiw6 & V2riw6);
assign Sbpiy6 = (~(W1piy6 ^ Euoiy6));
assign W1piy6 = (Uepiy6 & Cfpiy6);
assign Cfpiy6 = (~(Gfihw6 & X7wxx6));
assign Gfihw6 = (~(Kfpiy6 & Sfpiy6));
assign Sfpiy6 = (Agpiy6 & Igpiy6);
assign Igpiy6 = (Qgpiy6 & Ygpiy6);
assign Ygpiy6 = (~(Ts97x6 & Ntg7z6[3]));
assign Agpiy6 = (Ghpiy6 & Ohpiy6);
assign Ohpiy6 = (Dqr8v6 | Y8piy6);
assign Ghpiy6 = (Whpiy6 | K7piy6);
assign Kfpiy6 = (Eipiy6 & Mipiy6);
assign Mipiy6 = (Uipiy6 & Cjpiy6);
assign Cjpiy6 = (~(Qij7z6[3] & Ztaov6));
assign Uipiy6 = (Kjpiy6 & Sjpiy6);
assign Sjpiy6 = (~(O5h7z6[3] & G9piy6));
assign Kjpiy6 = (S7piy6 | Akpiy6);
assign Eipiy6 = (Uapiy6 & Ikpiy6);
assign Ikpiy6 = (~(E8h7z6[3] & Kbpiy6));
assign Uepiy6 = (~(Czoiy6 & Oac7z6[3]));
assign K3piy6 = (Qkpiy6 & Ykpiy6);
assign Ykpiy6 = (~(U2piy6 ^ Otoiy6));
assign U2piy6 = (Glpiy6 & Olpiy6);
assign Olpiy6 = (~(Qdihw6 & X7wxx6));
assign Qdihw6 = (!L937x6);
assign L937x6 = (Wlpiy6 & Empiy6);
assign Empiy6 = (Mmpiy6 & Umpiy6);
assign Umpiy6 = (Qgpiy6 & Cnpiy6);
assign Cnpiy6 = (Nnr8v6 | Y8piy6);
assign Qgpiy6 = (Ayaov6 & Elphw6);
assign Mmpiy6 = (Knpiy6 & Snpiy6);
assign Snpiy6 = (~(O5h7z6[2] & G9piy6));
assign Knpiy6 = (S7piy6 | Aopiy6);
assign Wlpiy6 = (Iopiy6 & Qopiy6);
assign Qopiy6 = (Yopiy6 & Gppiy6);
assign Gppiy6 = (Oppiy6 | K7piy6);
assign Yopiy6 = (Wppiy6 & Eqpiy6);
assign Eqpiy6 = (~(E8h7z6[2] & Kbpiy6));
assign Wppiy6 = (~(Ts97x6 & Ntg7z6[2]));
assign Iopiy6 = (Uapiy6 & Mqpiy6);
assign Mqpiy6 = (~(Qij7z6[2] & Ztaov6));
assign Uapiy6 = (Uqpiy6 & Crpiy6);
assign Crpiy6 = (Krpiy6 & G3a7x6);
assign G3a7x6 = (~(Eekiy6 & Uvvnv6));
assign Krpiy6 = (Snkiy6 & Qxknv6);
assign Qxknv6 = (~(Kophw6 & Ytlnv6));
assign Kophw6 = (Dwb7z6[4] & Kioov6);
assign Snkiy6 = (~(Srpiy6 & Vqihw6));
assign Srpiy6 = (Dioov6 & Dwb7z6[5]);
assign Uqpiy6 = (Aspiy6 & Ispiy6);
assign Ispiy6 = (~(Qij7z6[4] & Ztaov6));
assign Glpiy6 = (~(Czoiy6 & Oac7z6[2]));
assign Qkpiy6 = (~(C3piy6 ^ Uuoiy6));
assign C3piy6 = (Qspiy6 & Yspiy6);
assign Yspiy6 = (~(Vcihw6 & X7wxx6));
assign X7wxx6 = (~(Gtpiy6 & Otpiy6));
assign Otpiy6 = (Wtpiy6 & Elphw6);
assign Wtpiy6 = (~(R3h7z6[0] & Eupiy6));
assign Eupiy6 = (~(N3a7x6 & U3a7x6));
assign Gtpiy6 = (Mupiy6 & Uupiy6);
assign Uupiy6 = (~(Pi9ov6 & Vxihw6));
assign Mupiy6 = (~(M6a7x6 & Cvpiy6));
assign Cvpiy6 = (~(Kvpiy6 & Svpiy6));
assign Svpiy6 = (~(Zzihw6 & Awpiy6));
assign Awpiy6 = (~(I1d7x6 & Hjihw6));
assign I1d7x6 = (!Yckiy6);
assign Kvpiy6 = (~(Bh2et6 & Iwpiy6));
assign Iwpiy6 = (~(Qwpiy6 & Ywpiy6));
assign Ywpiy6 = (~(S2a7x6 & Ytlnv6));
assign Qwpiy6 = (Gxpiy6 & N3a7x6);
assign Gxpiy6 = (Oxpiy6 | Dwb7z6[3]);
assign M6a7x6 = (!Wbxdt6);
assign Vcihw6 = (!G337x6);
assign G337x6 = (Wxpiy6 & Eypiy6);
assign Eypiy6 = (Mypiy6 & Uypiy6);
assign Uypiy6 = (Czpiy6 & Ayaov6);
assign Ayaov6 = (~(Dophw6 & Vqihw6));
assign Czpiy6 = (Kzpiy6 & Elphw6);
assign Kzpiy6 = (~(Szpiy6 & Qij7z6[1]));
assign Szpiy6 = (Ztaov6 & Tdwxx6);
assign Mypiy6 = (A0qiy6 & I0qiy6);
assign I0qiy6 = (~(O5h7z6[1] & G9piy6));
assign G9piy6 = (~(Q0qiy6 | Y0qiy6));
assign Q0qiy6 = (Whxdt6 & Uebdt6);
assign A0qiy6 = (~(Ts97x6 & Ntg7z6[1]));
assign Ts97x6 = (Yckiy6 & G1qiy6);
assign Wxpiy6 = (O1qiy6 & W1qiy6);
assign W1qiy6 = (E2qiy6 & M2qiy6);
assign M2qiy6 = (Xkr8v6 | Y8piy6);
assign Y8piy6 = (~(U2qiy6 | Dihhw6));
assign U2qiy6 = (C3qiy6 & K3qiy6);
assign K3qiy6 = (S3qiy6 | A4qiy6);
assign E2qiy6 = (I4qiy6 & Q4qiy6);
assign Q4qiy6 = (S7piy6 | C8a7x6);
assign S7piy6 = (~(Y4qiy6 & G5qiy6));
assign G5qiy6 = (Vt97x6 & Uvvnv6);
assign Y4qiy6 = (Y0qiy6 & S2a7x6);
assign I4qiy6 = (O9kiy6 | K7piy6);
assign K7piy6 = (O5qiy6 & W5qiy6);
assign W5qiy6 = (E6qiy6 & M6qiy6);
assign M6qiy6 = (~(U6qiy6 & C3qiy6));
assign C3qiy6 = (Ruxxx6 & Luvnv6);
assign U6qiy6 = (~(S3qiy6 | A4qiy6));
assign A4qiy6 = (F6a7x6 & C7qiy6);
assign C7qiy6 = (~(Vxihw6 & K7qiy6));
assign K7qiy6 = (~(N6xiw6 & Bfo7v6));
assign F6a7x6 = (Glkiy6 | S7qiy6);
assign S7qiy6 = (!Mikiy6);
assign Mikiy6 = (Q9xdt6 & Zzihw6);
assign S3qiy6 = (!D5a7x6);
assign D5a7x6 = (~(Lxydt6 | Emhhw6));
assign Emhhw6 = (Wfxdt6 & Bfo7v6);
assign E6qiy6 = (T4jnv6 & Tulnv6);
assign O5qiy6 = (A8qiy6 & Mmkiy6);
assign Mmkiy6 = (~(I8qiy6 & Yckiy6));
assign I8qiy6 = (!G1qiy6);
assign G1qiy6 = (~(Iga7z6 & Q8qiy6));
assign A8qiy6 = (~(Y8qiy6 & Y0qiy6));
assign Y8qiy6 = (Cnkiy6 & S2a7x6);
assign Cnkiy6 = (!Vt97x6);
assign Vt97x6 = (~(Aga7z6 & Q8qiy6));
assign Q8qiy6 = (~(Hsa7x6 & Wjfhw6));
assign Wjfhw6 = (!Q9xdt6);
assign Hsa7x6 = (!Vxihw6);
assign O1qiy6 = (Aspiy6 & G9qiy6);
assign G9qiy6 = (~(E8h7z6[1] & Kbpiy6));
assign Kbpiy6 = (O9qiy6 & Whxdt6);
assign O9qiy6 = (~(Ijmov6 | Y0qiy6));
assign Y0qiy6 = (W9qiy6 & N3a7x6);
assign N3a7x6 = (Tpvxx6 | Dwb7z6[1]);
assign W9qiy6 = (U3a7x6 & Oxpiy6);
assign U3a7x6 = (!M2kiy6);
assign M2kiy6 = (Ltvxx6 & Vqihw6);
assign Aspiy6 = (Eaqiy6 & Maqiy6);
assign Maqiy6 = (Uaqiy6 & Cbqiy6);
assign Cbqiy6 = (~(Riuxx6 & Luvnv6));
assign Riuxx6 = (~(Zna7x6 | Sna7x6));
assign Uaqiy6 = (Kbqiy6 & X1a7x6);
assign X1a7x6 = (~(Ywaov6 & Dwb7z6[2]));
assign Kbqiy6 = (~(Tiphw6 & Kioov6));
assign Eaqiy6 = (Sbqiy6 & Acqiy6);
assign Acqiy6 = (~(Icqiy6 & Vqihw6));
assign Icqiy6 = (Nvvnv6 & Gvvnv6);
assign Sbqiy6 = (Q1a7x6 & Ix97x6);
assign Ix97x6 = (~(Qcqiy6 & Dioov6));
assign Qcqiy6 = (Fxaov6 & Dwb7z6[5]);
assign Q1a7x6 = (~(Ckphw6 & Fulnv6));
assign Ckphw6 = (Lpwxx6 & Uvvnv6);
assign Qspiy6 = (~(Czoiy6 & Oac7z6[1]));
assign Czoiy6 = (Ycqiy6 & Ixfov6);
assign Ixfov6 = (Gdqiy6 & Jm8iw6);
assign Jm8iw6 = (!Zjb7z6[9]);
assign Gdqiy6 = (~(Pxfov6 & Odqiy6));
assign Odqiy6 = (~(Wdqiy6 & Eeqiy6));
assign Eeqiy6 = (~(Meqiy6 & Ueqiy6));
assign Ueqiy6 = (Cfqiy6 & Kfqiy6);
assign Kfqiy6 = (~(Sfqiy6 & Notiw6));
assign Sfqiy6 = (V9riw6 & Oo07x6);
assign V9riw6 = (Agqiy6 & Igqiy6);
assign Igqiy6 = (Qgqiy6 & Ygqiy6);
assign Ygqiy6 = (Ghqiy6 & Ohqiy6);
assign Ohqiy6 = (~(Uh2ov6 | M6jiy6));
assign Uh2ov6 = (J1gov6 & Wxkiy6);
assign Ghqiy6 = (Whqiy6 & D7u6x6);
assign D7u6x6 = (~(Doadt6 & Eiqiy6));
assign Eiqiy6 = (~(Miqiy6 & Tdxxx6));
assign Tdxxx6 = (Twphw6 & T4jnv6);
assign T4jnv6 = (!Cwlnv6);
assign Miqiy6 = (~(Dur7x6 | Fvr7x6));
assign Fvr7x6 = (Uiqiy6 & Ydziw6);
assign Uiqiy6 = (~(Ketnv6 | Cngdt6));
assign Ketnv6 = (!Pxfov6);
assign Dur7x6 = (~(Tpvxx6 | Bwvnv6));
assign Tpvxx6 = (!Mahiy6);
assign Whqiy6 = (~(Cjqiy6 & Kjqiy6));
assign Kjqiy6 = (Sjqiy6 & Akqiy6);
assign Akqiy6 = (Ovbdt6 ^ Qwoiy6);
assign Sjqiy6 = (Uqd7z6[17] ^ Mqoiy6);
assign Cjqiy6 = (Ikqiy6 & Qkqiy6);
assign Qkqiy6 = (Uqd7z6[18] ^ Eyoiy6);
assign Ikqiy6 = (Uqd7z6[19] ^ Wtoiy6);
assign Qgqiy6 = (Ykqiy6 & Ydziw6);
assign Ykqiy6 = (Pxfov6 & Glqiy6);
assign Glqiy6 = (~(Olqiy6 & Wlqiy6));
assign Wlqiy6 = (Emqiy6 & Mmqiy6);
assign Mmqiy6 = (Zec7z6[0] ^ Qwoiy6);
assign Emqiy6 = (Zec7z6[1] ^ Mqoiy6);
assign Olqiy6 = (Umqiy6 & Cnqiy6);
assign Cnqiy6 = (Zec7z6[2] ^ Eyoiy6);
assign Umqiy6 = (Zec7z6[3] ^ Wtoiy6);
assign Agqiy6 = (Knqiy6 & Snqiy6);
assign Snqiy6 = (Aoqiy6 & Ioqiy6);
assign Ioqiy6 = (Z9nhw6 ^ Qwoiy6);
assign Qwoiy6 = (!Z8c7z6[0]);
assign Aoqiy6 = (Uyoiy6 & Oqviw6);
assign Oqviw6 = (Qoqiy6 & Q1ghw6);
assign Q1ghw6 = (!Q8onv6);
assign Qoqiy6 = (!Mhwiw6);
assign Mhwiw6 = (~(Yoqiy6 & X8onv6));
assign Yoqiy6 = (P8wiw6 & E9onv6);
assign Knqiy6 = (Gpqiy6 & Opqiy6);
assign Opqiy6 = (Zec7z6[30] ^ Eyoiy6);
assign Eyoiy6 = (!Z8c7z6[2]);
assign Gpqiy6 = (Wpqiy6 & Eqqiy6);
assign Eqqiy6 = (Zec7z6[31] ^ Wtoiy6);
assign Wpqiy6 = (M6nhw6 ^ Mqoiy6);
assign Mqoiy6 = (!Z8c7z6[1]);
assign Cfqiy6 = (~(A827x6 | Nvtiw6));
assign Nvtiw6 = (!Ot27x6);
assign Ot27x6 = (~(Mqqiy6 & Bdf7z6[0]));
assign Mqqiy6 = (Muhiy6 & D4aov6);
assign Muhiy6 = (~(Ju27x6 | Bdf7z6[1]));
assign A827x6 = (~(D4aov6 | Y4aov6));
assign Y4aov6 = (!G427x6);
assign G427x6 = (Bdf7z6[1] & Bdf7z6[0]);
assign Meqiy6 = (Uqqiy6 & Crqiy6);
assign Crqiy6 = (Ol8iw6 | Krqiy6);
assign Krqiy6 = (Ydziw6 & Nf4ov6);
assign Nf4ov6 = (!Oztiw6);
assign Oztiw6 = (Wxkiy6 & Xp07x6);
assign Ydziw6 = (!H827x6);
assign H827x6 = (J227x6 | Svziw6);
assign Svziw6 = (Srqiy6 & Dte7z6[15]);
assign Srqiy6 = (~(Zao6x6 | J227x6));
assign Zao6x6 = (!Xp07x6);
assign Xp07x6 = (Dte7z6[14] & Dte7z6[13]);
assign Ol8iw6 = (~(Asqiy6 & Ngxxx6));
assign Asqiy6 = (K4aov6 & Ju27x6);
assign Uqqiy6 = (~(Isqiy6 & Aetiw6));
assign Aetiw6 = (!Ehgdt6);
assign Isqiy6 = (Tdtiw6 | Qwkiy6);
assign Qwkiy6 = (Qsqiy6 & M5aov6);
assign Qsqiy6 = (Bdf7z6[0] & Oo07x6);
assign Oo07x6 = (!Vo07x6);
assign Vo07x6 = (~(Ysqiy6 | Djgdt6));
assign Ysqiy6 = (Bqziw6 & Wxkiy6);
assign Wxkiy6 = (~(J227x6 | Dte7z6[15]));
assign J227x6 = (~(Dte7z6[17] & Dte7z6[16]));
assign Bqziw6 = (!Kz17x6);
assign Kz17x6 = (Nzz6x6 | Dte7z6[13]);
assign Nzz6x6 = (!Dte7z6[14]);
assign Tdtiw6 = (!E4lhw6);
assign Wdqiy6 = (~(Ubhdt6 & Uqkiy6));
assign Uqkiy6 = (~(Gtqiy6 | Awkiy6));
assign Awkiy6 = (~(Otqiy6 & K537x6));
assign K537x6 = (Wtqiy6 ? Xwe7z6[0] : Oac7z6[0]);
assign Otqiy6 = (Z937x6 & X837x6);
assign X837x6 = (Wtqiy6 ? Xwe7z6[3] : Oac7z6[3]);
assign Z937x6 = (Euqiy6 ? Oac7z6[2] : Xwe7z6[2]);
assign Gtqiy6 = (B437x6 | Qg2nv6);
assign B437x6 = (Euqiy6 ? Oac7z6[1] : Xwe7z6[1]);
assign Euqiy6 = (!Wtqiy6);
assign Wtqiy6 = (~(Muqiy6 & Q8iiy6));
assign Q8iiy6 = (~(M5aov6 & R4aov6));
assign Muqiy6 = (~(Ehgdt6 & Uuqiy6));
assign Uuqiy6 = (~(Pbtiw6 & E4lhw6));
assign E4lhw6 = (~(Cvqiy6 & Ngxxx6));
assign Ngxxx6 = (R4aov6 & D4aov6);
assign D4aov6 = (!Bdf7z6[2]);
assign R4aov6 = (!Bdf7z6[0]);
assign Cvqiy6 = (Bdf7z6[1] & Bdf7z6[3]);
assign Pbtiw6 = (!Notiw6);
assign Notiw6 = (M5aov6 & K4aov6);
assign K4aov6 = (!Bdf7z6[1]);
assign M5aov6 = (Bdf7z6[2] & Ju27x6);
assign Ju27x6 = (!Bdf7z6[3]);
assign Ycqiy6 = (Ubhdt6 & Pxfov6);
assign Cgsiw6 = (Kvqiy6 & Svqiy6);
assign Svqiy6 = (~(Awqiy6 | Wpoiy6));
assign Wpoiy6 = (~(Iwqiy6 | Wtoiy6));
assign Wtoiy6 = (!Z8c7z6[3]);
assign Iwqiy6 = (~(Z8c7z6[2] & Z8c7z6[0]));
assign Awqiy6 = (Qwqiy6 & Xvlhw6);
assign Xvlhw6 = (Ywqiy6 & C8onv6);
assign C8onv6 = (~(Vulhw6 & Gxqiy6));
assign Vulhw6 = (~(Zilhw6 | Vsnov6));
assign Vsnov6 = (Oxqiy6 & Gxqiy6);
assign Oxqiy6 = (Kssov6 & Uqd7z6[17]);
assign Zilhw6 = (Wxqiy6 & Ijtov6);
assign Ijtov6 = (Eyqiy6 & Hftov6);
assign Eyqiy6 = (Uqd7z6[18] & Fjohw6);
assign Wxqiy6 = (Gxqiy6 & Qjwiw6);
assign Gxqiy6 = (Myqiy6 & Uyqiy6);
assign Uyqiy6 = (Buihw6 & Qtnov6);
assign Myqiy6 = (Czqiy6 & Kzqiy6);
assign Ywqiy6 = (~(Szqiy6 & A0riy6));
assign A0riy6 = (~(I0riy6 | Q0riy6));
assign Szqiy6 = (~(Y0riy6 | G1riy6));
assign Qwqiy6 = (O1riy6 & Zplhw6);
assign Zplhw6 = (~(Oulhw6 & W1riy6));
assign Oulhw6 = (~(Silhw6 | Jtnov6));
assign Jtnov6 = (E2riy6 & W1riy6);
assign E2riy6 = (E3fhw6 & Xeinv6);
assign Silhw6 = (M2riy6 & U2riy6);
assign U2riy6 = (Qtnov6 & Zpehw6);
assign M2riy6 = (Ttehw6 & W1riy6);
assign W1riy6 = (~(C3riy6 | K3riy6));
assign C3riy6 = (~(Z3fhw6 & S3riy6));
assign O1riy6 = (~(A4riy6 & I4riy6));
assign I4riy6 = (Q4riy6 & E6jiy6);
assign E6jiy6 = (~(Dte7z6[18] | Dte7z6[19]));
assign Q4riy6 = (W4onv6 & A2sov6);
assign W4onv6 = (~(Y4riy6 & Z3fhw6));
assign Y4riy6 = (S3riy6 & K3riy6);
assign A4riy6 = (G5riy6 & M6jiy6);
assign M6jiy6 = (O5riy6 & W5riy6);
assign W5riy6 = (Wqfov6 & Drfov6);
assign O5riy6 = (E6riy6 & M6riy6);
assign M6riy6 = (~(U6riy6 & Ohe7z6[6]));
assign U6riy6 = (Ohe7z6[5] & Ohe7z6[7]);
assign E6riy6 = (~(C7riy6 ^ K7riy6));
assign K7riy6 = (N0gdt6 ^ Ohe7z6[4]);
assign G5riy6 = (Buxxx6 & Z9onv6);
assign Z9onv6 = (~(S7riy6 & Z3fhw6));
assign S7riy6 = (I5fhw6 & Bainv6);
assign Buxxx6 = (~(Ii9ov6 & Kvbov6));
assign Kvbov6 = (!T3cdt6);
assign Kvqiy6 = (Uyoiy6 & A8riy6);
assign A8riy6 = (~(I8riy6 & Gtiiy6));
assign Gtiiy6 = (Q8riy6 & Y8riy6);
assign Y8riy6 = (G9riy6 & Adohw6);
assign G9riy6 = (~(O9riy6 & W9riy6));
assign W9riy6 = (Eariy6 & Mariy6);
assign Mariy6 = (!Zec7z6[19]);
assign Eariy6 = (!Zec7z6[18]);
assign O9riy6 = (Uariy6 & Cbriy6);
assign Cbriy6 = (!Zec7z6[17]);
assign Uariy6 = (!Zec7z6[16]);
assign I8riy6 = (Uiiiy6 & Kbriy6);
assign Uiiiy6 = (Sbriy6 & Zec7z6[25]);
assign Sbriy6 = (Ubsiw6 & Zec7z6[31]);
assign Uyoiy6 = (Acriy6 & Icriy6);
assign Icriy6 = (Qcriy6 & Vzvnv6);
assign Vzvnv6 = (!Zgadt6);
assign Qcriy6 = (Qg2nv6 & C0wnv6);
assign C0wnv6 = (!Nneet6);
assign Acriy6 = (W6u6x6 & Mjhov6);
assign Tka7x6 = (~(Mulnv6 & Oxpiy6));
assign Qgoiy6 = (~(Tiphw6 & Ycriy6));
assign Ycriy6 = (~(Hbo7v6 & Cziiy6));
assign Hbo7v6 = (!Y3jnv6);
assign Icoiy6 = (Gdriy6 & Odriy6);
assign Odriy6 = (Wdriy6 & Eeriy6);
assign Eeriy6 = (~(Meriy6 & Kioov6));
assign Meriy6 = (Ueriy6 & Cfriy6);
assign Cfriy6 = (~(Kfriy6 & Dwb7z6[5]));
assign Kfriy6 = (Lxydt6 & Uvvnv6);
assign Ueriy6 = (~(Dioov6 & Bfo7v6));
assign Wdriy6 = (Sfriy6 & Agriy6);
assign Agriy6 = (~(Bhoov6 & Y3jnv6));
assign Y3jnv6 = (~(Igriy6 & Qgriy6));
assign Qgriy6 = (Ygriy6 & G2oov6);
assign G2oov6 = (!Iladt6);
assign Ygriy6 = (~(U5u6x6 & M7mov6));
assign Igriy6 = (P6u6x6 & Ghriy6);
assign Ghriy6 = (~(Lqfxx6 & Eqfxx6));
assign Eqfxx6 = (~(Z1oov6 & V4jhw6));
assign Sfriy6 = (~(Dwb7z6[1] & Ohriy6));
assign Ohriy6 = (~(Sga7x6 & Zna7x6));
assign Sga7x6 = (!Dioov6);
assign Gdriy6 = (Whriy6 & Eiriy6);
assign Eiriy6 = (Dwb7z6[4] ? Uiriy6 : Miriy6);
assign Uiriy6 = (~(Dwb7z6[0] & Cjriy6));
assign Cjriy6 = (~(Dwb7z6[2] & Lxydt6));
assign Miriy6 = (~(Kjriy6 & Sjriy6));
assign Sjriy6 = (Dioov6 & Akriy6);
assign Akriy6 = (~(Pdlhw6 & Qg2nv6));
assign Kjriy6 = (J8a7x6 & Bh2et6);
assign J8a7x6 = (Ikriy6 & Ntg7z6[3]);
assign Ikriy6 = (Ntg7z6[2] & Ntg7z6[0]);
assign Whriy6 = (Qkriy6 & Ykriy6);
assign Ykriy6 = (~(Glriy6 & Luvnv6));
assign Glriy6 = (~(Olriy6 & Wlriy6));
assign Wlriy6 = (~(Emriy6 & Mmriy6));
assign Emriy6 = (~(Bfo7v6 & Gvvnv6));
assign Olriy6 = (Umriy6 & Cnriy6);
assign Cnriy6 = (~(Bhoov6 & Knriy6));
assign Knriy6 = (~(Uuinv6 & O5a7z6));
assign Uuinv6 = (~(Dwinv6 | Iga7z6));
assign Dwinv6 = (!Cziiy6);
assign Cziiy6 = (~(Snriy6 & Aoriy6));
assign Aoriy6 = (Ioriy6 & Qoriy6);
assign Qoriy6 = (Brriw6 | Yoriy6);
assign Yoriy6 = (Gpriy6 & Yzriw6);
assign Yzriw6 = (Opriy6 & Mjq6x6);
assign Mjq6x6 = (!Zeihw6);
assign Zeihw6 = (~(Wpriy6 & Eqriy6));
assign Eqriy6 = (Mqriy6 & Uqriy6);
assign Uqriy6 = (Crriy6 & Krriy6);
assign Krriy6 = (~(Zec7z6[0] & Srriy6));
assign Mqriy6 = (Asriy6 & Isriy6);
assign Isriy6 = (Wkriw6 | Fcinv6);
assign Asriy6 = (~(Ovbdt6 & Qsriy6));
assign Wpriy6 = (Ysriy6 & Gtriy6);
assign Gtriy6 = (Otriy6 & Wtriy6);
assign Wtriy6 = (~(Mynhw6 & Zec7z6[24]));
assign Otriy6 = (U2ohw6 | Qvlhw6);
assign Ysriy6 = (Qsoiy6 & E7phw6);
assign Qsoiy6 = (Euriy6 & Muriy6);
assign Muriy6 = (Uuriy6 & Cvriy6);
assign Cvriy6 = (~(Kvriy6 & Zec7z6[8]));
assign Uuriy6 = (Svriy6 & G1kxx6);
assign Svriy6 = (~(Zec7z6[0] & Gdpiy6));
assign Euriy6 = (Awriy6 & Iwriy6);
assign Iwriy6 = (Ctnov6 | Y447x6);
assign Awriy6 = (Qwriy6 & Ywriy6);
assign Ywriy6 = (Gxriy6 | Kfa7z6);
assign Qwriy6 = (~(Vuehw6 & Zec7z6[6]));
assign Opriy6 = (Nfihw6 & Xdihw6);
assign Xdihw6 = (~(Oxriy6 & Wxriy6));
assign Wxriy6 = (Eyriy6 & Myriy6);
assign Myriy6 = (Crriy6 & Uyriy6);
assign Uyriy6 = (~(Zec7z6[2] & Srriy6));
assign Eyriy6 = (Czriy6 & Kzriy6);
assign Kzriy6 = (Wkriw6 | Bainv6);
assign Czriy6 = (~(Uqd7z6[18] & Qsriy6));
assign Oxriy6 = (Szriy6 & A0siy6);
assign A0siy6 = (I0siy6 & Q0siy6);
assign Q0siy6 = (~(Mynhw6 & Zec7z6[26]));
assign I0siy6 = (Zpehw6 | Qvlhw6);
assign Szriy6 = (Otoiy6 & E7phw6);
assign Otoiy6 = (Y0siy6 & G1siy6);
assign G1siy6 = (O1siy6 & W1siy6);
assign W1siy6 = (Adohw6 | Gxriy6);
assign O1siy6 = (E2siy6 & G1kxx6);
assign E2siy6 = (~(Zec7z6[2] & Gdpiy6));
assign Y0siy6 = (M2siy6 & U2siy6);
assign U2siy6 = (Jbqiw6 | Y447x6);
assign M2siy6 = (C3siy6 & K3siy6);
assign K3siy6 = (~(Kvriy6 & Zec7z6[10]));
assign C3siy6 = (~(Vuehw6 & Zec7z6[8]));
assign Nfihw6 = (~(S3siy6 & A4siy6));
assign A4siy6 = (I4siy6 & Q4siy6);
assign Q4siy6 = (Crriy6 & G1kxx6);
assign Crriy6 = (Onlhw6 & I1wiw6);
assign I4siy6 = (Y4siy6 & G5siy6);
assign G5siy6 = (~(Zec7z6[3] & O5siy6));
assign O5siy6 = (~(Mquiw6 & Hffhw6));
assign Mquiw6 = (~(Bvuiw6 | V0nhw6));
assign Y4siy6 = (~(Uqd7z6[19] & Qsriy6));
assign S3siy6 = (W5siy6 & E6siy6);
assign E6siy6 = (M6siy6 & U6siy6);
assign U6siy6 = (~(Mynhw6 & Zec7z6[27]));
assign M6siy6 = (~(Zec7z6[6] & C7siy6));
assign C7siy6 = (K7siy6 | G5sov6);
assign G5sov6 = (!Amtov6);
assign W5siy6 = (Euoiy6 & E7phw6);
assign Euoiy6 = (S7siy6 & A8siy6);
assign A8siy6 = (Fjohw6 | Y447x6);
assign S7siy6 = (Elviw6 | Gxriy6);
assign Gpriy6 = (Ltq6x6 & F4ihw6);
assign F4ihw6 = (~(I8siy6 & Q8siy6));
assign Q8siy6 = (Y8siy6 & G9siy6);
assign G9siy6 = (O9siy6 & I1wiw6);
assign O9siy6 = (Qtnov6 | Qvlhw6);
assign Y8siy6 = (W9siy6 & Easiy6);
assign Easiy6 = (~(Uqd7z6[17] & Qsriy6));
assign W9siy6 = (Wkriw6 | Xeinv6);
assign I8siy6 = (Masiy6 & Uasiy6);
assign Uasiy6 = (Cbsiy6 & Kbsiy6);
assign Kbsiy6 = (~(Mynhw6 & Zec7z6[25]));
assign Cbsiy6 = (~(Zec7z6[1] & Srriy6));
assign Srriy6 = (~(Sbsiy6 & A7onv6));
assign Masiy6 = (Uuoiy6 & E7phw6);
assign Uuoiy6 = (Acsiy6 & Icsiy6);
assign Icsiy6 = (Qcsiy6 & Ycsiy6);
assign Ycsiy6 = (~(Kvriy6 & Zec7z6[9]));
assign Qcsiy6 = (Gdsiy6 & G1kxx6);
assign Gdsiy6 = (~(Zec7z6[1] & Gdpiy6));
assign Acsiy6 = (Odsiy6 & Wdsiy6);
assign Wdsiy6 = (Jgtov6 | Y447x6);
assign Odsiy6 = (Eesiy6 & Mesiy6);
assign Mesiy6 = (Gxriy6 | Bat8v6);
assign Bat8v6 = (!M6nhw6);
assign Eesiy6 = (~(Vuehw6 & Zec7z6[7]));
assign Ltq6x6 = (~(Uesiy6 & Cfsiy6));
assign Cfsiy6 = (Kfsiy6 & Sfsiy6);
assign Sfsiy6 = (Agsiy6 & Igsiy6);
assign Igsiy6 = (Wkriw6 & Irsov6);
assign Agsiy6 = (~(Gxriw6 | Bmwiw6));
assign Bmwiw6 = (!M6onv6);
assign Gxriw6 = (Vuehw6 & Qgsiy6);
assign Qgsiy6 = (~(Gginv6 & Ygsiy6));
assign Ygsiy6 = (!Cvehw6);
assign Kfsiy6 = (Ghsiy6 & Ohsiy6);
assign Ohsiy6 = (~(Rzriw6 & Gginv6));
assign Rzriw6 = (~(Nrqiw6 & Whsiy6));
assign Ghsiy6 = (Eisiy6 & F0fhw6);
assign Eisiy6 = (~(V0nhw6 & Misiy6));
assign Misiy6 = (~(Hwpiw6 & E3fhw6));
assign Hwpiw6 = (!Mxuiw6);
assign Mxuiw6 = (~(Uisiy6 & D4ohw6));
assign D4ohw6 = (~(M6nhw6 | Z9nhw6));
assign Uisiy6 = (Nqlhw6 & Adohw6);
assign Uesiy6 = (Cjsiy6 & Kjsiy6);
assign Kjsiy6 = (Sjsiy6 & Aksiy6);
assign Aksiy6 = (Iksiy6 & Qksiy6);
assign Qksiy6 = (~(Yksiy6 & Kzriw6));
assign Iksiy6 = (~(Auehw6 & Rktov6));
assign Sjsiy6 = (Bouiw6 & Sbsiy6);
assign Sbsiy6 = (Glsiy6 & Smuiw6);
assign Smuiw6 = (Buviw6 & Dssov6);
assign Glsiy6 = (Hffhw6 & A2sov6);
assign Hffhw6 = (~(Olsiy6 & Wlsiy6));
assign Wlsiy6 = (Lofhw6 & Buihw6);
assign Olsiy6 = (Emsiy6 & Hxviw6);
assign Bouiw6 = (Mmsiy6 & Nqehw6);
assign Mmsiy6 = (T6onv6 & D0riw6);
assign Cjsiy6 = (Umsiy6 & Jvriw6);
assign Umsiy6 = (Qvlhw6 & Cgfhw6);
assign Cgfhw6 = (Cnsiy6 & Knsiy6);
assign Knsiy6 = (Snsiy6 & Onlhw6);
assign Onlhw6 = (!P3vxx6);
assign Snsiy6 = (I1wiw6 & Vnlhw6);
assign Cnsiy6 = (Gqehw6 & Aosiy6);
assign Aosiy6 = (~(Rdfhw6 & Yksiy6));
assign Rdfhw6 = (!Nrqiw6);
assign Qvlhw6 = (Iosiy6 & Emiiy6);
assign Iosiy6 = (C3riw6 & Amtov6);
assign C3riw6 = (Qosiy6 & Yosiy6);
assign Yosiy6 = (~(Gpsiy6 & Yksiy6));
assign Qosiy6 = (Ayuiw6 & Stuiw6);
assign Stuiw6 = (~(Opsiy6 & Wpsiy6));
assign Opsiy6 = (Gginv6 & Eqsiy6);
assign Ayuiw6 = (~(Gpsiy6 & Ydfhw6));
assign Gpsiy6 = (Mqsiy6 & Uqsiy6);
assign Brriw6 = (Crsiy6 & Npfhw6);
assign Npfhw6 = (~(B2xxx6 | Eofhw6));
assign Eofhw6 = (!Sofhw6);
assign Sofhw6 = (~(Krsiy6 & Srsiy6));
assign Srsiy6 = (Assiy6 & Issiy6);
assign Issiy6 = (Qssiy6 & Yssiy6);
assign Yssiy6 = (~(Zec7z6[4] & Nxlhw6));
assign Qssiy6 = (Gtsiy6 & Z0kxx6);
assign Gtsiy6 = (~(Zec7z6[9] & Oipiw6));
assign Assiy6 = (Otsiy6 & Wtsiy6);
assign Wtsiy6 = (S8ohw6 | D447x6);
assign Otsiy6 = (~(Bvuiw6 & Uqd7z6[17]));
assign Krsiy6 = (Eusiy6 & Musiy6);
assign Musiy6 = (~(Iwoiy6 | Uusiy6));
assign Uusiy6 = (~(A7onv6 | Buihw6));
assign Iwoiy6 = (~(Cvsiy6 & Kvsiy6));
assign Kvsiy6 = (Svsiy6 & G1kxx6);
assign Svsiy6 = (~(Zec7z6[4] & Cniiy6));
assign Cvsiy6 = (Awsiy6 & Iwsiy6);
assign Iwsiy6 = (~(Zec7z6[1] & Qwsiy6));
assign Awsiy6 = (~(Odpiy6 & Zec7z6[9]));
assign Eusiy6 = (Asiiy6 & Jvlhw6);
assign Asiiy6 = (Hulhw6 & Ywsiy6);
assign Ywsiy6 = (S8ohw6 | Emiiy6);
assign B2xxx6 = (!Xnfhw6);
assign Xnfhw6 = (Gxsiy6 & Oxsiy6);
assign Oxsiy6 = (Wxsiy6 & Eysiy6);
assign Eysiy6 = (Mysiy6 & Uysiy6);
assign Uysiy6 = (~(Zec7z6[0] & Czsiy6));
assign Mysiy6 = (~(Zec7z6[8] & Oipiw6));
assign Wxsiy6 = (Kzsiy6 & Szsiy6);
assign Szsiy6 = (~(Bvuiw6 & Ovbdt6));
assign Kzsiy6 = (~(V0nhw6 & Zec7z6[24]));
assign Gxsiy6 = (A0tiy6 & I0tiy6);
assign A0tiy6 = (~(Ywoiy6 | Q0tiy6));
assign Q0tiy6 = (Zec7z6[3] & Nxlhw6);
assign Ywoiy6 = (~(Y0tiy6 & G1tiy6));
assign G1tiy6 = (O1tiy6 & W1tiy6);
assign W1tiy6 = (~(Zec7z6[3] & Cniiy6));
assign O1tiy6 = (~(Zec7z6[0] & Qwsiy6));
assign Y0tiy6 = (Fefhw6 & E2tiy6);
assign E2tiy6 = (~(Odpiy6 & Zec7z6[8]));
assign Crsiy6 = (Omfhw6 & Rrfhw6);
assign Rrfhw6 = (~(M2tiy6 & U2tiy6));
assign U2tiy6 = (C3tiy6 & K3tiy6);
assign K3tiy6 = (S3tiy6 & A4tiy6);
assign A4tiy6 = (~(Zec7z6[2] & Czsiy6));
assign Czsiy6 = (~(D447x6 & Emiiy6));
assign Emiiy6 = (I4tiy6 & Q4tiy6);
assign Q4tiy6 = (~(K7siy6 | Mtehw6));
assign Mtehw6 = (Zrwiw6 & V1fhw6);
assign I4tiy6 = (K4uiw6 & Anriw6);
assign Anriw6 = (Y4tiy6 & G5tiy6);
assign G5tiy6 = (O5tiy6 & Uh37x6);
assign Uh37x6 = (~(W5tiy6 & Obwiw6));
assign O5tiy6 = (Lpsov6 & Xhriw6);
assign Xhriw6 = (~(E6tiy6 & M6tiy6));
assign Lpsov6 = (!Gh37x6);
assign Gh37x6 = (M6tiy6 & Oyuiw6);
assign Y4tiy6 = (U6tiy6 & Ydsiw6);
assign Ydsiw6 = (C7tiy6 & K7tiy6);
assign K7tiy6 = (S7tiy6 & A4wiw6);
assign A4wiw6 = (~(Hyuiw6 & P5fhw6));
assign S7tiy6 = (Ldwiw6 & H4wiw6);
assign H4wiw6 = (~(E6tiy6 & Hyuiw6));
assign Ldwiw6 = (~(W5tiy6 & Sywiw6));
assign C7tiy6 = (Ekwiw6 & Wdriw6);
assign Wdriw6 = (~(A8tiy6 | Q6viw6));
assign Q6viw6 = (I8tiy6 & Hyuiw6);
assign I8tiy6 = (Sywiw6 & Fcinv6);
assign A8tiy6 = (Hyuiw6 & Q8tiy6);
assign Ekwiw6 = (Y8tiy6 & G2uiw6);
assign G2uiw6 = (!Zbsov6);
assign Zbsov6 = (Q8tiy6 & M6tiy6);
assign Q8tiy6 = (~(G9tiy6 | Bainv6));
assign G9tiy6 = (!Ttehw6);
assign Y8tiy6 = (~(W5tiy6 & B0xiw6));
assign W5tiy6 = (M6tiy6 & Fcinv6);
assign U6tiy6 = (X9fhw6 & Epsov6);
assign Epsov6 = (~(M6tiy6 & P5fhw6));
assign X9fhw6 = (~(O9tiy6 & M6tiy6));
assign M6tiy6 = (W9tiy6 & V1fhw6);
assign K4uiw6 = (Eatiy6 & Matiy6);
assign Matiy6 = (~(P5fhw6 & Uatiy6));
assign P5fhw6 = (~(M2xiw6 | Zec7z6[6]));
assign M2xiw6 = (!Zdwiw6);
assign Eatiy6 = (Pyehw6 & N4fhw6);
assign N4fhw6 = (~(Uatiy6 & Oyuiw6));
assign Oyuiw6 = (Obwiw6 & Zec7z6[6]);
assign Pyehw6 = (~(E6tiy6 & Uatiy6));
assign Uatiy6 = (Cbtiy6 & V1fhw6);
assign Cbtiy6 = (I5fhw6 & Zec7z6[11]);
assign E6tiy6 = (Ttehw6 & Bainv6);
assign Ttehw6 = (~(Fcinv6 | Zec7z6[7]));
assign S3tiy6 = (~(Zec7z6[10] & Oipiw6));
assign Oipiw6 = (!Aulhw6);
assign Aulhw6 = (~(Nh37x6 | V8fhw6));
assign V8fhw6 = (~(W5siw6 | Kbtiy6));
assign Nh37x6 = (~(W5siw6 | Yksiy6));
assign W5siw6 = (~(Mqsiy6 & Zec7z6[13]));
assign Mqsiy6 = (Sbtiy6 & Eqsiy6);
assign C3tiy6 = (Actiy6 & Ictiy6);
assign Ictiy6 = (~(Bvuiw6 & Uqd7z6[18]));
assign Actiy6 = (~(V0nhw6 & Zec7z6[26]));
assign M2tiy6 = (Qctiy6 & I0tiy6);
assign Qctiy6 = (~(Myoiy6 | Yctiy6));
assign Yctiy6 = (Zec7z6[5] & Nxlhw6);
assign Nxlhw6 = (~(Gdtiy6 & Buviw6));
assign Buviw6 = (Odtiy6 & Wdtiy6);
assign Wdtiy6 = (~(Hyuiw6 & Obwiw6));
assign Odtiy6 = (Xzuiw6 & Ltuiw6);
assign Ltuiw6 = (~(Eetiy6 & Hyuiw6));
assign Eetiy6 = (B0xiw6 & Fcinv6);
assign Xzuiw6 = (~(O9tiy6 & Hyuiw6));
assign Hyuiw6 = (W9tiy6 & Kdfhw6);
assign O9tiy6 = (Sywiw6 & Zec7z6[6]);
assign Gdtiy6 = (V2riw6 & Wkriw6);
assign Wkriw6 = (~(Zafhw6 & Metiy6));
assign Metiy6 = (Kdfhw6 | V1fhw6);
assign V2riw6 = (Uetiy6 & C6viw6);
assign C6viw6 = (~(Cftiy6 & Z3fhw6));
assign Cftiy6 = (Wpsiy6 & Eqsiy6);
assign Uetiy6 = (~(Zafhw6 & Gbfhw6));
assign Zafhw6 = (Kftiy6 & Wpsiy6);
assign Kftiy6 = (Zec7z6[11] & Eqsiy6);
assign Myoiy6 = (~(Sftiy6 & Agtiy6));
assign Agtiy6 = (Igtiy6 & Qgtiy6);
assign Qgtiy6 = (~(Odpiy6 & Zec7z6[10]));
assign Odpiy6 = (!O8fhw6);
assign Igtiy6 = (~(Zec7z6[5] & Cniiy6));
assign Cniiy6 = (!I4ghw6);
assign Sftiy6 = (Fefhw6 & Ygtiy6);
assign Ygtiy6 = (~(Zec7z6[2] & Qwsiy6));
assign Omfhw6 = (!Wqfhw6);
assign Wqfhw6 = (Ghtiy6 & Ohtiy6);
assign Ohtiy6 = (Whtiy6 & Eitiy6);
assign Eitiy6 = (~(V0nhw6 & Zec7z6[27]));
assign V0nhw6 = (!A7onv6);
assign Whtiy6 = (Mitiy6 & R447x6);
assign R447x6 = (~(Zec7z6[7] & K7siy6));
assign K7siy6 = (~(Uitiy6 & Cjtiy6));
assign Cjtiy6 = (Q9fhw6 & Kjtiy6);
assign Uitiy6 = (Rlriw6 & B5siw6);
assign B5siw6 = (~(Sjtiy6 & Aktiy6));
assign Rlriw6 = (~(Iktiy6 & W9tiy6));
assign Iktiy6 = (Gbfhw6 & Zec7z6[8]);
assign Mitiy6 = (~(Bvuiw6 & Uqd7z6[19]));
assign Bvuiw6 = (!Dssov6);
assign Dssov6 = (~(Qktiy6 & Yktiy6));
assign Qktiy6 = (Qjwiw6 & Xeinv6);
assign Ghtiy6 = (Gltiy6 & I0tiy6);
assign I0tiy6 = (Oltiy6 & Jvlhw6);
assign Jvlhw6 = (S9nhw6 & I1wiw6);
assign I1wiw6 = (~(Wltiy6 & Gqlhw6));
assign Gqlhw6 = (Emtiy6 & Uqd7z6[21]);
assign Emtiy6 = (Jolhw6 & E9onv6);
assign Jolhw6 = (Czqiy6 & Zec7z6[4]);
assign Czqiy6 = (Mmtiy6 & Erwiw6);
assign Erwiw6 = (E3fhw6 & Sywiw6);
assign Mmtiy6 = (Umtiy6 & V1fhw6);
assign Wltiy6 = (Uqd7z6[22] & Sfa7z6);
assign Oltiy6 = (Wcsiw6 & Ddsiw6);
assign Ddsiw6 = (Cntiy6 & Z0kxx6);
assign Z0kxx6 = (Kbtiy6 | Kntiy6);
assign Cntiy6 = (~(Sntiy6 & Ydfhw6));
assign Wcsiw6 = (Hulhw6 & Hcviw6);
assign Hcviw6 = (~(Zrwiw6 & Kdfhw6));
assign Zrwiw6 = (Aotiy6 & I5fhw6);
assign Aotiy6 = (Gginv6 & Bainv6);
assign Hulhw6 = (E7phw6 & A2sov6);
assign E7phw6 = (Sfohw6 & T1sov6);
assign Gltiy6 = (~(Wxoiy6 | Iotiy6));
assign Iotiy6 = (~(U2ohw6 | D447x6));
assign D447x6 = (Qotiy6 & Irsov6);
assign Qotiy6 = (!Qsriy6);
assign Qsriy6 = (~(Yotiy6 & Gptiy6));
assign Gptiy6 = (~(Kvviw6 | X8onv6));
assign X8onv6 = (!Vnlhw6);
assign Vnlhw6 = (~(Optiy6 & Wptiy6));
assign Wptiy6 = (Eqtiy6 & Kktov6);
assign Eqtiy6 = (Hxviw6 & Qtnov6);
assign Optiy6 = (Mqtiy6 & Zec7z6[9]);
assign Mqtiy6 = (~(Y1xiw6 | I0riy6));
assign Y1xiw6 = (!B0xiw6);
assign Yotiy6 = (Inviw6 & M6onv6);
assign M6onv6 = (~(Uqtiy6 & Crtiy6));
assign Crtiy6 = (Krtiy6 & Oenhw6);
assign Krtiy6 = (Glpiw6 & Fcinv6);
assign Uqtiy6 = (Yktiy6 & Zec7z6[7]);
assign Inviw6 = (Srtiy6 & Astiy6);
assign Astiy6 = (Istiy6 & T6onv6);
assign T6onv6 = (~(Qstiy6 & Ystiy6));
assign Ystiy6 = (Oenhw6 & Xeinv6);
assign Qstiy6 = (Yktiy6 & K0riw6);
assign Yktiy6 = (Gttiy6 & Ottiy6);
assign Ottiy6 = (~(I0riy6 | Zec7z6[8]));
assign Gttiy6 = (Q8onv6 & Zec7z6[9]);
assign Istiy6 = (Prsov6 & L4riw6);
assign Srtiy6 = (Wttiy6 & Gqehw6);
assign Gqehw6 = (~(Xjwiw6 | S6wiw6));
assign S6wiw6 = (Eutiy6 & Mutiy6);
assign Mutiy6 = (Uutiy6 & Zec7z6[6]);
assign Uutiy6 = (~(I0riy6 | Zec7z6[4]));
assign Eutiy6 = (Qjwiw6 & Cvtiy6);
assign Xjwiw6 = (Kvtiy6 & Svtiy6);
assign Kvtiy6 = (Qjwiw6 & Qtnov6);
assign Wttiy6 = (Awtiy6 & Nqehw6);
assign Nqehw6 = (~(Iwtiy6 & Qwtiy6));
assign Qwtiy6 = (Ywtiy6 & Svtiy6);
assign Svtiy6 = (Gxtiy6 & Cvtiy6);
assign Gxtiy6 = (~(I0riy6 | Zec7z6[6]));
assign Ywtiy6 = (Zec7z6[4] & Uqd7z6[22]);
assign Iwtiy6 = (Uqd7z6[20] & Fqohw6);
assign Fqohw6 = (Uqd7z6[21] & Oenhw6);
assign Awtiy6 = (D0riw6 | Kvviw6);
assign D0riw6 = (!Owpiw6);
assign Wxoiy6 = (~(Fefhw6 & Oxtiy6));
assign Oxtiy6 = (~(Zec7z6[3] & Qwsiy6));
assign Qwsiy6 = (~(Y447x6 & Gxriy6));
assign Gxriy6 = (F547x6 & W347x6);
assign W347x6 = (!Igviw6);
assign Igviw6 = (~(Rsriw6 & Wxtiy6));
assign Wxtiy6 = (~(Eytiy6 & Qtnov6));
assign Rsriw6 = (Cvmiy6 & Mytiy6);
assign F547x6 = (!Pgviw6);
assign Pgviw6 = (~(Uytiy6 & Cztiy6));
assign Cztiy6 = (~(Eytiy6 & Zec7z6[4]));
assign Uytiy6 = (Kztiy6 & Sztiy6);
assign Kztiy6 = (~(Auehw6 & A0uiy6));
assign Y447x6 = (F0fhw6 & I0uiy6);
assign I0uiy6 = (~(Wdpiy6 & Auehw6));
assign Wdpiy6 = (!A0uiy6);
assign A0uiy6 = (~(Q0uiy6 & Y0uiy6));
assign Y0uiy6 = (G1uiy6 & O1uiy6);
assign O1uiy6 = (W1uiy6 & L4riw6);
assign L4riw6 = (~(E2uiy6 & M2uiy6));
assign E2uiy6 = (Elviw6 & Qeinv6);
assign W1uiy6 = (~(I2phw6 | Eytiy6));
assign Eytiy6 = (!Yzehw6);
assign I2phw6 = (~(T1riw6 | U2uiy6));
assign G1uiy6 = (~(Mynhw6 | Kvviw6));
assign Kvviw6 = (C3uiy6 & Lzviw6);
assign Lzviw6 = (Zdwiw6 & Nbfhw6);
assign C3uiy6 = (Owpiw6 & K0riw6);
assign Owpiw6 = (V1fhw6 & Zhmhw6);
assign V1fhw6 = (Zec7z6[9] & Painv6);
assign Mynhw6 = (!Irsov6);
assign Irsov6 = (~(K3uiy6 & S3uiy6));
assign K3uiy6 = (Zec7z6[6] & Bainv6);
assign Q0uiy6 = (A4uiy6 & I4uiy6);
assign I4uiy6 = (~(Q4uiy6 | Axihw6));
assign Axihw6 = (Auehw6 & Zec7z6[27]);
assign Q4uiy6 = (P3vxx6 & Y4uiy6);
assign Y4uiy6 = (~(M7siw6 & G5uiy6));
assign G5uiy6 = (~(Ehtov6 & F4vxx6));
assign F4vxx6 = (O5uiy6 & Qjwiw6);
assign O5uiy6 = (Uqd7z6[19] & Jbqiw6);
assign Ehtov6 = (Uqd7z6[17] & Ctnov6);
assign M7siw6 = (N99iw6 | Tnzdt6);
assign P3vxx6 = (Qzuiw6 & Emsiy6);
assign Emsiy6 = (!Fquiw6);
assign Fquiw6 = (~(W5uiy6 & E6uiy6));
assign E6uiy6 = (M6uiy6 & U6uiy6);
assign M6uiy6 = (Kfa7z6 & Qtnov6);
assign W5uiy6 = (H2riw6 & Cvtiy6);
assign A4uiy6 = (Oe37x6 & Mefhw6);
assign Mefhw6 = (B2phw6 & Cvmiy6);
assign B2phw6 = (Mytiy6 & Sztiy6);
assign Oe37x6 = (C7uiy6 & S9nhw6);
assign S9nhw6 = (~(L4sov6 | Wpnhw6));
assign Wpnhw6 = (Umtiy6 & K7uiy6);
assign Umtiy6 = (S7uiy6 & U6uiy6);
assign S7uiy6 = (Kfa7z6 & Adohw6);
assign L4sov6 = (U6uiy6 & Z9nhw6);
assign C7uiy6 = (Prsov6 & A7onv6);
assign A7onv6 = (~(A8uiy6 & S3uiy6));
assign A8uiy6 = (Zec7z6[8] & Qtnov6);
assign Prsov6 = (~(I8uiy6 & S3uiy6));
assign S3uiy6 = (Q8uiy6 & M2uiy6);
assign Q8uiy6 = (Zec7z6[9] & Elviw6);
assign I8uiy6 = (Fcinv6 & Bainv6);
assign Fefhw6 = (~(Ioiiy6 | Mqiiy6));
assign Ioriy6 = (Qalhw6 & Whhov6);
assign Qalhw6 = (~(Y8uiy6 & G9uiy6));
assign G9uiy6 = (Md37x6 & O9uiy6);
assign O9uiy6 = (~(Ryfhw6 & Llyxx6));
assign Llyxx6 = (Qtnov6 | L6wiw6);
assign L6wiw6 = (P8wiw6 & W9uiy6);
assign Ryfhw6 = (!Mytiy6);
assign Mytiy6 = (~(Eauiy6 & Mauiy6));
assign Mauiy6 = (Qzuiw6 | Uauiy6);
assign Uauiy6 = (Zec7z6[6] & Zec7z6[8]);
assign Md37x6 = (F0fhw6 & Kjtiy6);
assign Kjtiy6 = (!Znvnv6);
assign F0fhw6 = (!Nkyxx6);
assign Nkyxx6 = (Cbuiy6 & Kktov6);
assign Y8uiy6 = (Kbuiy6 & Sbuiy6);
assign Sbuiy6 = (!Tlyxx6);
assign Tlyxx6 = (~(Acuiy6 & I4ghw6));
assign I4ghw6 = (~(Gdpiy6 | Vuehw6));
assign Vuehw6 = (~(Icuiy6 | D6siw6));
assign Gdpiy6 = (~(Wyehw6 & Nrqiw6));
assign Nrqiw6 = (~(Qcuiy6 & Zec7z6[14]));
assign Qcuiy6 = (Zec7z6[13] & Eqsiy6);
assign Wyehw6 = (!K1qiw6);
assign K1qiw6 = (Kzriw6 & Ycuiy6);
assign Kzriw6 = (Gduiy6 & Zec7z6[15]);
assign Acuiy6 = (~(Ioiiy6 | Lsihw6));
assign Lsihw6 = (~(Oduiy6 & Wduiy6));
assign Wduiy6 = (Eeuiy6 | Jvriw6);
assign Jvriw6 = (Sztiy6 & Yzehw6);
assign Eeuiy6 = (Zec7z6[4] ? Ueuiy6 : Meuiy6);
assign Meuiy6 = (~(Cfuiy6 & Kfuiy6));
assign Kfuiy6 = (~(Sfuiy6 & Aguiy6));
assign Aguiy6 = (Ovbdt6 & Sztiy6);
assign Sztiy6 = (~(Iguiy6 & Zdwiw6));
assign Zdwiw6 = (Xeinv6 & Bainv6);
assign Iguiy6 = (Eauiy6 & Nbfhw6);
assign Sfuiy6 = (Uqd7z6[19] & Uqd7z6[18]);
assign Cfuiy6 = (~(Ubsiw6 & Yzehw6));
assign Yzehw6 = (~(Qguiy6 & Yguiy6));
assign Yguiy6 = (Nbfhw6 & Qolhw6);
assign Qolhw6 = (Ghuiy6 & Uqd7z6[22]);
assign Ghuiy6 = (Sfa7z6 & Dsehw6);
assign Dsehw6 = (!Uqd7z6[21]);
assign Qguiy6 = (Eauiy6 & Obwiw6);
assign Ubsiw6 = (!P8wiw6);
assign P8wiw6 = (~(Ohuiy6 & Zec7z6[27]));
assign Ohuiy6 = (Zec7z6[26] & Zec7z6[24]);
assign Oduiy6 = (~(Auehw6 & Whuiy6));
assign Whuiy6 = (~(Eiuiy6 & J1ghw6));
assign Eiuiy6 = (~(Yyfhw6 | Lofhw6));
assign Yyfhw6 = (~(Miuiy6 & Uiuiy6));
assign Uiuiy6 = (Cjuiy6 & Kjuiy6);
assign Kjuiy6 = (Z9nhw6 ^ Baohw6);
assign Cjuiy6 = (M6nhw6 ^ S8ohw6);
assign Miuiy6 = (Sjuiy6 & Akuiy6);
assign Akuiy6 = (Zec7z6[2] ^ Adohw6);
assign Sjuiy6 = (Zec7z6[31] ^ U2ohw6);
assign Auehw6 = (!T1riw6);
assign T1riw6 = (~(Ikuiy6 & Qkuiy6));
assign Qkuiy6 = (~(Q0riy6 | Ykuiy6));
assign Ykuiy6 = (!Y0riy6);
assign Y0riy6 = (~(Q8onv6 & Gluiy6));
assign Gluiy6 = (~(Oluiy6 & Zec7z6[4]));
assign Oluiy6 = (~(Hxviw6 | E3fhw6));
assign Q8onv6 = (Ueuiy6 & M6nhw6);
assign M6nhw6 = (Zec7z6[29] & Otiiy6);
assign Ueuiy6 = (!W9uiy6);
assign W9uiy6 = (~(Wluiy6 & Zec7z6[31]));
assign Wluiy6 = (Zec7z6[30] & Z9nhw6);
assign Q0riy6 = (Zec7z6[8] & Emuiy6);
assign Emuiy6 = (Qtnov6 | Nbfhw6);
assign Ikuiy6 = (~(G1riy6 | I0riy6));
assign I0riy6 = (~(Shmhw6 & Painv6));
assign Shmhw6 = (Mmuiy6 & Zec7z6[12]);
assign Mmuiy6 = (Zec7z6[11] & Otiiy6);
assign G1riy6 = (~(Umuiy6 & Cnuiy6));
assign Cnuiy6 = (J1ghw6 | Knuiy6);
assign Knuiy6 = (Snuiy6 & Aouiy6);
assign Aouiy6 = (~(K0riw6 & Qtnov6));
assign Snuiy6 = (Hxihw6 | P2ihw6);
assign P2ihw6 = (Iouiy6 & Qouiy6);
assign Iouiy6 = (Nqlhw6 & Xeinv6);
assign J1ghw6 = (Youiy6 & U2uiy6);
assign Youiy6 = (Zec7z6[27] & Utihw6);
assign Umuiy6 = (~(Qzuiw6 | Zec7z6[9]));
assign Ioiiy6 = (!G3ghw6);
assign G3ghw6 = (Whsiy6 & G1kxx6);
assign G1kxx6 = (!Zwriw6);
assign Zwriw6 = (Ydfhw6 & Gpuiy6);
assign Whsiy6 = (!Kvriy6);
assign Kvriy6 = (Wpsiy6 & Zec7z6[15]);
assign Wpsiy6 = (Gduiy6 & Zec7z6[12]);
assign Gduiy6 = (Uqsiy6 & Sbtiy6);
assign Kbuiy6 = (!Vkyxx6);
assign Vkyxx6 = (~(Opuiy6 & Wpuiy6));
assign Wpuiy6 = (Bylhw6 | Equiy6);
assign Equiy6 = (Mquiy6 & Uquiy6);
assign Uquiy6 = (Qtnov6 & Xeinv6);
assign Qtnov6 = (!Zec7z6[4]);
assign Mquiy6 = (~(K3riy6 | Q2fhw6));
assign Q2fhw6 = (!Hxviw6);
assign Hxviw6 = (Zpehw6 & Fcinv6);
assign K3riy6 = (~(Cruiy6 & Kruiy6));
assign Kruiy6 = (T5ohw6 & U2ohw6);
assign U2ohw6 = (!Zec7z6[3]);
assign T5ohw6 = (!Zec7z6[2]);
assign Cruiy6 = (Baohw6 & S8ohw6);
assign S8ohw6 = (!Zec7z6[1]);
assign Baohw6 = (!Zec7z6[0]);
assign Bylhw6 = (O8fhw6 & Sruiy6);
assign Sruiy6 = (!Mqiiy6);
assign O8fhw6 = (~(Xgmhw6 & Ycuiy6));
assign Ycuiy6 = (~(Jdviw6 & Kbtiy6));
assign Jdviw6 = (!Ydfhw6);
assign Opuiy6 = (Kjmiy6 & Asuiy6);
assign Asuiy6 = (~(Zofhw6 & Isuiy6));
assign Isuiy6 = (~(Qsuiy6 & Ysuiy6));
assign Ysuiy6 = (Gtuiy6 & Kfa7z6);
assign Kfa7z6 = (!Z9nhw6);
assign Z9nhw6 = (Zec7z6[28] & Otiiy6);
assign Gtuiy6 = (Adohw6 & Elviw6);
assign Qsuiy6 = (Otuiy6 & Kssov6);
assign Kssov6 = (Gitov6 & Qjwiw6);
assign Qjwiw6 = (Kktov6 & E9onv6);
assign E9onv6 = (!Uqd7z6[20]);
assign Uqd7z6[20] = (Zec7z6[20] & Otiiy6);
assign Kktov6 = (~(K4ohw6 | Uqd7z6[21]));
assign Uqd7z6[21] = (Zec7z6[21] & Otiiy6);
assign K4ohw6 = (!Nqlhw6);
assign Nqlhw6 = (Glpiw6 & Sfa7z6);
assign Sfa7z6 = (!Oenhw6);
assign Oenhw6 = (Zec7z6[23] & Otiiy6);
assign Glpiw6 = (!Uqd7z6[22]);
assign Uqd7z6[22] = (Zec7z6[22] & Otiiy6);
assign Gitov6 = (Jbqiw6 & Fjohw6);
assign Fjohw6 = (!Uqd7z6[19]);
assign Uqd7z6[19] = (Zec7z6[19] & Otiiy6);
assign Jbqiw6 = (!Uqd7z6[18]);
assign Uqd7z6[18] = (Zec7z6[18] & Otiiy6);
assign Otuiy6 = (Hftov6 & Qouiy6);
assign Qouiy6 = (Wtuiy6 & Kzqiy6);
assign Wtuiy6 = (Buihw6 & Offhw6);
assign Offhw6 = (!Zec7z6[27]);
assign Hftov6 = (Jgtov6 & Ctnov6);
assign Ctnov6 = (!Ovbdt6);
assign Ovbdt6 = (Zec7z6[16] & Otiiy6);
assign Jgtov6 = (!Uqd7z6[17]);
assign Uqd7z6[17] = (Zec7z6[17] & Otiiy6);
assign Zofhw6 = (!Cvmiy6);
assign Kjmiy6 = (~(Mqiiy6 & Zec7z6[8]));
assign Snriy6 = (A8jiy6 & W6u6x6);
assign W6u6x6 = (!M7mov6);
assign M7mov6 = (~(Euuiy6 & Muuiy6));
assign Muuiy6 = (~(Uuuiy6 | L9cdt6));
assign Uuuiy6 = (Cvuiy6 & Kvuiy6);
assign Kvuiy6 = (~(A3ddt6 & Svuiy6));
assign Svuiy6 = (~(Awuiy6 & Iwuiy6));
assign Iwuiy6 = (~(Yiaov6 & Qwuiy6));
assign Qwuiy6 = (Ywuiy6 | Gxuiy6);
assign Awuiy6 = (~(Fjaov6 & Oxuiy6));
assign Oxuiy6 = (~(Wxuiy6 & Eyuiy6));
assign Eyuiy6 = (Kbriy6 | Ghiiy6);
assign Cvuiy6 = (Myuiy6 | IFLUSH);
assign Euuiy6 = (K3jnv6 & Ldo7v6);
assign A8jiy6 = (~(Cta7x6 | Tjhov6));
assign Tjhov6 = (!Lybdt6);
assign Cta7x6 = (!Mjhov6);
assign Mjhov6 = (D6mov6 & Y6mov6);
assign Y6mov6 = (~(Gxuiy6 | Uyuiy6));
assign Uyuiy6 = (~(Wxuiy6 | Ywuiy6));
assign Wxuiy6 = (Kbriy6 | Ohiiy6);
assign Ohiiy6 = (Czuiy6 & Kzuiy6);
assign Kzuiy6 = (~(Gcd7z6[3] & L9d7z6[4]));
assign Czuiy6 = (Szuiy6 & A0viy6);
assign A0viy6 = (~(Gcd7z6[5] & L9d7z6[0]));
assign Szuiy6 = (~(Gcd7z6[1] & L9d7z6[2]));
assign D6mov6 = (~(Ywuiy6 | I0viy6));
assign I0viy6 = (Q0viy6 & Otiiy6);
assign Q0viy6 = (~(Gxuiy6 | Ghiiy6));
assign Ghiiy6 = (Y0viy6 & G1viy6);
assign G1viy6 = (~(Gcd7z6[1] & L9d7z6[3]));
assign Y0viy6 = (O1viy6 & W1viy6);
assign W1viy6 = (~(Gcd7z6[3] & L9d7z6[5]));
assign O1viy6 = (~(Gcd7z6[5] & L9d7z6[1]));
assign Gxuiy6 = (~(E2viy6 & M2viy6));
assign M2viy6 = (~(L9d7z6[2] & U2viy6));
assign E2viy6 = (C3viy6 & K3viy6);
assign K3viy6 = (~(L9d7z6[0] & S3viy6));
assign C3viy6 = (~(L9d7z6[4] & A4viy6));
assign Ywuiy6 = (~(I4viy6 & Q4viy6));
assign Q4viy6 = (~(L9d7z6[3] & U2viy6));
assign U2viy6 = (Gcd7z6[2] | Gcd7z6[3]);
assign I4viy6 = (Y4viy6 & G5viy6);
assign G5viy6 = (~(L9d7z6[1] & S3viy6));
assign S3viy6 = (Gcd7z6[0] | Gcd7z6[1]);
assign Y4viy6 = (~(L9d7z6[5] & A4viy6));
assign A4viy6 = (Gcd7z6[4] | Gcd7z6[5]);
assign Umriy6 = (~(Nvvnv6 & O5viy6));
assign O5viy6 = (~(Txinv6 & W5viy6));
assign W5viy6 = (~(E6viy6 & Yl2et6));
assign E6viy6 = (~(Szc7x6 | Ii9ov6));
assign Txinv6 = (~(M6viy6 | Z6xxx6));
assign Z6xxx6 = (Vgwxx6 | Lhwxx6);
assign Lhwxx6 = (Kihhw6 & U6viy6);
assign U6viy6 = (~(Ajphw6 & J0q6x6));
assign J0q6x6 = (!V1c7z6[12]);
assign Vgwxx6 = (C7viy6 & Rihhw6);
assign C7viy6 = (~(Yihhw6 & K7viy6));
assign K7viy6 = (~(V1c7z6[14] & Ajphw6));
assign M6viy6 = (~(F8xxx6 & S7viy6));
assign S7viy6 = (!R6xxx6);
assign R6xxx6 = (A8viy6 & V1c7z6[15]);
assign A8viy6 = (Szc7x6 & Ajphw6);
assign Szc7x6 = (Rihhw6 | Hir8v6);
assign F8xxx6 = (!Dhwxx6);
assign Dhwxx6 = (B6xxx6 | L5xxx6);
assign L5xxx6 = (I8viy6 & V1c7z6[11]);
assign I8viy6 = (Q8viy6 & Ajphw6);
assign Q8viy6 = (~(Ikmiy6 & Y8viy6));
assign Y8viy6 = (~(Hir8v6 & Nnr8v6));
assign B6xxx6 = (~(G9viy6 & Xjwxx6));
assign Xjwxx6 = (O9viy6 & W9viy6);
assign W9viy6 = (N4wxx6 & Vkwxx6);
assign Vkwxx6 = (!P3wxx6);
assign P3wxx6 = (Eaviy6 & Ycniy6);
assign Eaviy6 = (Maviy6 & Uaviy6);
assign Uaviy6 = (~(Ajphw6 & G8phw6));
assign G8phw6 = (!V1c7z6[3]);
assign Maviy6 = (~(Pxmov6 & Xumov6));
assign N4wxx6 = (~(Cbviy6 & Xkr8v6));
assign Cbviy6 = (Ycniy6 & Kbviy6);
assign Kbviy6 = (~(Ajphw6 & N7s6x6));
assign N7s6x6 = (!V1c7z6[2]);
assign O9viy6 = (F4wxx6 & X3wxx6);
assign X3wxx6 = (~(G1niy6 | Pzwxx6));
assign Pzwxx6 = (Sbviy6 & V1c7z6[4]);
assign Sbviy6 = (Ycniy6 & Ajphw6);
assign G1niy6 = (!Hzwxx6);
assign Hzwxx6 = (~(Acviy6 & V1c7z6[5]));
assign Acviy6 = (Icviy6 & Qcviy6);
assign Qcviy6 = (~(Y8niy6 & Pxmov6));
assign F4wxx6 = (Bywxx6 & Txwxx6);
assign Txwxx6 = (!Qgniy6);
assign Qgniy6 = (Ycviy6 & Qtvnv6);
assign Qtvnv6 = (!Yl2et6);
assign Ycviy6 = (~(J6jnv6 & Ajphw6));
assign J6jnv6 = (!V1c7z6[0]);
assign Bywxx6 = (!Ohniy6);
assign Ohniy6 = (Gdviy6 & Odviy6);
assign Odviy6 = (~(Ajphw6 & C6jnv6));
assign C6jnv6 = (!V1c7z6[1]);
assign G9viy6 = (X7xxx6 & Wdviy6);
assign Wdviy6 = (!Tlwxx6);
assign Tlwxx6 = (~(Fwwxx6 & Nwwxx6));
assign Nwwxx6 = (~(Eeviy6 & V1c7z6[7]));
assign Eeviy6 = (Meviy6 & Ueviy6);
assign Ueviy6 = (~(Cfviy6 & Y8niy6));
assign Cfviy6 = (Pxmov6 & Xumov6);
assign Fwwxx6 = (~(V1c7z6[6] & Icviy6));
assign Icviy6 = (Meviy6 & Kfviy6);
assign Kfviy6 = (~(Y8niy6 & Xumov6));
assign X7xxx6 = (Sfviy6 & Ziwxx6);
assign Ziwxx6 = (!Gtmiy6);
assign Gtmiy6 = (Meviy6 & V1c7z6[8]);
assign Meviy6 = (Dqr8v6 & Ajphw6);
assign Sfviy6 = (Hjwxx6 & Agviy6);
assign Agviy6 = (!Pjwxx6);
assign Pjwxx6 = (Igviy6 & V1c7z6[10]);
assign Igviy6 = (Qgviy6 & Ajphw6);
assign Hjwxx6 = (!Dxwxx6);
assign Dxwxx6 = (Ygviy6 & V1c7z6[9]);
assign Ygviy6 = (Mumiy6 & Ajphw6);
assign Mumiy6 = (Qgviy6 & Ghviy6);
assign Ghviy6 = (~(Pxmov6 & Xlaov6));
assign Qgviy6 = (!Ikmiy6);
assign Ikmiy6 = (~(Kihhw6 & Ohviy6));
assign Ohviy6 = (~(Xumov6 & Xlaov6));
assign Qkriy6 = (~(Whviy6 & Eiviy6));
assign Eiviy6 = (Mlfov6 & Gvvnv6);
assign Mlfov6 = (!Yfadt6);
assign Whviy6 = (Ytlnv6 & Fulnv6);
assign Y0oiy6 = (~(Miviy6 | A8mov6));
assign A8mov6 = (Tlmov6 & Uiviy6);
assign Uiviy6 = (~(Cjviy6 & Sosiw6));
assign Sosiw6 = (!Wkb7z6[2]);
assign Miviy6 = (Xsddt6 & Qg2nv6);
assign Kzniy6 = (S6cdt6 & S2onv6);
assign S2onv6 = (~(Nhonv6 & Kjviy6));
assign Kjviy6 = (Vglhw6 | Atmov6);
assign Atmov6 = (Fulnv6 & Mahiy6);
assign Hwr7x6 = (~(Teliw6 | S1wnv6));
assign Teliw6 = (!Kkmhw6);
assign Kkmhw6 = (~(Tlmov6 & Sjviy6));
assign Sjviy6 = (Dqnov6 | Y2piw6);
assign Y2piw6 = (!Dxvnv6);
assign Dxvnv6 = (S1wnv6 | Q0wnv6);
assign S1wnv6 = (Akviy6 & Tlmov6);
assign Akviy6 = (Ikviy6 & Xsinv6);
assign Ikviy6 = (~(Qkviy6 & Cjviy6));
assign Cjviy6 = (K6mov6 & Vmsiw6);
assign Vmsiw6 = (Ykviy6 & Glviy6);
assign Ykviy6 = (Olviy6 & Wlviy6);
assign Olviy6 = (M697z6 & Emviy6);
assign K6mov6 = (~(Tlb7z6[0] | Wkb7z6[0]));
assign Qkviy6 = (Mmviy6 & Jnsiw6);
assign Jnsiw6 = (!Ffadt6);
assign Mmviy6 = (~(Umviy6 & V6l8v6));
assign V6l8v6 = (Cnviy6 & K9d7x6);
assign Cnviy6 = (~(Knviy6 & Snviy6));
assign Snviy6 = (Qolov6 ? Ioviy6 : Aoviy6);
assign Qolov6 = (Qoviy6 & Yoviy6);
assign Yoviy6 = (~(D9d7x6 & E3c7z6[3]));
assign Qoviy6 = (~(D6c7z6[3] & Cubdt6));
assign Ioviy6 = (Ad9iw6 & Gpviy6);
assign Gpviy6 = (~(Umviy6 & Ea2nv6));
assign Ad9iw6 = (Opviy6 & Wpviy6);
assign Wpviy6 = (~(D9d7x6 & E3c7z6[2]));
assign Opviy6 = (~(D6c7z6[2] & Cubdt6));
assign Aoviy6 = (Ea2nv6 | Aqadt6);
assign Knviy6 = (E6d7x6 & C5d7x6);
assign C5d7x6 = (~(Eqviy6 & Mqviy6));
assign Mqviy6 = (~(D9d7x6 & E3c7z6[0]));
assign Eqviy6 = (~(Cubdt6 & D6c7z6[0]));
assign E6d7x6 = (Uqviy6 & Crviy6);
assign Crviy6 = (~(D9d7x6 & E3c7z6[1]));
assign Uqviy6 = (~(D6c7z6[1] & Cubdt6));
assign Umviy6 = (~(Ev2nv6 | Dxgov6));
assign Dqnov6 = (Krviy6 & Yfadt6);
assign Krviy6 = (Srviy6 & O5a7z6);
assign Kd2nv6 = (Asviy6 & Isviy6);
assign Isviy6 = (~(Qsviy6 | Lafov6));
assign Lafov6 = (Ysviy6 & Y5o7x6);
assign Y5o7x6 = (Gtviy6 & Otviy6);
assign Otviy6 = (~(Wtviy6 & Euviy6));
assign Euviy6 = (~(Y94iw6 | W22ft6));
assign Y94iw6 = (!Lhmov6);
assign Wtviy6 = (~(Muviy6 | Uuviy6));
assign Uuviy6 = (Po4ft6 & Mdo7x6);
assign Muviy6 = (R25yx6 ? I7p7z6[0] : K5o7x6);
assign R25yx6 = (!D5o7x6);
assign K5o7x6 = (I7p7z6[1] | P35yx6);
assign Gtviy6 = (~(Cvviy6 | Cx5ov6));
assign Cx5ov6 = (Cq2ft6 & Kvviy6);
assign Kvviy6 = (~(Svviy6 & Awviy6));
assign Awviy6 = (~(Iwviy6 & Tv5ov6));
assign Tv5ov6 = (!Bup7z6[1]);
assign Svviy6 = (~(Qwviy6 & Aw5ov6));
assign Aw5ov6 = (!Wrp7z6[1]);
assign Cvviy6 = (Ywviy6 & Gxviy6);
assign Gxviy6 = (~(Po4ft6 & Mdo7x6));
assign Ywviy6 = (~(Oxviy6 & Fs4ft6));
assign Oxviy6 = (Wxviy6 & Eyviy6);
assign Eyviy6 = (~(Myviy6 & Uyviy6));
assign Myviy6 = (~(I7p7z6[0] | I7p7z6[1]));
assign Wxviy6 = (Czviy6 | W22ft6);
assign Czviy6 = (Gjdiw6 & Kzviy6);
assign Kzviy6 = (~(Szviy6 & A0wiy6));
assign A0wiy6 = (D5o7x6 ^ I7p7z6[0]);
assign D5o7x6 = (~(I0wiy6 & I7p7z6[3]));
assign I0wiy6 = (I7p7z6[2] & HTMDHBURST[0]);
assign Szviy6 = (~(Lhmov6 | P35yx6));
assign P35yx6 = (Uyviy6 & HTMDHBURST[0]);
assign Uyviy6 = (~(I7p7z6[2] | I7p7z6[3]));
assign Ysviy6 = (~(L9o7x6 | I7p7z6[3]));
assign L9o7x6 = (!I7p7z6[2]);
assign Qsviy6 = (X9fov6 | Eafov6);
assign Eafov6 = (Q0wiy6 & Hmp7z6[2]);
assign Q0wiy6 = (~(N2a8x6 | Hmp7z6[3]));
assign N2a8x6 = (Y0wiy6 & G1wiy6);
assign G1wiy6 = (~(O1wiy6 & J95ft6));
assign O1wiy6 = (Mdo7x6 & B4fiw6);
assign Y0wiy6 = (~(W1wiy6 & E2wiy6));
assign E2wiy6 = (M2wiy6 & U2wiy6);
assign U2wiy6 = (~(C3wiy6 & Veo7x6));
assign Veo7x6 = (~(K3wiy6 & HTMDHBURST[0]));
assign K3wiy6 = (~(Hmp7z6[2] | Hmp7z6[3]));
assign C3wiy6 = (Lhmov6 ? Jfo7x6 : Cfo7x6);
assign Jfo7x6 = (!S3wiy6);
assign S3wiy6 = (By4yx6 ? Hmp7z6[0] : Hmp7z6[1]);
assign Cfo7x6 = (~(By4yx6 ^ Hmp7z6[0]));
assign By4yx6 = (!Mko7x6);
assign Mko7x6 = (~(A4wiy6 & Hmp7z6[3]));
assign A4wiy6 = (Hmp7z6[2] & HTMDHBURST[0]);
assign M2wiy6 = (I4wiy6 & B4fiw6);
assign B4fiw6 = (~(Cq2ft6 & Q4wiy6));
assign Q4wiy6 = (~(Y4wiy6 & G5wiy6));
assign G5wiy6 = (~(Bup7z6[1] & Iwviy6));
assign Iwviy6 = (!Bup7z6[0]);
assign Y4wiy6 = (~(Wrp7z6[1] & Qwviy6));
assign Qwviy6 = (!Wrp7z6[0]);
assign I4wiy6 = (~(O5wiy6 & Zy4yx6));
assign Zy4yx6 = (!Hmp7z6[0]);
assign O5wiy6 = (~(Hmp7z6[1] | Hmp7z6[2]));
assign W1wiy6 = (Zc5ft6 & Gjdiw6);
assign X9fov6 = (W5wiy6 & Hyp7z6[2]);
assign W5wiy6 = (V0fiw6 & E6wiy6);
assign V0fiw6 = (~(M6wiy6 & U6wiy6));
assign U6wiy6 = (~(C7wiy6 & K7wiy6));
assign K7wiy6 = (S7wiy6 & Gjdiw6);
assign S7wiy6 = (~(Lx6ov6 | Cq2ft6));
assign Lx6ov6 = (A8wiy6 & I8wiy6);
assign A8wiy6 = (Q1fiw6 & Vz98x6);
assign C7wiy6 = (Q8wiy6 & Q35ft6);
assign Q8wiy6 = (!Y8wiy6);
assign Y8wiy6 = (Lhmov6 ? V18ov6 : O18ov6);
assign V18ov6 = (!Dco7x6);
assign Dco7x6 = (G9wiy6 & O9wiy6);
assign O9wiy6 = (~(E2fiw6 & I8wiy6));
assign I8wiy6 = (!Hyp7z6[0]);
assign G9wiy6 = (~(X1fiw6 & Q1fiw6));
assign Q1fiw6 = (!Hyp7z6[1]);
assign O18ov6 = (Hyp7z6[0] ? E2fiw6 : X1fiw6);
assign X1fiw6 = (~(E2fiw6 | D15yx6));
assign D15yx6 = (W9wiy6 & HTMDHBURST[0]);
assign W9wiy6 = (Vz98x6 & E6wiy6);
assign E6wiy6 = (!Hyp7z6[3]);
assign Vz98x6 = (!Hyp7z6[2]);
assign E2fiw6 = (Eawiy6 & Hyp7z6[3]);
assign Eawiy6 = (Hyp7z6[2] & HTMDHBURST[0]);
assign M6wiy6 = (Mawiy6 & Xch7v6);
assign Mawiy6 = (~(A05ft6 & Mdo7x6));
assign Asviy6 = (~(Sn8iw6 | L99ov6));
assign L99ov6 = (Uawiy6 & Sgp7z6[2]);
assign Uawiy6 = (~(Wxeiw6 | Sgp7z6[3]));
assign Wxeiw6 = (Cbwiy6 & Kbwiy6);
assign Kbwiy6 = (~(Sbwiy6 & Hk5ft6));
assign Sbwiy6 = (Mdo7x6 & D5fiw6);
assign Mdo7x6 = (Ke2ft6 & Cpsnv6);
assign Cbwiy6 = (~(Acwiy6 & Icwiy6));
assign Icwiy6 = (Qcwiy6 & Ycwiy6);
assign Ycwiy6 = (~(Gdwiy6 & F6fiw6));
assign F6fiw6 = (~(Odwiy6 & HTMDHBURST[0]));
assign Odwiy6 = (~(Sgp7z6[2] | Sgp7z6[3]));
assign Gdwiy6 = (Lhmov6 ? T6fiw6 : M6fiw6);
assign T6fiw6 = (!Wdwiy6);
assign Wdwiy6 = (Tzeiw6 ? Sgp7z6[0] : Sgp7z6[1]);
assign M6fiw6 = (~(Tzeiw6 ^ Sgp7z6[0]));
assign Tzeiw6 = (Eewiy6 & Sgp7z6[3]);
assign Eewiy6 = (Sgp7z6[2] & HTMDHBURST[0]);
assign Qcwiy6 = (Mewiy6 & D5fiw6);
assign D5fiw6 = (~(Cq2ft6 & Uewiy6));
assign Uewiy6 = (~(Cfwiy6 & Kfwiy6));
assign Kfwiy6 = (~(Bup7z6[0] & Bup7z6[1]));
assign Cfwiy6 = (~(Wrp7z6[0] & Wrp7z6[1]));
assign Mewiy6 = (Sfwiy6 | Sgp7z6[0]);
assign Sfwiy6 = (Sgp7z6[1] | Sgp7z6[2]);
assign Acwiy6 = (Xn5ft6 & Gjdiw6);
assign Gjdiw6 = (~(Shmov6 | Nhonv6));
assign Shmov6 = (!Vfmov6);
assign Vfmov6 = (Gr2et6 & Vb4iw6);
assign Gr2et6 = (O5a7z6 & Aeonv6);
assign Aeonv6 = (~(Wcmov6 & Agwiy6));
assign Agwiy6 = (~(Igwiy6 & Qgwiy6));
assign Igwiy6 = (~(Ygwiy6 & Ghwiy6));
assign Ghwiy6 = (~(Ohwiy6 & HREADYD));
assign Ohwiy6 = (Whwiy6 & Ibonv6);
assign Ygwiy6 = (Eiwiy6 & Miwiy6);
assign Miwiy6 = (~(Uiwiy6 & Gyjiw6));
assign Uiwiy6 = (Cjwiy6 & Vd2iw6);
assign Eiwiy6 = (~(Kjwiy6 & Sjwiy6));
assign Kjwiy6 = (HREADYS & Uaonv6);
assign Sn8iw6 = (Akwiy6 | EDBGRQ);
assign Akwiy6 = (~(Ikwiy6 & Edh7v6));
assign Ikwiy6 = (!Mq97z6);
assign Q7hov6 = (!V9m7x6);
assign V9m7x6 = (~(Qkwiy6 & Ykwiy6));
assign Ykwiy6 = (~(Glwiy6 | Yd2nv6));
assign Yd2nv6 = (Olwiy6 & Wlwiy6);
assign Wlwiy6 = (~(Emwiy6 & Mmwiy6));
assign Mmwiy6 = (~(Umwiy6 & Cnwiy6));
assign Olwiy6 = (Knwiy6 & Izs7x6);
assign Izs7x6 = (~(Ea2nv6 & Jm98x6));
assign Ea2nv6 = (!Snwiy6);
assign Knwiy6 = (~(Y0t7x6 & Aowiy6));
assign Aowiy6 = (~(Iowiy6 & Pahov6));
assign Iowiy6 = (Umwiy6 & Cnwiy6);
assign Cnwiy6 = (~(Qowiy6 & Yowiy6));
assign Yowiy6 = (Gpwiy6 & Cehov6);
assign Gpwiy6 = (~(Jehov6 & B6t7x6));
assign Qowiy6 = (Rwl8v6 & N5t7x6);
assign Umwiy6 = (B6t7x6 | Jehov6);
assign Glwiy6 = (Fe2nv6 | Nmadt6);
assign Fe2nv6 = (!Amg7x6);
assign Qkwiy6 = (E1cet6 & Te2nv6);
assign Te2nv6 = (Etinv6 & Opwiy6);
assign Opwiy6 = (~(Wpwiy6 & Eqwiy6));
assign Wpwiy6 = (Mqwiy6 & Uqwiy6);
assign Uqwiy6 = (~(Crwiy6 & Emwiy6));
assign Emwiy6 = (!Pahov6);
assign Crwiy6 = (~(Krwiy6 & Ldr7x6));
assign Mqwiy6 = (Ldr7x6 | Krwiy6);
assign Krwiy6 = (Srwiy6 & Aswiy6);
assign Aswiy6 = (~(Iswiy6 & Qswiy6));
assign Qswiy6 = (CURRPRI[5] & Cehov6);
assign Cehov6 = (!Nbj7z6[0]);
assign Iswiy6 = (Rwl8v6 & Yswiy6);
assign Yswiy6 = (~(Jehov6 & Bfr7x6));
assign Srwiy6 = (~(Ger7x6 & Adhov6));
assign Adhov6 = (!Jehov6);
assign Awniy6 = (~(Lh18x6 & Ykliy6));
assign Sln7v6 = (W3e7v6 ^ Gtwiy6);
assign Gtwiy6 = (Vuf7v6 & Twhiw6);
assign Lln7v6 = (Kygnv6 ? Otwiy6 : Imh7v6);
assign Otwiy6 = (!W597z6);
assign Eln7v6 = (Kygnv6 ? We6ft6 : Wtwiy6);
assign Wtwiy6 = (Ci6ft6 & Euwiy6);
assign Euwiy6 = (~(W597z6 & Og6ft6));
assign Xkn7v6 = (Kygnv6 ? Qb6ft6 : Muwiy6);
assign Muwiy6 = (Uuwiy6 & We6ft6);
assign Uuwiy6 = (Og6ft6 & Ci6ft6);
assign Qkn7v6 = (P7fyx6 ? Nks7z6[1] : Iuvmz6[5]);
assign Jkn7v6 = (P7fyx6 ? Nks7z6[2] : Iuvmz6[6]);
assign Ckn7v6 = (P7fyx6 ? Nks7z6[3] : Iuvmz6[7]);
assign Vjn7v6 = (P7fyx6 ? Nks7z6[4] : Iuvmz6[8]);
assign Ojn7v6 = (P7fyx6 ? Nks7z6[0] : Iuvmz6[4]);
assign P7fyx6 = (V4byx6 & Cvwiy6);
assign Cvwiy6 = (~(Kvwiy6 & Eifnv6));
assign Kvwiy6 = (~(E46ft6 | Ur37v6));
assign V4byx6 = (!Fo4yx6);
assign Fo4yx6 = (~(Svwiy6 & Awwiy6));
assign Awwiy6 = (Iwwiy6 & Qwwiy6);
assign Qwwiy6 = (~(Ywwiy6 & Jafyx6));
assign Jafyx6 = (O2wmz6[0] ^ Z6fyx6);
assign Z6fyx6 = (!Y4wmz6[0]);
assign Ywwiy6 = (Gxwiy6 & X7fyx6);
assign X7fyx6 = (Oxwiy6 | Wxwiy6);
assign Wxwiy6 = (~(Eywiy6 & Mywiy6));
assign Mywiy6 = (~(Iuvmz6[5] & Yo37v6));
assign Eywiy6 = (~(Iuvmz6[7] & Uywiy6));
assign Oxwiy6 = (~(Czwiy6 & Kzwiy6));
assign Kzwiy6 = (~(Iuvmz6[6] & Szwiy6));
assign Czwiy6 = (~(A0xiy6 | Iuvmz6[4]));
assign A0xiy6 = (Iuvmz6[8] & I0xiy6);
assign Gxwiy6 = (~(Y4wmz6[1] ^ L56yx6));
assign L56yx6 = (!O2wmz6[1]);
assign Iwwiy6 = (Q0xiy6 & Y0xiy6);
assign Y0xiy6 = (~(G1xiy6 & T1gyx6));
assign T1gyx6 = (A3xmz6[0] ^ H76yx6);
assign H76yx6 = (!K5xmz6[0]);
assign G1xiy6 = (O1xiy6 & Zifyx6);
assign Zifyx6 = (~(W1xiy6 & E2xiy6));
assign E2xiy6 = (M2xiy6 & U2xiy6);
assign U2xiy6 = (~(Iuvmz6[5] & Szwiy6));
assign M2xiy6 = (~(C3xiy6 | Iuvmz6[8]));
assign C3xiy6 = (Iuvmz6[7] & I0xiy6);
assign W1xiy6 = (K3xiy6 & S3xiy6);
assign S3xiy6 = (~(Iuvmz6[6] & Uywiy6));
assign K3xiy6 = (~(Iuvmz6[4] & Yo37v6));
assign O1xiy6 = (~(K5xmz6[1] ^ Zm3yx6));
assign Zm3yx6 = (!A3xmz6[1]);
assign Q0xiy6 = (~(A4xiy6 & Pffyx6));
assign Pffyx6 = (Ukwmz6[0] ^ Vc6yx6);
assign Vc6yx6 = (!Enwmz6[0]);
assign A4xiy6 = (I4xiy6 & Ldfyx6);
assign Ldfyx6 = (~(Q4xiy6 & Y4xiy6));
assign Y4xiy6 = (G5xiy6 & O5xiy6);
assign O5xiy6 = (~(Iuvmz6[5] & I0xiy6));
assign G5xiy6 = (~(W5xiy6 | Iuvmz6[6]));
assign W5xiy6 = (Iuvmz6[8] & Szwiy6);
assign Q4xiy6 = (E6xiy6 & M6xiy6);
assign M6xiy6 = (~(Iuvmz6[7] & Yo37v6));
assign E6xiy6 = (~(Iuvmz6[4] & Uywiy6));
assign I4xiy6 = (~(Enwmz6[1] ^ Ze6yx6));
assign Ze6yx6 = (!Ukwmz6[1]);
assign Svwiy6 = (U6xiy6 & C7xiy6);
assign C7xiy6 = (~(K7xiy6 & Vcfyx6));
assign Vcfyx6 = (Rbwmz6[0] ^ Vg6yx6);
assign Vg6yx6 = (!Bewmz6[0]);
assign K7xiy6 = (S7xiy6 & Zafyx6);
assign Zafyx6 = (~(A8xiy6 & I8xiy6));
assign I8xiy6 = (Q8xiy6 & Y8xiy6);
assign Y8xiy6 = (~(Iuvmz6[4] & I0xiy6));
assign Q8xiy6 = (~(G9xiy6 | Iuvmz6[5]));
assign G9xiy6 = (Szwiy6 & Iuvmz6[7]);
assign A8xiy6 = (O9xiy6 & W9xiy6);
assign W9xiy6 = (~(Iuvmz6[8] & Uywiy6));
assign O9xiy6 = (~(Iuvmz6[6] & Yo37v6));
assign S7xiy6 = (~(Bewmz6[1] ^ Hj6yx6));
assign Hj6yx6 = (!Rbwmz6[1]);
assign U6xiy6 = (~(Eaxiy6 & Jifyx6));
assign Jifyx6 = (Xtwmz6[0] ^ V86yx6);
assign V86yx6 = (!Hwwmz6[0]);
assign Eaxiy6 = (Maxiy6 & Fgfyx6);
assign Fgfyx6 = (~(Uaxiy6 & Cbxiy6));
assign Cbxiy6 = (Kbxiy6 & Sbxiy6);
assign Sbxiy6 = (~(Iuvmz6[4] & Szwiy6));
assign Szwiy6 = (Uywiy6 & Acxiy6);
assign Acxiy6 = (M6s7z6[0] | Yo37v6);
assign Kbxiy6 = (~(Icxiy6 | Iuvmz6[7]));
assign Icxiy6 = (Iuvmz6[6] & I0xiy6);
assign I0xiy6 = (Uywiy6 | M6s7z6[0]);
assign M6s7z6[0] = (~(Qcxiy6 & Ycxiy6));
assign Ycxiy6 = (Gdxiy6 & Odxiy6);
assign Odxiy6 = (~(Wdxiy6 & X9s7z6[0]));
assign Wdxiy6 = (L17yx6 & Eexiy6);
assign Eexiy6 = (!X9s7z6[1]);
assign Gdxiy6 = (~(H77yx6 | Xz7yx6));
assign Xz7yx6 = (Ju5yx6 & Hnayx6);
assign H77yx6 = (~(Mexiy6 | Uexiy6));
assign Mexiy6 = (!J27yx6);
assign Qcxiy6 = (Cfxiy6 & Kfxiy6);
assign Kfxiy6 = (~(Rmayx6 & Rq9yx6));
assign Cfxiy6 = (Sfxiy6 & Agxiy6);
assign Agxiy6 = (~(Cu5ft6 & Vkfyx6));
assign Vkfyx6 = (!L1dyx6);
assign Sfxiy6 = (~(Be7yx6 & Igxiy6));
assign Uaxiy6 = (Qgxiy6 & Ygxiy6);
assign Ygxiy6 = (~(Iuvmz6[8] & Yo37v6));
assign Qgxiy6 = (~(Iuvmz6[5] & Uywiy6));
assign Uywiy6 = (M6s7z6[1] | Yo37v6);
assign Yo37v6 = (~(Ghxiy6 & Ohxiy6));
assign Ohxiy6 = (~(Jmayx6 | R27yx6));
assign R27yx6 = (~(L1dyx6 | Cu5ft6));
assign L1dyx6 = (~(Ra5yx6 & Hnayx6));
assign Ra5yx6 = (!Xnayx6);
assign Xnayx6 = (~(Whxiy6 & Eixiy6));
assign Whxiy6 = (~(F85yx6 | Ju5yx6));
assign Jmayx6 = (~(Dt8yx6 | Xy5ft6));
assign Dt8yx6 = (!N47yx6);
assign Ghxiy6 = (Mixiy6 & Uixiy6);
assign Uixiy6 = (~(X9s7z6[0] & Tp9yx6));
assign Mixiy6 = (~(Xcr7z6[1] & Rmayx6));
assign Rmayx6 = (~(Dd7yx6 | Xcr7z6[0]));
assign M6s7z6[1] = (~(Cjxiy6 & Kjxiy6));
assign Kjxiy6 = (Nw7yx6 & Sjxiy6);
assign Sjxiy6 = (~(Akxiy6 & Xcr7z6[0]));
assign Akxiy6 = (P37yx6 & Rq9yx6);
assign Rq9yx6 = (!Xcr7z6[1]);
assign P37yx6 = (!Dd7yx6);
assign Dd7yx6 = (~(Ikxiy6 & Ixr7z6[1]));
assign Ikxiy6 = (Hnayx6 & T1byx6);
assign T1byx6 = (!Xwadt6);
assign Nw7yx6 = (Qkxiy6 & Tt8yx6);
assign Tt8yx6 = (!V47yx6);
assign V47yx6 = (F85yx6 & Hnayx6);
assign F85yx6 = (Ykxiy6 & Uur7z6[1]);
assign Ykxiy6 = (Eixiy6 & Ri5yx6);
assign Ri5yx6 = (!Ju5yx6);
assign Ju5yx6 = (C4s7z6[1] & Eixiy6);
assign Qkxiy6 = (~(Xy5ft6 & N47yx6));
assign N47yx6 = (Xwadt6 & Hnayx6);
assign Hnayx6 = (Glxiy6 & D5byx6);
assign Glxiy6 = (No4yx6 & Ld7yx6);
assign Cjxiy6 = (Olxiy6 & Wlxiy6);
assign Wlxiy6 = (~(Tp9yx6 & Emxiy6));
assign Emxiy6 = (!X9s7z6[0]);
assign Tp9yx6 = (X9s7z6[1] & L17yx6);
assign L17yx6 = (~(No4yx6 | Ur37v6));
assign No4yx6 = (!I96ft6);
assign Olxiy6 = (~(Be7yx6 & L94yx6));
assign Be7yx6 = (J27yx6 & V0dyx6);
assign V0dyx6 = (~(Mmxiy6 & Umxiy6));
assign Umxiy6 = (F84yx6 & Cnxiy6);
assign Cnxiy6 = (~(Vs27v6 | Nu27v6));
assign F84yx6 = (~(P7s7z6[13] | P7s7z6[14]));
assign Mmxiy6 = (Knxiy6 & D94yx6);
assign D94yx6 = (~(P7s7z6[11] | P7s7z6[12]));
assign Knxiy6 = (Igxiy6 & Snxiy6);
assign Snxiy6 = (~(Aoxiy6 & P7s7z6[9]));
assign Aoxiy6 = (P7s7z6[8] & P7s7z6[10]);
assign Igxiy6 = (!L94yx6);
assign L94yx6 = (~(Ioxiy6 & Qoxiy6));
assign Qoxiy6 = (Yoxiy6 & N44yx6);
assign N44yx6 = (~(P7s7z6[21] | P7s7z6[22]));
assign Yoxiy6 = (~(P7s7z6[19] | P7s7z6[20]));
assign Ioxiy6 = (Gpxiy6 & Opxiy6);
assign Opxiy6 = (~(P7s7z6[17] | P7s7z6[18]));
assign Gpxiy6 = (Uexiy6 & Z64yx6);
assign Z64yx6 = (!P7s7z6[16]);
assign Uexiy6 = (Wpxiy6 & Eqxiy6);
assign Eqxiy6 = (Mqxiy6 & Uqxiy6);
assign Uqxiy6 = (~(P7s7z6[29] | P7s7z6[30]));
assign Mqxiy6 = (~(P7s7z6[27] | P7s7z6[28]));
assign Wpxiy6 = (Crxiy6 & L54yx6);
assign L54yx6 = (!P7s7z6[24]);
assign Crxiy6 = (~(P7s7z6[25] | P7s7z6[26]));
assign J27yx6 = (Krxiy6 & E46ft6);
assign Krxiy6 = (Eifnv6 & Ld7yx6);
assign Ld7yx6 = (!Ur37v6);
assign Eifnv6 = (!Fho7v6);
assign Maxiy6 = (~(Hwwmz6[1] ^ Za6yx6));
assign Za6yx6 = (!Xtwmz6[1]);
assign Hjn7v6 = (Yfadt6 | Phhov6);
assign Phhov6 = (L8oov6 & Ouyiw6);
assign Ouyiw6 = (~(Srxiy6 & Asxiy6));
assign Asxiy6 = (~(Pj1ov6 & Isxiy6));
assign Isxiy6 = (Qsxiy6 | Szoiw6);
assign Szoiw6 = (!P51ov6);
assign P51ov6 = (~(X9mhw6 & Cgc7z6[2]));
assign X9mhw6 = (Ydmhw6 & V4jhw6);
assign Ydmhw6 = (~(Cgc7z6[1] | Cgc7z6[0]));
assign Qsxiy6 = (Gtxiy6 ? Ipnov6 : Ysxiy6);
assign Ysxiy6 = (C21ov6 & R537x6);
assign C21ov6 = (B51ov6 & V4jhw6);
assign Pj1ov6 = (!IFLUSH);
assign Srxiy6 = (~(Z1oov6 & Gtxiy6));
assign Gtxiy6 = (!Uicdt6);
assign Z1oov6 = (Otxiy6 & Cgc7z6[2]);
assign Otxiy6 = (Cgc7z6[1] & O4jhw6);
assign L8oov6 = (R537x6 & X0oov6);
assign X0oov6 = (!Rxnov6);
assign Rxnov6 = (B51ov6 & T3jhw6);
assign Ajn7v6 = (Euxiy6 ? Wtxiy6 : Ab57v6);
assign Euxiy6 = (Quthw6 & Npthw6);
assign Quthw6 = (Muxiy6 & Hixhw6);
assign Hixhw6 = (Oqwhw6 & Uzxmz6[2]);
assign Muxiy6 = (Uzxmz6[0] & Uzxmz6[1]);
assign Wtxiy6 = (~(Uuxiy6 & Cvxiy6));
assign Cvxiy6 = (~(Dnxhw6 & Ds57v6));
assign Uuxiy6 = (~(Kvxiy6 | Eothw6));
assign Eothw6 = (Dnxhw6 & Zhthw6);
assign Zhthw6 = (!Yn57v6);
assign Dnxhw6 = (~(Kp57v6 | Cl57v6));
assign Kvxiy6 = (Svxiy6 & Qazhw6);
assign Qazhw6 = (!Lc57v6);
assign Svxiy6 = (Dfrhw6 | Awxiy6);
assign Awxiy6 = (Iwxiy6 & Qwxiy6);
assign Qwxiy6 = (Ywxiy6 & Gxxiy6);
assign Gxxiy6 = (Oxxiy6 & Wxxiy6);
assign Wxxiy6 = (~(Njxmz6[9] | Ds57v6));
assign Oxxiy6 = (~(Njxmz6[7] | Njxmz6[8]));
assign Ywxiy6 = (~(Eyxiy6 | Njxmz6[4]));
assign Eyxiy6 = (Njxmz6[5] | Njxmz6[6]);
assign Iwxiy6 = (Myxiy6 & Uyxiy6);
assign Uyxiy6 = (Czxiy6 & Kzxiy6);
assign Kzxiy6 = (~(Njxmz6[2] | Njxmz6[3]));
assign Czxiy6 = (~(Njxmz6[11] | Njxmz6[1]));
assign Myxiy6 = (Szxiy6 & Kp57v6);
assign Szxiy6 = (~(Njxmz6[0] | Njxmz6[10]));
assign Dfrhw6 = (Hnzhw6 & Onzhw6);
assign Onzhw6 = (!R957v6);
assign Hnzhw6 = (!Ek47v6);
assign Tin7v6 = (A0yiy6 ? Aixmz6[4] : L5ymz6[7]);
assign Min7v6 = (A0yiy6 ? Aixmz6[5] : L5ymz6[8]);
assign Fin7v6 = (A0yiy6 ? Aixmz6[6] : L5ymz6[9]);
assign Yhn7v6 = (A0yiy6 ? Aixmz6[7] : L5ymz6[10]);
assign Rhn7v6 = (A0yiy6 ? Aixmz6[8] : L5ymz6[11]);
assign Khn7v6 = (A0yiy6 ? Aixmz6[9] : L5ymz6[12]);
assign Dhn7v6 = (A0yiy6 ? Aixmz6[10] : L5ymz6[13]);
assign Wgn7v6 = (A0yiy6 ? Aixmz6[11] : L5ymz6[14]);
assign Pgn7v6 = (A0yiy6 ? Aixmz6[22] : L5ymz6[25]);
assign Ign7v6 = (A0yiy6 ? Aixmz6[23] : L5ymz6[26]);
assign Bgn7v6 = (A0yiy6 ? Aixmz6[24] : L5ymz6[27]);
assign Ufn7v6 = (A0yiy6 ? Aixmz6[25] : L5ymz6[28]);
assign Nfn7v6 = (A0yiy6 ? Aixmz6[26] : L5ymz6[29]);
assign Gfn7v6 = (A0yiy6 ? Aixmz6[27] : L5ymz6[30]);
assign Zen7v6 = (A0yiy6 ? Aixmz6[28] : L5ymz6[31]);
assign Sen7v6 = (A0yiy6 ? Aixmz6[29] : L5ymz6[32]);
assign Len7v6 = (A0yiy6 ? Aixmz6[30] : L5ymz6[33]);
assign Een7v6 = (~(Sg1iw6 ^ Qs67z6));
assign Sg1iw6 = (I0yiy6 & Kh47v6);
assign I0yiy6 = (Gj47v6 & Q0yiy6);
assign Xdn7v6 = (T1zhw6 ? Y0yiy6 : Bmh7v6);
assign Qdn7v6 = (T1zhw6 ? Ye47v6 : Y0yiy6);
assign Y0yiy6 = (!Oh67z6);
assign Jdn7v6 = (T1zhw6 ? Up47v6 : G1yiy6);
assign G1yiy6 = (O1yiy6 & Ye47v6);
assign O1yiy6 = (Dbymz6[1] & E6qhw6);
assign Cdn7v6 = (~(W8qhw6 ^ Is67z6));
assign Vcn7v6 = (Xzvhw6 ? Fduhw6 : W1yiy6);
assign Xzvhw6 = (~(Ft1nv6 | Gq1nv6));
assign Ft1nv6 = (~(E2yiy6 & R9ymz6[2]));
assign E2yiy6 = (Nq1nv6 & K3whw6);
assign Nq1nv6 = (!R9ymz6[0]);
assign Fduhw6 = (~(P2whw6 & M2yiy6));
assign M2yiy6 = (R9qhw6 & U2yiy6);
assign U2yiy6 = (~(W8qhw6 & W6ymz6[0]));
assign W8qhw6 = (S367v6 & Ek47v6);
assign R9qhw6 = (Qs67z6 ^ Is67z6);
assign P2whw6 = (W6ymz6[1] & Co1nv6);
assign Ocn7v6 = (~(C3yiy6 | K9qhw6));
assign C3yiy6 = (~(Uu57v6 | K3yiy6));
assign K3yiy6 = (By1nv6 & W1yiy6);
assign Hcn7v6 = (T1zhw6 ? S3yiy6 : Ulh7v6);
assign Acn7v6 = (T1zhw6 ? Ee47v6 : S3yiy6);
assign S3yiy6 = (!Gh67z6);
assign Tbn7v6 = (I4yiy6 ? Fvzet6 : A4yiy6);
assign Mbn7v6 = (A0yiy6 ? Aixmz6[31] : L5ymz6[34]);
assign Fbn7v6 = (Q4yiy6 ? U3o7z6[31] : Fvb7z6[31]);
assign Yan7v6 = (Y4yiy6 ? U42nv6 : A0fet6);
assign Y4yiy6 = (Awbet6 & Zhg7x6);
assign Ran7v6 = (T8lov6 ? X4eet6 : Is5iw6);
assign Kan7v6 = (X27iw6 ? Fuadt6 : U47iw6);
assign X27iw6 = (~(G5yiy6 & R58iw6));
assign G5yiy6 = (Z4m7x6 & Bqi7z6[1]);
assign Dan7v6 = (O5yiy6 ? U42nv6 : Aqadt6);
assign W9n7v6 = (O5yiy6 ? W52nv6 : Esadt6);
assign P9n7v6 = (O5yiy6 ? P52nv6 : Dradt6);
assign O5yiy6 = (!W5yiy6);
assign I9n7v6 = (W5yiy6 ? O6cet6 : B52nv6);
assign W5yiy6 = (~(Zh18x6 & Z4m7x6));
assign B9n7v6 = (!E6yiy6);
assign E6yiy6 = (Wc0iw6 ? M6yiy6 : Ygqhw6);
assign U8n7v6 = (I4yiy6 ? R0bdt6 : U6yiy6);
assign U6yiy6 = (C7yiy6 | K7yiy6);
assign C7yiy6 = (S7yiy6 | A4yiy6);
assign A4yiy6 = (A8yiy6 & Ee47v6);
assign A8yiy6 = (Dbymz6[1] & Dbymz6[0]);
assign N8n7v6 = (~(I8yiy6 & Q8yiy6));
assign Q8yiy6 = (~(Y8yiy6 & Y9o7z6[1]));
assign I8yiy6 = (~(G9yiy6 & Ugo7z6[1]));
assign G8n7v6 = (O9yiy6 | W9yiy6);
assign O9yiy6 = (Wc0iw6 ? Eayiy6 : Oeo7z6[0]);
assign Eayiy6 = (~(Mayiy6 & Uayiy6));
assign Uayiy6 = (~(Oeo7z6[2] & Cbyiy6));
assign Cbyiy6 = (~(Kbyiy6 & Aiqhw6));
assign Mayiy6 = (~(Sbyiy6 & Acyiy6));
assign Z7n7v6 = (Icyiy6 ? L3bdt6 : F61iw6);
assign F61iw6 = (~(R1yhw6 | Qcyiy6));
assign Qcyiy6 = (Ycyiy6 & Gdyiy6);
assign Gdyiy6 = (Odyiy6 | Oh77z6);
assign Ycyiy6 = (~(On47v6 & Wdyiy6));
assign R1yhw6 = (~(Qjqhw6 ^ Xjqhw6));
assign Xjqhw6 = (JTAGNSW ? Hhxmz6[0] : Blxmz6[0]);
assign Qjqhw6 = (!Jjqhw6);
assign Jjqhw6 = (JTAGNSW ? Hhxmz6[1] : Blxmz6[1]);
assign S7n7v6 = (Q4yiy6 ? U3o7z6[11] : Fvb7z6[11]);
assign L7n7v6 = (~(Eeyiy6 & Meyiy6));
assign Meyiy6 = (~(Y8yiy6 & Y9o7z6[0]));
assign Eeyiy6 = (~(G9yiy6 & Ugo7z6[0]));
assign E7n7v6 = (Ueyiy6 ? Cxxmz6[1] : Ulxmz6[1]);
assign X6n7v6 = (!Cfyiy6);
assign Cfyiy6 = (V6wnv6 ? Kfyiy6 : M6giy6);
assign Kfyiy6 = (~(Pl0ft6 & Sfyiy6));
assign Q6n7v6 = (Q4yiy6 ? U3o7z6[10] : Fvb7z6[10]);
assign J6n7v6 = (Agyiy6 ? S2uhw6 : Ds57v6);
assign Agyiy6 = (~(Nwthw6 | J1uhw6));
assign Nwthw6 = (~(Rgxhw6 & Ccxhw6));
assign Ccxhw6 = (!Uzxmz6[3]);
assign Rgxhw6 = (Igyiy6 & Tbwhw6);
assign Igyiy6 = (Uzxmz6[1] & Axwhw6);
assign C6n7v6 = (Atthw6 ? Kp57v6 : S2uhw6);
assign Atthw6 = (Uwthw6 | J1uhw6);
assign Uwthw6 = (~(L4zhw6 & Oqwhw6));
assign Oqwhw6 = (~(Uzxmz6[3] | Uzxmz6[4]));
assign L4zhw6 = (Crwhw6 & L6xhw6);
assign Crwhw6 = (Uzxmz6[1] & Twwhw6);
assign Twwhw6 = (!Uzxmz6[0]);
assign S2uhw6 = (!Sdqhw6);
assign Sdqhw6 = (Dz1nv6 & K3a7z6);
assign K3a7z6 = (!SWDITMS);
assign V5n7v6 = (~(Qgyiy6 & Ygyiy6));
assign Ygyiy6 = (Ghyiy6 | Yg67z6);
assign O5n7v6 = (Ueyiy6 ? Cxxmz6[4] : Ulxmz6[4]);
assign H5n7v6 = (Ueyiy6 ? Cxxmz6[6] : Ulxmz6[6]);
assign A5n7v6 = (Ueyiy6 ? Cxxmz6[7] : Ulxmz6[7]);
assign T4n7v6 = (Ueyiy6 ? Cxxmz6[9] : Ulxmz6[9]);
assign M4n7v6 = (Ueyiy6 ? Cxxmz6[10] : Ulxmz6[10]);
assign F4n7v6 = (Ueyiy6 ? Cxxmz6[11] : Ulxmz6[11]);
assign Y3n7v6 = (Ueyiy6 ? Cxxmz6[12] : Ulxmz6[12]);
assign R3n7v6 = (Ueyiy6 ? Cxxmz6[28] : Ulxmz6[28]);
assign K3n7v6 = (Q4yiy6 ? U3o7z6[28] : Fvb7z6[28]);
assign D3n7v6 = (Ueyiy6 ? Cxxmz6[29] : Ulxmz6[29]);
assign W2n7v6 = (Q4yiy6 ? U3o7z6[29] : Fvb7z6[29]);
assign P2n7v6 = (Ueyiy6 ? Cxxmz6[30] : Ulxmz6[30]);
assign I2n7v6 = (Q4yiy6 ? U3o7z6[30] : Fvb7z6[30]);
assign B2n7v6 = (Ueyiy6 ? Cxxmz6[31] : Ulxmz6[31]);
assign U1n7v6 = (Ueyiy6 ? Cxxmz6[0] : Ulxmz6[0]);
assign N1n7v6 = (Qgyiy6 ? Usxmz6[0] : Yn57v6);
assign G1n7v6 = (Qgyiy6 ? Usxmz6[1] : Cl57v6);
assign Z0n7v6 = (Qgyiy6 ? E157v6 : Lothw6);
assign Qgyiy6 = (~(Ghyiy6 & Kp57v6));
assign Ghyiy6 = (Ekxhw6 & Bqthw6);
assign Bqthw6 = (Xh1nv6 & Npthw6);
assign Npthw6 = (!J1uhw6);
assign J1uhw6 = (B1ymz6[0] & Uc1nv6);
assign Uc1nv6 = (!Uia7z6);
assign Uia7z6 = (~(Ohyiy6 & Whyiy6));
assign Whyiy6 = (~(Eiyiy6 | Tzthw6));
assign Tzthw6 = (!B1ymz6[1]);
assign Eiyiy6 = (B1ymz6[2] | B1ymz6[3]);
assign Ohyiy6 = (B1ymz6[5] & B1ymz6[4]);
assign Xh1nv6 = (Tbwhw6 & Iuwhw6);
assign Iuwhw6 = (Uj1nv6 & Vbxhw6);
assign Vbxhw6 = (!Uzxmz6[1]);
assign Uj1nv6 = (~(Axwhw6 | Uzxmz6[3]));
assign Axwhw6 = (!Uzxmz6[4]);
assign Tbwhw6 = (Uzxmz6[0] & L6xhw6);
assign L6xhw6 = (!Uzxmz6[2]);
assign Ekxhw6 = (R7zhw6 & Qh1nv6);
assign Qh1nv6 = (!D857v6);
assign R7zhw6 = (Hf57v6 & Wd1nv6);
assign Wd1nv6 = (!Tq57v6);
assign Lothw6 = (!Ds57v6);
assign S0n7v6 = (Ueyiy6 ? Cxxmz6[2] : Ulxmz6[2]);
assign L0n7v6 = (Ueyiy6 ? Cxxmz6[23] : Ulxmz6[23]);
assign E0n7v6 = (Q4yiy6 ? U3o7z6[23] : Fvb7z6[23]);
assign Xzm7v6 = (Ueyiy6 ? Cxxmz6[22] : Ulxmz6[22]);
assign Qzm7v6 = (Q4yiy6 ? U3o7z6[22] : Fvb7z6[22]);
assign Jzm7v6 = (Ueyiy6 ? Cxxmz6[21] : Ulxmz6[21]);
assign Czm7v6 = (A0yiy6 ? Aixmz6[21] : L5ymz6[24]);
assign Vym7v6 = (Q4yiy6 ? U3o7z6[21] : Fvb7z6[21]);
assign Oym7v6 = (A0yiy6 ? Aixmz6[20] : L5ymz6[23]);
assign Hym7v6 = (Ueyiy6 ? Cxxmz6[20] : Ulxmz6[20]);
assign Aym7v6 = (Q4yiy6 ? U3o7z6[20] : Fvb7z6[20]);
assign Txm7v6 = (Ueyiy6 ? Cxxmz6[19] : Ulxmz6[19]);
assign Mxm7v6 = (A0yiy6 ? Aixmz6[19] : L5ymz6[22]);
assign Fxm7v6 = (Q4yiy6 ? U3o7z6[19] : Fvb7z6[19]);
assign Ywm7v6 = (A0yiy6 ? Aixmz6[18] : L5ymz6[21]);
assign Rwm7v6 = (Ueyiy6 ? Cxxmz6[18] : Ulxmz6[18]);
assign Kwm7v6 = (Q4yiy6 ? U3o7z6[18] : Fvb7z6[18]);
assign Dwm7v6 = (Ueyiy6 ? Cxxmz6[17] : Ulxmz6[17]);
assign Wvm7v6 = (A0yiy6 ? Aixmz6[17] : L5ymz6[20]);
assign Pvm7v6 = (Q4yiy6 ? U3o7z6[17] : Fvb7z6[17]);
assign Ivm7v6 = (A0yiy6 ? Aixmz6[16] : L5ymz6[19]);
assign Bvm7v6 = (Ueyiy6 ? Cxxmz6[16] : Ulxmz6[16]);
assign Uum7v6 = (Q4yiy6 ? U3o7z6[16] : Fvb7z6[16]);
assign Num7v6 = (Ueyiy6 ? Cxxmz6[15] : Ulxmz6[15]);
assign Gum7v6 = (A0yiy6 ? Aixmz6[15] : L5ymz6[18]);
assign Ztm7v6 = (Q4yiy6 ? U3o7z6[15] : Fvb7z6[15]);
assign Stm7v6 = (A0yiy6 ? Aixmz6[14] : L5ymz6[17]);
assign Ltm7v6 = (Ueyiy6 ? Cxxmz6[14] : Ulxmz6[14]);
assign Etm7v6 = (Q4yiy6 ? U3o7z6[14] : Fvb7z6[14]);
assign Xsm7v6 = (Ueyiy6 ? Cxxmz6[13] : Ulxmz6[13]);
assign Qsm7v6 = (A0yiy6 ? Aixmz6[13] : L5ymz6[16]);
assign Jsm7v6 = (Q4yiy6 ? U3o7z6[13] : Fvb7z6[13]);
assign Csm7v6 = (A0yiy6 ? Aixmz6[12] : L5ymz6[15]);
assign Vrm7v6 = (Q4yiy6 ? U3o7z6[12] : Fvb7z6[12]);
assign Orm7v6 = (~(Xczet6 ^ Aglov6));
assign Aglov6 = (~(Miyiy6 & Ejo7z6[0]));
assign Miyiy6 = (Ejo7z6[1] & Q7wnv6);
assign Hrm7v6 = (!Uiyiy6);
assign Uiyiy6 = (Kr97z6 ? Ua77z6 : Ma77z6);
assign Arm7v6 = (Zuixx6 ? O3uet6 : Cjyiy6);
assign Cjyiy6 = (~(Wp9ov6 | Dconv6));
assign Wp9ov6 = (~(Kjyiy6 & Sjyiy6));
assign Sjyiy6 = (Akyiy6 & Ikyiy6);
assign Akyiy6 = (~(Njkiw6 | Meoet6));
assign Kjyiy6 = (Qkyiy6 & Lbkiw6);
assign Qkyiy6 = (Ykyiy6 & Cfliy6);
assign Tqm7v6 = (Ueyiy6 ? Cxxmz6[3] : Ulxmz6[3]);
assign Mqm7v6 = (A0yiy6 ? Aixmz6[3] : L5ymz6[6]);
assign Fqm7v6 = (A0yiy6 ? Aixmz6[2] : L5ymz6[5]);
assign Ypm7v6 = (A0yiy6 ? Aixmz6[1] : L5ymz6[4]);
assign Rpm7v6 = (A0yiy6 ? Aixmz6[0] : L5ymz6[3]);
assign Kpm7v6 = (A0yiy6 ? Uixmz6[3] : L5ymz6[2]);
assign Dpm7v6 = (A0yiy6 ? Uixmz6[2] : L5ymz6[1]);
assign A0yiy6 = (!Q0yiy6);
assign Wom7v6 = (Icyiy6 ? Zn0ft6 : Cozet6);
assign Pom7v6 = (!Glyiy6);
assign Glyiy6 = (Wc0iw6 ? Olyiy6 : Rgqhw6);
assign Rgqhw6 = (!Oeo7z6[1]);
assign Iom7v6 = (Iownv6 ? Ekoet6 : Wlyiy6);
assign Wlyiy6 = (Ee3iw6 & M52iw6);
assign Ee3iw6 = (Emyiy6 & Mmyiy6);
assign Mmyiy6 = (~(M52iw6 & Umyiy6));
assign Umyiy6 = (~(Cnyiy6 & Knyiy6));
assign Knyiy6 = (~(Khoet6 | Wmoet6));
assign Cnyiy6 = (~(Snyiy6 | Aoyiy6));
assign Snyiy6 = (Ewyet6 & Ioyiy6);
assign Ioyiy6 = (Qln7z6[0] | Qln7z6[1]);
assign M52iw6 = (Qoyiy6 & Yoyiy6);
assign Qoyiy6 = (Hz1iw6 & Gpyiy6);
assign Gpyiy6 = (!Se3iw6);
assign Emyiy6 = (Se3iw6 ? Cjwiy6 : Opyiy6);
assign Se3iw6 = (Gyjiw6 & Wcmov6);
assign Gyjiw6 = (!Lgonv6);
assign Cjwiy6 = (Wpyiy6 & Eqyiy6);
assign Eqyiy6 = (Mqyiy6 & Uqyiy6);
assign Mqyiy6 = (~(Bzjiw6 | Qboet6));
assign Wpyiy6 = (Cryiy6 & Kryiy6);
assign Opyiy6 = (Yoyiy6 & Hz1iw6);
assign Bom7v6 = (~(Sryiy6 & Asyiy6));
assign Asyiy6 = (~(Isyiy6 & Ppzet6));
assign Isyiy6 = (O4qhw6 & Kr97z6);
assign Sryiy6 = (~(Tszet6 & Qsyiy6));
assign Qsyiy6 = (T1zhw6 | O4qhw6);
assign O4qhw6 = (~(Ysyiy6 | Silov6));
assign Silov6 = (Gtyiy6 & Wc0iw6);
assign Gtyiy6 = (~(K7yiy6 | S7yiy6));
assign S7yiy6 = (Olyiy6 & M6yiy6);
assign K7yiy6 = (M6yiy6 & Otyiy6);
assign M6yiy6 = (Wtyiy6 & Euyiy6);
assign Wtyiy6 = (Oeo7z6[2] ? Uuyiy6 : Muyiy6);
assign Uuyiy6 = (~(Cvyiy6 & Kvyiy6));
assign Kvyiy6 = (Svyiy6 & Naonv6);
assign Naonv6 = (!O7o7z6[2]);
assign Svyiy6 = (Ic0iw6 & Awyiy6);
assign Awyiy6 = (!Oeo7z6[0]);
assign Ic0iw6 = (!Gco7z6[4]);
assign Cvyiy6 = (Gco7z6[5] & Aiqhw6);
assign Aiqhw6 = (!Frzet6);
assign Muyiy6 = (Otyiy6 | Acyiy6);
assign Acyiy6 = (~(Cb77z6 & Sfyiy6));
assign Unm7v6 = (!Iwyiy6);
assign Iwyiy6 = (V6wnv6 ? Qwyiy6 : Jie7x6);
assign Qwyiy6 = (~(O7o7z6[2] | Ywyiy6));
assign Nnm7v6 = (He1iw6 ? Hhxmz6[0] : L5ymz6[5]);
assign Gnm7v6 = (He1iw6 ? Hhxmz6[1] : L5ymz6[6]);
assign Zmm7v6 = (He1iw6 ? Ogxmz6[0] : L5ymz6[11]);
assign Smm7v6 = (He1iw6 ? Ogxmz6[1] : L5ymz6[12]);
assign Lmm7v6 = (He1iw6 ? Ogxmz6[2] : L5ymz6[13]);
assign Emm7v6 = (He1iw6 ? Ogxmz6[3] : L5ymz6[14]);
assign Xlm7v6 = (He1iw6 ? Qf47v6 : L5ymz6[29]);
assign Qlm7v6 = (He1iw6 ? Mg47v6 : L5ymz6[33]);
assign Jlm7v6 = (He1iw6 ? Kh47v6 : L5ymz6[31]);
assign Clm7v6 = (He1iw6 ? Ez57v6 : L5ymz6[3]);
assign He1iw6 = (~(Gxyiy6 & Oxyiy6));
assign Oxyiy6 = (Qo1nv6 & Wxyiy6);
assign Gxyiy6 = (L5ymz6[1] & Su1iw6);
assign Vkm7v6 = (Eyyiy6 ? Uixmz6[25] : L5ymz6[28]);
assign Okm7v6 = (Eyyiy6 ? Uixmz6[26] : L5ymz6[29]);
assign Hkm7v6 = (Eyyiy6 ? Uixmz6[27] : L5ymz6[30]);
assign Akm7v6 = (Eyyiy6 ? Uixmz6[28] : L5ymz6[31]);
assign Tjm7v6 = (Eyyiy6 ? Uixmz6[29] : L5ymz6[32]);
assign Eyyiy6 = (!Myyiy6);
assign Mjm7v6 = (Myyiy6 ? L5ymz6[33] : Uixmz6[30]);
assign Fjm7v6 = (Myyiy6 ? L5ymz6[34] : Uixmz6[31]);
assign Yim7v6 = (Myyiy6 ? L5ymz6[7] : Uixmz6[4]);
assign Rim7v6 = (Myyiy6 ? L5ymz6[8] : Uixmz6[5]);
assign Kim7v6 = (Ueyiy6 ? Cxxmz6[25] : Ulxmz6[25]);
assign Dim7v6 = (Q4yiy6 ? U3o7z6[25] : Fvb7z6[25]);
assign Whm7v6 = (Vjqnv6 ? Aym7z6[1] : Hjqnv6);
assign Phm7v6 = (Vjqnv6 ? Aym7z6[2] : Yhqnv6);
assign Ihm7v6 = (Vjqnv6 ? Aym7z6[3] : Pgqnv6);
assign Bhm7v6 = (Iownv6 ? Dtm7z6[3] : Az1iw6);
assign Iownv6 = (~(Q7wnv6 | L1bdt6));
assign Q7wnv6 = (~(Uyyiy6 & Czyiy6));
assign Czyiy6 = (Kzyiy6 & Szyiy6);
assign Szyiy6 = (~(Dtm7z6[2] & Vd2iw6));
assign Kzyiy6 = (A0ziy6 & I0ziy6);
assign I0ziy6 = (~(Dtm7z6[0] & HREADYD));
assign A0ziy6 = (~(Dtm7z6[3] & Q0ziy6));
assign Uyyiy6 = (I6oet6 & Y0ziy6);
assign Y0ziy6 = (~(Dtm7z6[1] & HREADYS));
assign Az1iw6 = (~(G1ziy6 & O1ziy6));
assign O1ziy6 = (Bownv6 | Go9ov6);
assign Bownv6 = (K7giy6 | Yoyiy6);
assign Yoyiy6 = (!Oz1iw6);
assign G1ziy6 = (W1ziy6 & E2ziy6);
assign W1ziy6 = (~(Aoyiy6 & I2yet6));
assign Ugm7v6 = (Ueyiy6 ? Cxxmz6[27] : Ulxmz6[27]);
assign Ngm7v6 = (Q4yiy6 ? U3o7z6[27] : Fvb7z6[27]);
assign Ggm7v6 = (Ueyiy6 ? Cxxmz6[26] : Ulxmz6[26]);
assign Zfm7v6 = (Q4yiy6 ? U3o7z6[26] : Fvb7z6[26]);
assign Sfm7v6 = (Ueyiy6 ? Cxxmz6[5] : Ulxmz6[5]);
assign Lfm7v6 = (Q4yiy6 ? U3o7z6[9] : Fvb7z6[9]);
assign Efm7v6 = (Q4yiy6 ? U3o7z6[8] : Fvb7z6[8]);
assign Xem7v6 = (Ueyiy6 ? Cxxmz6[8] : Ulxmz6[8]);
assign Qem7v6 = (Q4yiy6 ? U3o7z6[7] : Fvb7z6[7]);
assign Jem7v6 = (Q4yiy6 ? U3o7z6[6] : Fvb7z6[6]);
assign Cem7v6 = (Q4yiy6 ? U3o7z6[5] : Fvb7z6[5]);
assign Vdm7v6 = (Q4yiy6 ? U3o7z6[4] : Fvb7z6[4]);
assign Odm7v6 = (M2ziy6 | U2ziy6);
assign U2ziy6 = (Y8yiy6 & Y9o7z6[3]);
assign M2ziy6 = (G9yiy6 ? Fvb7z6[3] : C3ziy6);
assign C3ziy6 = (Ib1iw6 & F5o7z6[3]);
assign Hdm7v6 = (K3ziy6 | S3ziy6);
assign S3ziy6 = (Y8yiy6 & Y9o7z6[2]);
assign Y8yiy6 = (~(Ib1iw6 | G9yiy6));
assign Ib1iw6 = (!A4ziy6);
assign K3ziy6 = (G9yiy6 ? Fvb7z6[2] : I4ziy6);
assign I4ziy6 = (~(A4ziy6 | X11iw6));
assign X11iw6 = (!F5o7z6[2]);
assign A4ziy6 = (~(F5o7z6[4] & Pb1iw6));
assign Pb1iw6 = (~(Q4ziy6 | F5o7z6[5]));
assign Q4ziy6 = (F5o7z6[6] | F5o7z6[7]);
assign Adm7v6 = (Icyiy6 ? K2bdt6 : Qmzet6);
assign Tcm7v6 = (Ueyiy6 ? Cxxmz6[24] : Ulxmz6[24]);
assign Ueyiy6 = (~(Werhw6 | Yg67z6));
assign Werhw6 = (!M257v6);
assign Mcm7v6 = (Q4yiy6 ? U3o7z6[24] : Fvb7z6[24]);
assign Q4yiy6 = (!G9yiy6);
assign G9yiy6 = (Y4ziy6 & Icyiy6);
assign Icyiy6 = (!V6wnv6);
assign V6wnv6 = (~(Dnh7v6 ^ Hgzet6));
assign Y4ziy6 = (Wmh7v6 ^ Mezet6);
assign Fcm7v6 = (Myyiy6 ? L5ymz6[9] : Uixmz6[6]);
assign Ybm7v6 = (Myyiy6 ? L5ymz6[10] : Uixmz6[7]);
assign Rbm7v6 = (Myyiy6 ? L5ymz6[27] : Uixmz6[24]);
assign Myyiy6 = (G5ziy6 & O5ziy6);
assign O5ziy6 = (Qo1nv6 & W5ziy6);
assign Qo1nv6 = (!L5ymz6[0]);
assign G5ziy6 = (L5ymz6[2] & Su1iw6);
assign Kbm7v6 = (!E6ziy6);
assign E6ziy6 = (Q0yiy6 ? L5ymz6[0] : Oh77z6);
assign Q0yiy6 = (M6ziy6 & Xf1iw6);
assign Xf1iw6 = (~(F267v6 | S067v6));
assign M6ziy6 = (K9qhw6 & Eg1iw6);
assign Eg1iw6 = (~(Sx57v6 & Ez57v6));
assign K9qhw6 = (U6ziy6 & C7ziy6);
assign U6ziy6 = (W6ymz6[0] & W6ymz6[1]);
assign Dbm7v6 = (Dc1iw6 ? Q2ymz6[1] : K7ziy6);
assign K7ziy6 = (~(L5ymz6[1] & Wxyiy6));
assign Wxyiy6 = (!L5ymz6[2]);
assign Wam7v6 = (Dc1iw6 ? Q2ymz6[0] : S7ziy6);
assign Dc1iw6 = (!Su1iw6);
assign Su1iw6 = (Tm1nv6 & C7ziy6);
assign C7ziy6 = (A8ziy6 & By1nv6);
assign By1nv6 = (I8ziy6 & Lw1nv6);
assign Lw1nv6 = (R9ymz6[0] & Gq1nv6);
assign Gq1nv6 = (!R9ymz6[1]);
assign I8ziy6 = (R9ymz6[2] & K3whw6);
assign K3whw6 = (!R9ymz6[3]);
assign A8ziy6 = (Co1nv6 & W1yiy6);
assign W1yiy6 = (!Wh77z6);
assign Co1nv6 = (W6ymz6[3] & Mm1nv6);
assign Mm1nv6 = (!W6ymz6[2]);
assign Tm1nv6 = (W6ymz6[1] & Jo1nv6);
assign Jo1nv6 = (!W6ymz6[0]);
assign S7ziy6 = (~(L5ymz6[2] & W5ziy6));
assign W5ziy6 = (!L5ymz6[1]);
assign Pam7v6 = (P9get6 ? Qmj7z6[5] : Jqj7z6[5]);
assign Qmj7z6[5] = (~(Q8ziy6 | Y8ziy6));
assign Iam7v6 = (Cpsnv6 ? G9ziy6 : N6c7v6);
assign Cpsnv6 = (~(O9ziy6 & Wfo7v6));
assign O9ziy6 = (Kgbdt6 & Jgliw6);
assign G9ziy6 = (H8c7v6 & Detnv6);
assign Detnv6 = (!W9c7v6);
assign Bam7v6 = (P9get6 ? Pnfet6 : Jqj7z6[2]);
assign Pnfet6 = (~(Y8ziy6 | W9ziy6));
assign Y8ziy6 = (!Ykliy6);
assign U9m7v6 = (Otshy6 ? Xfymz6[11] : Pjb7z6[11]);
assign N9m7v6 = (Otshy6 ? Xfymz6[10] : Pjb7z6[10]);
assign G9m7v6 = (Otshy6 ? Xfymz6[9] : Pjb7z6[9]);
assign Z8m7v6 = (Otshy6 ? Xfymz6[8] : Pjb7z6[8]);
assign S8m7v6 = (Otshy6 ? Xfymz6[7] : Pjb7z6[7]);
assign L8m7v6 = (Otshy6 ? Xfymz6[6] : Pjb7z6[6]);
assign E8m7v6 = (Otshy6 ? Xfymz6[5] : Pjb7z6[5]);
assign X7m7v6 = (Otshy6 ? Xfymz6[4] : Pjb7z6[4]);
assign Q7m7v6 = (Otshy6 ? Xfymz6[3] : Pjb7z6[3]);
assign J7m7v6 = (Maziy6 ? Ti2nz6[4] : Eaziy6);
assign Eaziy6 = (Uaziy6 & Cbziy6);
assign Cbziy6 = (~(Kbziy6 | Pjb7z6[7]));
assign Kbziy6 = (Pjb7z6[8] | Pjb7z6[9]);
assign Uaziy6 = (~(Sbziy6 | Pjb7z6[10]));
assign Sbziy6 = (Pjb7z6[11] | Pjb7z6[6]);
assign C7m7v6 = (Maziy6 ? Ti2nz6[3] : Pjb7z6[5]);
assign V6m7v6 = (Cjliy6 ? Pjb7z6[4] : Ti2nz6[2]);
assign O6m7v6 = (Cjliy6 ? Pjb7z6[3] : Ti2nz6[1]);
assign H6m7v6 = (Qgnhy6 ? J02nz6[3] : Pjb7z6[3]);
assign A6m7v6 = (Qgnhy6 ? J02nz6[4] : Pjb7z6[4]);
assign T5m7v6 = (Qgnhy6 ? J02nz6[5] : Pjb7z6[5]);
assign M5m7v6 = (Qgnhy6 ? J02nz6[6] : Pjb7z6[6]);
assign F5m7v6 = (Qgnhy6 ? J02nz6[7] : Pjb7z6[7]);
assign Y4m7v6 = (Qgnhy6 ? J02nz6[8] : Pjb7z6[8]);
assign R4m7v6 = (Qgnhy6 ? J02nz6[9] : Pjb7z6[9]);
assign K4m7v6 = (Qgnhy6 ? J02nz6[10] : Pjb7z6[10]);
assign D4m7v6 = (Qgnhy6 ? J02nz6[11] : Pjb7z6[11]);
assign W3m7v6 = (Kr97z6 ? Acziy6 : Rjzet6);
assign Acziy6 = (L6qhw6 & Icziy6);
assign Icziy6 = (~(Wc0iw6 & Qcziy6));
assign Qcziy6 = (~(Olyiy6 & Otyiy6));
assign Otyiy6 = (!Sbyiy6);
assign Sbyiy6 = (Pc0iw6 & Ycziy6);
assign Olyiy6 = (Euyiy6 & Gdziy6);
assign Gdziy6 = (~(Odziy6 & Pc0iw6));
assign Odziy6 = (Wdziy6 & Ygqhw6);
assign Ygqhw6 = (!Oeo7z6[2]);
assign Wdziy6 = (~(Ycziy6 & Eeziy6));
assign Eeziy6 = (~(Cb77z6 & Ywyiy6));
assign Euyiy6 = (~(Meziy6 & Ueziy6));
assign Ueziy6 = (~(W9yiy6 | Frzet6));
assign Meziy6 = (Oeo7z6[2] & Cfziy6);
assign Cfziy6 = (Kbyiy6 | Oeo7z6[1]);
assign Kbyiy6 = (O7o7z6[0] & Oeo7z6[0]);
assign O7o7z6[0] = (~(O7o7z6[2] | Pl0ft6));
assign Wc0iw6 = (!I4yiy6);
assign I4yiy6 = (L6qhw6 ? Sfziy6 : Kfziy6);
assign Sfziy6 = (~(Kr97z6 & Agziy6));
assign Agziy6 = (~(Pc0iw6 & Igziy6));
assign Igziy6 = (~(Qgziy6 & Kgqhw6));
assign Kgqhw6 = (~(Ygziy6 & Ghziy6));
assign Ghziy6 = (~(Ohziy6 & Whziy6));
assign Whziy6 = (Eiziy6 & Miziy6);
assign Miziy6 = (~(Uiziy6 | Omxmz6[29]));
assign Uiziy6 = (Omxmz6[30] | Omxmz6[31]);
assign Eiziy6 = (~(Omxmz6[27] | Omxmz6[28]));
assign Ohziy6 = (Cjziy6 & Kjziy6);
assign Kjziy6 = (~(Omxmz6[25] | Omxmz6[26]));
assign Cjziy6 = (S397z6 & Wdyiy6);
assign Ygziy6 = (~(Sjziy6 & Akziy6));
assign Akziy6 = (Ikziy6 & Qkziy6);
assign Qkziy6 = (~(Ykziy6 | Uixmz6[29]));
assign Ykziy6 = (Uixmz6[30] | Uixmz6[31]);
assign Ikziy6 = (~(Uixmz6[27] | Uixmz6[28]));
assign Sjziy6 = (Glziy6 & Olziy6);
assign Olziy6 = (~(Uixmz6[25] | Uixmz6[26]));
assign Glziy6 = (~(Odyiy6 | Uixmz6[24]));
assign Odyiy6 = (!Wlziy6);
assign Qgziy6 = (~(Emziy6 & Ycziy6));
assign Ycziy6 = (Swzhw6 & Mmziy6);
assign Mmziy6 = (~(Umziy6 & Cnziy6));
assign Cnziy6 = (Knziy6 & Wmqhw6);
assign Knziy6 = (Knqhw6 & Pmqhw6);
assign Umziy6 = (Imqhw6 & Dnqhw6);
assign Swzhw6 = (~(Snziy6 & Aoziy6));
assign Aoziy6 = (!Pmqhw6);
assign Snziy6 = (~(Ioziy6 | Imqhw6));
assign Imqhw6 = (~(Qoziy6 & Yoziy6));
assign Yoziy6 = (~(Uixmz6[3] & Wlziy6));
assign Qoziy6 = (~(Omxmz6[3] & Wdyiy6));
assign Emziy6 = (Gpziy6 & Sfyiy6);
assign Sfyiy6 = (!Ywyiy6);
assign Ywyiy6 = (Opziy6 & Pmqhw6);
assign Pmqhw6 = (~(Wpziy6 & Eqziy6));
assign Eqziy6 = (~(Uixmz6[4] & Wlziy6));
assign Wpziy6 = (~(Omxmz6[4] & Wdyiy6));
assign Gpziy6 = (~(Opziy6 & Ulqhw6));
assign Ulqhw6 = (~(Mqziy6 & Uqziy6));
assign Uqziy6 = (~(Uixmz6[2] & Wlziy6));
assign Mqziy6 = (~(Omxmz6[2] & Wdyiy6));
assign Opziy6 = (!Ioziy6);
assign Ioziy6 = (~(Crziy6 & Krziy6));
assign Krziy6 = (!Knqhw6);
assign Knqhw6 = (~(Srziy6 & Asziy6));
assign Asziy6 = (~(Uixmz6[7] & Wlziy6));
assign Srziy6 = (~(Omxmz6[7] & Wdyiy6));
assign Crziy6 = (~(Wmqhw6 | Dnqhw6));
assign Dnqhw6 = (~(Isziy6 & Qsziy6));
assign Qsziy6 = (~(Uixmz6[6] & Wlziy6));
assign Isziy6 = (~(Omxmz6[6] & Wdyiy6));
assign Wmqhw6 = (~(Ysziy6 & Gtziy6));
assign Gtziy6 = (~(Uixmz6[5] & Wlziy6));
assign Wlziy6 = (~(E6qhw6 | Dz1nv6));
assign Ysziy6 = (~(Omxmz6[5] & Wdyiy6));
assign Wdyiy6 = (~(E6qhw6 | JTAGNSW));
assign E6qhw6 = (!Dbymz6[0]);
assign Pc0iw6 = (~(Oeo7z6[1] | Oeo7z6[0]));
assign Kfziy6 = (~(Kr97z6 & Otziy6));
assign Otziy6 = (Ysyiy6 | Tszet6);
assign Ysyiy6 = (Ua77z6 ^ Ma77z6);
assign L6qhw6 = (~(Oeo7z6[2] | W9yiy6));
assign W9yiy6 = (Oeo7z6[1] & Oeo7z6[0]);
assign P3m7v6 = (Wtziy6 ? Cx4iw6 : H1j7z6[23]);
assign I3m7v6 = (Wtziy6 ? D85iw6 : H1j7z6[22]);
assign B3m7v6 = (Wtziy6 ? Ej5iw6 : H1j7z6[21]);
assign U2m7v6 = (Wtziy6 ? Bl5iw6 : H1j7z6[20]);
assign N2m7v6 = (Wtziy6 ? Mn5iw6 : H1j7z6[19]);
assign G2m7v6 = (Wtziy6 ? Jp5iw6 : H1j7z6[18]);
assign Z1m7v6 = (Wtziy6 ? Gr5iw6 : H1j7z6[17]);
assign S1m7v6 = (Euziy6 ? Z0iov6 : H1j7z6[15]);
assign L1m7v6 = (Euziy6 ? Bk6iw6 : H1j7z6[14]);
assign E1m7v6 = (Euziy6 ? Guhov6 : H1j7z6[13]);
assign X0m7v6 = (Euziy6 ? Emhov6 : H1j7z6[12]);
assign Q0m7v6 = (Euziy6 ? Dz6iw6 : H1j7z6[11]);
assign J0m7v6 = (Euziy6 ? H17iw6 : H1j7z6[10]);
assign C0m7v6 = (Euziy6 ? J27iw6 : H1j7z6[9]);
assign Vzl7v6 = (Muziy6 ? U42nv6 : H1j7z6[0]);
assign Ozl7v6 = (Muziy6 ? R62nv6 : H1j7z6[7]);
assign Hzl7v6 = (Muziy6 ? K62nv6 : H1j7z6[6]);
assign Azl7v6 = (Muziy6 ? D62nv6 : H1j7z6[5]);
assign Tyl7v6 = (Muziy6 ? W52nv6 : H1j7z6[4]);
assign Myl7v6 = (Muziy6 ? P52nv6 : H1j7z6[3]);
assign Fyl7v6 = (Muziy6 ? B52nv6 : H1j7z6[1]);
assign Yxl7v6 = (~(Uuziy6 & Cvziy6));
assign Cvziy6 = (~(T7j7z6[0] & Kvziy6));
assign Uuziy6 = (~(Svziy6 & Hq3iw6));
assign Rxl7v6 = (~(Awziy6 & Iwziy6));
assign Iwziy6 = (~(T7j7z6[2] & Kvziy6));
assign Awziy6 = (~(Svziy6 & Gg2iw6));
assign Kxl7v6 = (~(Qwziy6 & Ywziy6));
assign Ywziy6 = (~(T7j7z6[1] & Kvziy6));
assign Kvziy6 = (~(Svziy6 & Bqi7z6[3]));
assign Qwziy6 = (~(Svziy6 & Nf3iw6));
assign Dxl7v6 = (~(Gxziy6 & Oxziy6));
assign Oxziy6 = (~(Z8j7z6[0] & Wxziy6));
assign Gxziy6 = (~(Svziy6 & T95iw6));
assign Wwl7v6 = (~(Eyziy6 & Myziy6));
assign Myziy6 = (~(Z8j7z6[2] & Wxziy6));
assign Eyziy6 = (~(Svziy6 & Qj4iw6));
assign Pwl7v6 = (~(Uyziy6 & Czziy6));
assign Czziy6 = (~(Z8j7z6[1] & Wxziy6));
assign Wxziy6 = (~(Svziy6 & Bqi7z6[2]));
assign Uyziy6 = (~(Svziy6 & Zy4iw6));
assign Iwl7v6 = (~(Kzziy6 & Szziy6));
assign Szziy6 = (~(Nbj7z6[0] & A00jy6));
assign Kzziy6 = (~(Svziy6 & X18iw6));
assign Bwl7v6 = (~(I00jy6 & Q00jy6));
assign Q00jy6 = (~(Nbj7z6[2] & A00jy6));
assign I00jy6 = (~(Svziy6 & O87iw6));
assign Uvl7v6 = (~(Y00jy6 & G10jy6));
assign G10jy6 = (~(Nbj7z6[1] & A00jy6));
assign A00jy6 = (~(Svziy6 & Bqi7z6[0]));
assign Y00jy6 = (~(Svziy6 & Np7iw6));
assign Svziy6 = (O10jy6 & Eec7x6);
assign O10jy6 = (Wdm7x6 & Pb8iw6);
assign Nvl7v6 = (W10jy6 ? Micet6 : Jp5iw6);
assign Gvl7v6 = (W10jy6 ? Sjcet6 : Gr5iw6);
assign Zul7v6 = (P9get6 ? Oqbet6 : Jqj7z6[7]);
assign Oqbet6 = (Q0hov6 & W14iw6);
assign Q0hov6 = (E20jy6 & Wdm7x6);
assign E20jy6 = (Z4m7x6 & Bqi7z6[3]);
assign Sul7v6 = (M20jy6 ? D5cet6 : B52nv6);
assign Lul7v6 = (M20jy6 ? L2cet6 : W52nv6);
assign Eul7v6 = (U20jy6 ? A8cet6 : U42nv6);
assign Xtl7v6 = (U20jy6 ? E9cet6 : B52nv6);
assign Qtl7v6 = (Ijeet6 & Nbmov6);
assign Nbmov6 = (!Mleet6);
assign Jtl7v6 = (T8lov6 ? Qij7z6[6] : K62nv6);
assign Ctl7v6 = (T8lov6 ? Qij7z6[5] : D62nv6);
assign Vsl7v6 = (T8lov6 ? Qij7z6[4] : W52nv6);
assign Osl7v6 = (T8lov6 ? Qij7z6[3] : P52nv6);
assign Hsl7v6 = (T8lov6 ? Qij7z6[1] : B52nv6);
assign T8lov6 = (!Knniy6);
assign Asl7v6 = (Knniy6 ? U42nv6 : Qij7z6[0]);
assign Trl7v6 = (~(C30jy6 & K30jy6));
assign K30jy6 = (~(S30jy6 & Hq3iw6));
assign C30jy6 = (~(Gaj7z6[0] & A40jy6));
assign Mrl7v6 = (~(I40jy6 & Q40jy6));
assign Q40jy6 = (~(S30jy6 & Gg2iw6));
assign Gg2iw6 = (~(Dv3iw6 | Fcgiw6));
assign I40jy6 = (~(Gaj7z6[2] & A40jy6));
assign Frl7v6 = (~(Y40jy6 & G50jy6));
assign G50jy6 = (~(S30jy6 & Nf3iw6));
assign Nf3iw6 = (~(Dv3iw6 | Wagiw6));
assign Y40jy6 = (~(Gaj7z6[1] & A40jy6));
assign A40jy6 = (~(S30jy6 & Bqi7z6[3]));
assign S30jy6 = (L28iw6 & Z4m7x6);
assign Z4m7x6 = (O50jy6 & Pi8iw6);
assign O50jy6 = (G42nv6 & Toi7z6[2]);
assign Yql7v6 = (W50jy6 ? Wf4iw6 : HTMDHBURST[0]);
assign W50jy6 = (E60jy6 & Bqi7z6[3]);
assign Rql7v6 = (~(K94iw6 & M60jy6));
assign M60jy6 = (~(HTMDHREADY & Kygnv6));
assign Kql7v6 = (Kygnv6 ? HTMDHRESP[1] : U60jy6);
assign U60jy6 = (C70jy6 & K70jy6);
assign K70jy6 = (~(S70jy6 & A80jy6));
assign A80jy6 = (~(HRESPS[1] & Ad47x6));
assign S70jy6 = (~(HRESPD[1] & Mc47x6));
assign Dql7v6 = (Kygnv6 ? HTMDHRESP[0] : I80jy6);
assign I80jy6 = (Ihnet6 | A0onv6);
assign A0onv6 = (!Qvkiw6);
assign Qvkiw6 = (~(C70jy6 & Q80jy6));
assign Q80jy6 = (~(Y80jy6 & G90jy6));
assign G90jy6 = (O90jy6 & W90jy6);
assign W90jy6 = (~(Zmoyx6 & Qhlov6));
assign Qhlov6 = (~(Ea0jy6 & Ma0jy6));
assign Ma0jy6 = (~(Ua0jy6 & Cb0jy6));
assign Cb0jy6 = (~(Kb0jy6 | Sb0jy6));
assign Ua0jy6 = (Ac0jy6 & Ic0jy6);
assign Ic0jy6 = (!Ozixx6);
assign Ea0jy6 = (Qc0jy6 | W5eiw6);
assign W5eiw6 = (~(Yc0jy6 & Gd0jy6));
assign Gd0jy6 = (Ac0jy6 | Teyet6);
assign Yc0jy6 = (~(Qmonv6 | Sjyet6));
assign Qc0jy6 = (~(Znn7z6[3] & Od0jy6));
assign Od0jy6 = (Vugxx6 | Znn7z6[0]);
assign O90jy6 = (~(Kfdiy6 & Xhlov6));
assign Xhlov6 = (~(Wd0jy6 & Ee0jy6));
assign Ee0jy6 = (~(Euget6 & Klo7z6[5]));
assign Wd0jy6 = (Me0jy6 & Ue0jy6);
assign Ue0jy6 = (~(Ja1ft6 & Cf0jy6));
assign Me0jy6 = (~(P8adt6 & Ngqyx6));
assign Y80jy6 = (Kf0jy6 & Sf0jy6);
assign Sf0jy6 = (~(HRESPS[0] & Ad47x6));
assign Kf0jy6 = (~(HRESPD[0] & Mc47x6));
assign C70jy6 = (~(Suixx6 | Yg77z6));
assign Wpl7v6 = (~(Nlh7v6 & K94iw6));
assign K94iw6 = (!Ob4iw6);
assign Ob4iw6 = (HTMDHBURST[0] & O5a7z6);
assign O5a7z6 = (Senet6 & Rsdiw6);
assign Rsdiw6 = (Qgwiy6 | Suixx6);
assign Suixx6 = (!Ag0jy6);
assign Qgwiy6 = (~(Ig0jy6 & Qg0jy6));
assign Qg0jy6 = (Yg0jy6 & Gh0jy6);
assign Gh0jy6 = (~(HREADYS & Ad47x6));
assign Ad47x6 = (Rnm7z6[1] & Oh0jy6);
assign Yg0jy6 = (~(Wh0jy6 | Yg77z6));
assign Wh0jy6 = (Ei0jy6 & Mi0jy6);
assign Mi0jy6 = (Ui0jy6 & Cj0jy6);
assign Cj0jy6 = (~(Kj0jy6 & Zuixx6));
assign Kj0jy6 = (~(HREADYD & Sj0jy6));
assign Sj0jy6 = (~(Ak0jy6 & Ik0jy6));
assign Ak0jy6 = (Qk0jy6 & Ag0jy6);
assign Ui0jy6 = (~(Yk0jy6 & Gl0jy6));
assign Ei0jy6 = (D6eiw6 & Zmoyx6);
assign Zmoyx6 = (Kryiy6 & Ol0jy6);
assign Ol0jy6 = (~(I497z6 & Wl0jy6));
assign Ig0jy6 = (Em0jy6 & Mm0jy6);
assign Mm0jy6 = (~(Kfdiy6 & Vd2iw6));
assign Vd2iw6 = (~(Um0jy6 & Cn0jy6));
assign Cn0jy6 = (Kn0jy6 & Xneiw6);
assign Xneiw6 = (Sn0jy6 | Ngqyx6);
assign Sn0jy6 = (Cf0jy6 | Klo7z6[5]);
assign Cf0jy6 = (~(Ao0jy6 & I4fiy6));
assign Kn0jy6 = (~(Klo7z6[5] & Orget6));
assign Um0jy6 = (Io0jy6 & Qo0jy6);
assign Qo0jy6 = (~(O9adt6 & Ngqyx6));
assign Ngqyx6 = (Klo7z6[4] | Klo7z6[6]);
assign Io0jy6 = (A497z6 | Yo0jy6);
assign Yo0jy6 = (Ao0jy6 & Gp0jy6);
assign Gp0jy6 = (I4fiy6 | D16ft6);
assign I4fiy6 = (!Klo7z6[3]);
assign Ao0jy6 = (Op0jy6 & F41zx6);
assign F41zx6 = (!Klo7z6[0]);
assign Op0jy6 = (~(Klo7z6[1] | Klo7z6[2]));
assign Kfdiy6 = (Rnm7z6[2] & Oh0jy6);
assign Em0jy6 = (~(Mc47x6 & HREADYD));
assign Mc47x6 = (Rnm7z6[0] & Oh0jy6);
assign Oh0jy6 = (Kryiy6 & Wl0jy6);
assign Wl0jy6 = (~(Wp0jy6 & Styet6));
assign Wp0jy6 = (~(Eq0jy6 | A9gxx6));
assign Ppl7v6 = (Mq0jy6 ? J27iw6 : X0eet6);
assign Ipl7v6 = (Mq0jy6 ? H17iw6 : W2eet6);
assign Bpl7v6 = (Mq0jy6 ? U47iw6 : Yydet6);
assign Mq0jy6 = (~(Uq0jy6 | Nq6iw6));
assign Uol7v6 = (Cr0jy6 ? Brdet6 : W52nv6);
assign Nol7v6 = (~(Kr0jy6 & Sr0jy6));
assign Sr0jy6 = (~(Zsdet6 & Cr0jy6));
assign Kr0jy6 = (~(X18iw6 & E60jy6));
assign Gol7v6 = (~(As0jy6 & Is0jy6));
assign Is0jy6 = (~(Zudet6 & Cr0jy6));
assign As0jy6 = (~(Np7iw6 & E60jy6));
assign Znl7v6 = (~(Qs0jy6 & Ys0jy6));
assign Ys0jy6 = (~(Ywdet6 & Cr0jy6));
assign Qs0jy6 = (~(O87iw6 & E60jy6));
assign Snl7v6 = (Cr0jy6 ? Zodet6 : U42nv6);
assign Cr0jy6 = (Uq0jy6 | Twaiw6);
assign Lnl7v6 = (Hyhov6 ? Mn5iw6 : Nybet6);
assign Enl7v6 = (Hyhov6 ? Jp5iw6 : Vzbet6);
assign Xml7v6 = (~(Gt0jy6 & Ot0jy6));
assign Ot0jy6 = (~(Tcj7z6[0] & Wt0jy6));
assign Gt0jy6 = (~(Eu0jy6 & T95iw6));
assign T95iw6 = (~(Ie5iw6 | Tyfiw6));
assign Qml7v6 = (~(Mu0jy6 & Uu0jy6));
assign Uu0jy6 = (~(Tcj7z6[2] & Wt0jy6));
assign Mu0jy6 = (~(Eu0jy6 & Qj4iw6));
assign Qj4iw6 = (~(Ie5iw6 | L1giw6));
assign Jml7v6 = (~(Cv0jy6 & Kv0jy6));
assign Kv0jy6 = (~(Tcj7z6[1] & Wt0jy6));
assign Wt0jy6 = (~(Eu0jy6 & Bqi7z6[2]));
assign Cv0jy6 = (~(Eu0jy6 & Zy4iw6));
assign Cml7v6 = (~(Sv0jy6 & Aw0jy6));
assign Aw0jy6 = (~(Ffj7z6[0] & Iw0jy6));
assign Sv0jy6 = (~(Eu0jy6 & X18iw6));
assign X18iw6 = (~(Twaiw6 | Tdfiw6));
assign Vll7v6 = (~(Qw0jy6 & Yw0jy6));
assign Yw0jy6 = (~(Ffj7z6[2] & Iw0jy6));
assign Qw0jy6 = (~(Eu0jy6 & O87iw6));
assign O87iw6 = (~(Twaiw6 | Egfiw6));
assign Oll7v6 = (~(Gx0jy6 & Ox0jy6));
assign Ox0jy6 = (~(Ffj7z6[1] & Iw0jy6));
assign Iw0jy6 = (~(Eu0jy6 & Bqi7z6[0]));
assign Gx0jy6 = (~(Eu0jy6 & Np7iw6));
assign Np7iw6 = (~(Twaiw6 | Gbeiw6));
assign Hll7v6 = (~(Wx0jy6 & Ey0jy6));
assign Ey0jy6 = (~(Zdj7z6[0] & My0jy6));
assign Wx0jy6 = (~(Eu0jy6 & Rl6iw6));
assign Rl6iw6 = (~(Nq6iw6 | Gofiw6));
assign All7v6 = (~(Uy0jy6 & Cz0jy6));
assign Cz0jy6 = (~(Zdj7z6[2] & My0jy6));
assign Uy0jy6 = (~(Eu0jy6 & Hv5iw6));
assign Hv5iw6 = (~(Nq6iw6 | Yqfiw6));
assign Tkl7v6 = (~(Kz0jy6 & Sz0jy6));
assign Sz0jy6 = (~(Zdj7z6[1] & My0jy6));
assign My0jy6 = (~(Eu0jy6 & Bqi7z6[1]));
assign Kz0jy6 = (~(Eu0jy6 & Qa6iw6));
assign Qa6iw6 = (~(Nq6iw6 | Ppfiw6));
assign Nq6iw6 = (!Bqi7z6[1]);
assign Eu0jy6 = (Hvjiw6 & L28iw6);
assign L28iw6 = (~(Wnaiw6 | X22nv6));
assign Mkl7v6 = (A01jy6 ? Doadt6 : U42nv6);
assign Fkl7v6 = (A01jy6 ? O7adt6 : B52nv6);
assign A01jy6 = (!I01jy6);
assign Yjl7v6 = (Q01jy6 ? U42nv6 : Rip7z6[0]);
assign Rjl7v6 = (Q01jy6 ? P52nv6 : Rip7z6[3]);
assign Kjl7v6 = (Q01jy6 ? B52nv6 : Rip7z6[1]);
assign Q01jy6 = (!Y01jy6);
assign Djl7v6 = (G11jy6 ? U42nv6 : G0q7z6[0]);
assign Wil7v6 = (G11jy6 ? P52nv6 : G0q7z6[3]);
assign Pil7v6 = (G11jy6 ? B52nv6 : G0q7z6[1]);
assign Iil7v6 = (O11jy6 ? R62nv6 : W22ft6);
assign Bil7v6 = (O11jy6 ? P52nv6 : I7p7z6[3]);
assign Uhl7v6 = (O11jy6 ? B52nv6 : I7p7z6[1]);
assign Nhl7v6 = (O11jy6 ? U42nv6 : I7p7z6[0]);
assign Ghl7v6 = (O11jy6 ? D62nv6 : M12ft6);
assign Zgl7v6 = (W11jy6 ? U42nv6 : E6p7z6[0]);
assign Sgl7v6 = (W11jy6 ? X0hov6 : E6p7z6[31]);
assign Lgl7v6 = (W11jy6 ? Ro3iw6 : E6p7z6[30]);
assign Egl7v6 = (W11jy6 ? Zz3iw6 : E6p7z6[29]);
assign Xfl7v6 = (W11jy6 ? W14iw6 : E6p7z6[28]);
assign Qfl7v6 = (W11jy6 ? H44iw6 : E6p7z6[27]);
assign Jfl7v6 = (W11jy6 ? E64iw6 : E6p7z6[26]);
assign Cfl7v6 = (W11jy6 ? Iklov6 : E6p7z6[25]);
assign Vel7v6 = (W11jy6 ? Wf4iw6 : E6p7z6[24]);
assign Oel7v6 = (W11jy6 ? Cx4iw6 : E6p7z6[23]);
assign Hel7v6 = (W11jy6 ? D85iw6 : E6p7z6[22]);
assign Ael7v6 = (W11jy6 ? Ej5iw6 : E6p7z6[21]);
assign Tdl7v6 = (W11jy6 ? Bl5iw6 : E6p7z6[20]);
assign Mdl7v6 = (W11jy6 ? Mn5iw6 : E6p7z6[19]);
assign Fdl7v6 = (W11jy6 ? Jp5iw6 : E6p7z6[18]);
assign Ycl7v6 = (W11jy6 ? Gr5iw6 : E6p7z6[17]);
assign Rcl7v6 = (W11jy6 ? Is5iw6 : E6p7z6[16]);
assign Kcl7v6 = (W11jy6 ? Z0iov6 : E6p7z6[15]);
assign Dcl7v6 = (W11jy6 ? Bk6iw6 : E6p7z6[14]);
assign Wbl7v6 = (W11jy6 ? Guhov6 : E6p7z6[13]);
assign Pbl7v6 = (W11jy6 ? Emhov6 : E6p7z6[12]);
assign Ibl7v6 = (W11jy6 ? Dz6iw6 : E6p7z6[11]);
assign Bbl7v6 = (W11jy6 ? H17iw6 : E6p7z6[10]);
assign Ual7v6 = (W11jy6 ? J27iw6 : E6p7z6[9]);
assign Nal7v6 = (W11jy6 ? U47iw6 : E6p7z6[8]);
assign Gal7v6 = (W11jy6 ? R62nv6 : E6p7z6[7]);
assign Z9l7v6 = (W11jy6 ? K62nv6 : E6p7z6[6]);
assign S9l7v6 = (W11jy6 ? D62nv6 : E6p7z6[5]);
assign L9l7v6 = (W11jy6 ? W52nv6 : E6p7z6[4]);
assign E9l7v6 = (W11jy6 ? P52nv6 : E6p7z6[3]);
assign X8l7v6 = (W11jy6 ? B52nv6 : E6p7z6[1]);
assign Q8l7v6 = (E21jy6 ? U42nv6 : Bqp7z6[0]);
assign J8l7v6 = (E21jy6 ? X0hov6 : Bqp7z6[31]);
assign C8l7v6 = (E21jy6 ? Ro3iw6 : Bqp7z6[30]);
assign V7l7v6 = (E21jy6 ? Zz3iw6 : Bqp7z6[29]);
assign O7l7v6 = (E21jy6 ? W14iw6 : Bqp7z6[28]);
assign H7l7v6 = (E21jy6 ? H44iw6 : Bqp7z6[27]);
assign A7l7v6 = (E21jy6 ? E64iw6 : Bqp7z6[26]);
assign T6l7v6 = (E21jy6 ? Iklov6 : Bqp7z6[25]);
assign M6l7v6 = (E21jy6 ? Wf4iw6 : Bqp7z6[24]);
assign F6l7v6 = (E21jy6 ? Cx4iw6 : Bqp7z6[23]);
assign Y5l7v6 = (E21jy6 ? D85iw6 : Bqp7z6[22]);
assign R5l7v6 = (E21jy6 ? Ej5iw6 : Bqp7z6[21]);
assign K5l7v6 = (E21jy6 ? Bl5iw6 : Bqp7z6[20]);
assign D5l7v6 = (E21jy6 ? Mn5iw6 : Bqp7z6[19]);
assign W4l7v6 = (E21jy6 ? Jp5iw6 : Bqp7z6[18]);
assign P4l7v6 = (E21jy6 ? Gr5iw6 : Bqp7z6[17]);
assign I4l7v6 = (E21jy6 ? Is5iw6 : Bqp7z6[16]);
assign B4l7v6 = (E21jy6 ? Z0iov6 : Bqp7z6[15]);
assign U3l7v6 = (E21jy6 ? Bk6iw6 : Bqp7z6[14]);
assign N3l7v6 = (E21jy6 ? Guhov6 : Bqp7z6[13]);
assign G3l7v6 = (E21jy6 ? Emhov6 : Bqp7z6[12]);
assign Z2l7v6 = (E21jy6 ? Dz6iw6 : Bqp7z6[11]);
assign S2l7v6 = (E21jy6 ? H17iw6 : Bqp7z6[10]);
assign L2l7v6 = (E21jy6 ? J27iw6 : Bqp7z6[9]);
assign E2l7v6 = (E21jy6 ? U47iw6 : Bqp7z6[8]);
assign X1l7v6 = (E21jy6 ? R62nv6 : Bqp7z6[7]);
assign Q1l7v6 = (E21jy6 ? K62nv6 : Bqp7z6[6]);
assign J1l7v6 = (E21jy6 ? D62nv6 : Bqp7z6[5]);
assign C1l7v6 = (E21jy6 ? W52nv6 : Bqp7z6[4]);
assign V0l7v6 = (E21jy6 ? P52nv6 : Bqp7z6[3]);
assign O0l7v6 = (E21jy6 ? B52nv6 : Bqp7z6[1]);
assign H0l7v6 = (Etgiw6 ? U42nv6 : Qb4ft6);
assign A0l7v6 = (Etgiw6 ? D85iw6 : Xkq7z6[22]);
assign Tzk7v6 = (Etgiw6 ? Ej5iw6 : Xkq7z6[21]);
assign Mzk7v6 = (Etgiw6 ? Bl5iw6 : Xkq7z6[20]);
assign Fzk7v6 = (Etgiw6 ? Mn5iw6 : Xkq7z6[19]);
assign Yyk7v6 = (Etgiw6 ? Jp5iw6 : Xkq7z6[18]);
assign Ryk7v6 = (Etgiw6 ? Gr5iw6 : Xkq7z6[17]);
assign Kyk7v6 = (Etgiw6 ? Is5iw6 : Xkq7z6[16]);
assign Dyk7v6 = (Etgiw6 ? Z0iov6 : Xkq7z6[15]);
assign Wxk7v6 = (Etgiw6 ? Bk6iw6 : Xkq7z6[14]);
assign Pxk7v6 = (Etgiw6 ? Guhov6 : Xkq7z6[13]);
assign Ixk7v6 = (Etgiw6 ? Emhov6 : Xkq7z6[12]);
assign Bxk7v6 = (Etgiw6 ? Dz6iw6 : W5q7z6[1]);
assign Uwk7v6 = (Etgiw6 ? H17iw6 : W5q7z6[0]);
assign Nwk7v6 = (Etgiw6 ? J27iw6 : Id4ft6);
assign Gwk7v6 = (Etgiw6 ? U47iw6 : X9q7z6[3]);
assign Zvk7v6 = (Etgiw6 ? R62nv6 : X9q7z6[2]);
assign Svk7v6 = (Etgiw6 ? K62nv6 : X9q7z6[1]);
assign Lvk7v6 = (Etgiw6 ? D62nv6 : X9q7z6[0]);
assign Evk7v6 = (Etgiw6 ? W52nv6 : Y7q7z6[3]);
assign Xuk7v6 = (Etgiw6 ? P52nv6 : Y7q7z6[2]);
assign Quk7v6 = (Etgiw6 ? B52nv6 : Y7q7z6[0]);
assign Juk7v6 = (M21jy6 ? D62nv6 : Dm2ft6);
assign Cuk7v6 = (M21jy6 ? P52nv6 : Hmp7z6[3]);
assign Vtk7v6 = (M21jy6 ? B52nv6 : Hmp7z6[1]);
assign Otk7v6 = (M21jy6 ? U42nv6 : Hmp7z6[0]);
assign Htk7v6 = (U21jy6 ? U42nv6 : Q8p7z6[0]);
assign Atk7v6 = (U21jy6 ? P52nv6 : Q8p7z6[3]);
assign Tsk7v6 = (U21jy6 ? B52nv6 : Q8p7z6[1]);
assign U21jy6 = (!C31jy6);
assign Msk7v6 = (K31jy6 ? U42nv6 : Gop7z6[0]);
assign Fsk7v6 = (K31jy6 ? P52nv6 : Gop7z6[3]);
assign Yrk7v6 = (K31jy6 ? B52nv6 : Gop7z6[1]);
assign Rrk7v6 = (S31jy6 ? D62nv6 : Ei2ft6);
assign Krk7v6 = (S31jy6 ? P52nv6 : Sgp7z6[3]);
assign Drk7v6 = (S31jy6 ? B52nv6 : Sgp7z6[1]);
assign Wqk7v6 = (S31jy6 ? U42nv6 : Sgp7z6[0]);
assign Pqk7v6 = (A41jy6 ? U42nv6 : B2q7z6[0]);
assign Iqk7v6 = (A41jy6 ? X0hov6 : B2q7z6[31]);
assign Bqk7v6 = (A41jy6 ? Ro3iw6 : B2q7z6[30]);
assign Upk7v6 = (A41jy6 ? Zz3iw6 : B2q7z6[29]);
assign Npk7v6 = (A41jy6 ? W14iw6 : B2q7z6[28]);
assign Gpk7v6 = (A41jy6 ? H44iw6 : B2q7z6[27]);
assign Zok7v6 = (A41jy6 ? E64iw6 : B2q7z6[26]);
assign Sok7v6 = (A41jy6 ? Iklov6 : B2q7z6[25]);
assign Lok7v6 = (A41jy6 ? Wf4iw6 : B2q7z6[24]);
assign Eok7v6 = (A41jy6 ? Cx4iw6 : B2q7z6[23]);
assign Xnk7v6 = (A41jy6 ? D85iw6 : B2q7z6[22]);
assign Qnk7v6 = (A41jy6 ? Ej5iw6 : B2q7z6[21]);
assign Jnk7v6 = (A41jy6 ? Bl5iw6 : B2q7z6[20]);
assign Cnk7v6 = (A41jy6 ? Mn5iw6 : B2q7z6[19]);
assign Vmk7v6 = (A41jy6 ? Jp5iw6 : B2q7z6[18]);
assign Omk7v6 = (A41jy6 ? Gr5iw6 : B2q7z6[17]);
assign Hmk7v6 = (A41jy6 ? Is5iw6 : B2q7z6[16]);
assign Amk7v6 = (A41jy6 ? Z0iov6 : B2q7z6[15]);
assign Tlk7v6 = (A41jy6 ? Bk6iw6 : B2q7z6[14]);
assign Mlk7v6 = (A41jy6 ? Guhov6 : B2q7z6[13]);
assign Flk7v6 = (A41jy6 ? Emhov6 : B2q7z6[12]);
assign Ykk7v6 = (A41jy6 ? Dz6iw6 : B2q7z6[11]);
assign Rkk7v6 = (A41jy6 ? H17iw6 : B2q7z6[10]);
assign Kkk7v6 = (A41jy6 ? J27iw6 : B2q7z6[9]);
assign Dkk7v6 = (A41jy6 ? U47iw6 : B2q7z6[8]);
assign Wjk7v6 = (A41jy6 ? R62nv6 : B2q7z6[7]);
assign Pjk7v6 = (A41jy6 ? K62nv6 : B2q7z6[6]);
assign Ijk7v6 = (A41jy6 ? D62nv6 : B2q7z6[5]);
assign Bjk7v6 = (A41jy6 ? W52nv6 : B2q7z6[4]);
assign Uik7v6 = (A41jy6 ? P52nv6 : B2q7z6[3]);
assign Nik7v6 = (A41jy6 ? B52nv6 : B2q7z6[1]);
assign Gik7v6 = (I41jy6 ? B52nv6 : Mkp7z6[1]);
assign Zhk7v6 = (I41jy6 ? P52nv6 : Mkp7z6[3]);
assign Shk7v6 = (I41jy6 ? W52nv6 : Mkp7z6[4]);
assign Lhk7v6 = (I41jy6 ? D62nv6 : Mkp7z6[5]);
assign Ehk7v6 = (I41jy6 ? K62nv6 : Mkp7z6[6]);
assign Xgk7v6 = (I41jy6 ? R62nv6 : Mkp7z6[7]);
assign Qgk7v6 = (I41jy6 ? U47iw6 : Mkp7z6[8]);
assign Jgk7v6 = (I41jy6 ? J27iw6 : Mkp7z6[9]);
assign Cgk7v6 = (I41jy6 ? H17iw6 : Mkp7z6[10]);
assign Vfk7v6 = (I41jy6 ? Dz6iw6 : Mkp7z6[11]);
assign Ofk7v6 = (I41jy6 ? Emhov6 : Mkp7z6[12]);
assign Hfk7v6 = (I41jy6 ? Guhov6 : Mkp7z6[13]);
assign Afk7v6 = (I41jy6 ? Bk6iw6 : Mkp7z6[14]);
assign Tek7v6 = (I41jy6 ? Z0iov6 : Mkp7z6[15]);
assign Mek7v6 = (I41jy6 ? Is5iw6 : Mkp7z6[16]);
assign Fek7v6 = (I41jy6 ? Gr5iw6 : Mkp7z6[17]);
assign Ydk7v6 = (I41jy6 ? Jp5iw6 : Mkp7z6[18]);
assign Rdk7v6 = (I41jy6 ? Mn5iw6 : Mkp7z6[19]);
assign Kdk7v6 = (I41jy6 ? Bl5iw6 : Mkp7z6[20]);
assign Ddk7v6 = (I41jy6 ? Ej5iw6 : Mkp7z6[21]);
assign Wck7v6 = (I41jy6 ? D85iw6 : Mkp7z6[22]);
assign Pck7v6 = (I41jy6 ? Cx4iw6 : Mkp7z6[23]);
assign Ick7v6 = (I41jy6 ? Wf4iw6 : Mkp7z6[24]);
assign Bck7v6 = (I41jy6 ? Iklov6 : Mkp7z6[25]);
assign Ubk7v6 = (I41jy6 ? E64iw6 : Mkp7z6[26]);
assign Nbk7v6 = (I41jy6 ? H44iw6 : Mkp7z6[27]);
assign Gbk7v6 = (I41jy6 ? W14iw6 : Mkp7z6[28]);
assign Zak7v6 = (I41jy6 ? Zz3iw6 : Mkp7z6[29]);
assign Sak7v6 = (I41jy6 ? Ro3iw6 : Mkp7z6[30]);
assign Lak7v6 = (I41jy6 ? X0hov6 : Mkp7z6[31]);
assign Eak7v6 = (I41jy6 ? U42nv6 : Mkp7z6[0]);
assign X9k7v6 = (Q41jy6 ? D62nv6 : Gs2ft6);
assign Q9k7v6 = (Q41jy6 ? P52nv6 : Hyp7z6[3]);
assign J9k7v6 = (Q41jy6 ? B52nv6 : Hyp7z6[1]);
assign C9k7v6 = (Q41jy6 ? U42nv6 : Hyp7z6[0]);
assign V8k7v6 = (Q41jy6 ? Dz6iw6 : Gwp7z6[1]);
assign O8k7v6 = (Q41jy6 ? Emhov6 : Bup7z6[0]);
assign H8k7v6 = (Q41jy6 ? Guhov6 : Bup7z6[1]);
assign A8k7v6 = (Q41jy6 ? Is5iw6 : Wrp7z6[0]);
assign T7k7v6 = (Q41jy6 ? Gr5iw6 : Wrp7z6[1]);
assign M7k7v6 = (Q41jy6 ? U47iw6 : Cq2ft6);
assign F7k7v6 = (Q41jy6 ? H17iw6 : Gwp7z6[0]);
assign Y6k7v6 = (Otshy6 ? Xfymz6[2] : Pjb7z6[2]);
assign Otshy6 = (!Mphiw6);
assign Mphiw6 = (Y41jy6 & G51jy6);
assign Y41jy6 = (O51jy6 & W51jy6);
assign W51jy6 = (~(E61jy6 | Pjb7z6[13]));
assign O51jy6 = (Pjb7z6[18] & Pjb7z6[12]);
assign R6k7v6 = (M61jy6 ? Z0iov6 : Unymz6[9]);
assign K6k7v6 = (M61jy6 ? R62nv6 : Unymz6[4]);
assign D6k7v6 = (M61jy6 ? Emhov6 : Unymz6[6]);
assign W5k7v6 = (M61jy6 ? Guhov6 : Unymz6[7]);
assign P5k7v6 = (M61jy6 ? U42nv6 : Unymz6[0]);
assign I5k7v6 = (M61jy6 ? B52nv6 : Unymz6[1]);
assign B5k7v6 = (M61jy6 ? D62nv6 : Unymz6[2]);
assign U4k7v6 = (M61jy6 ? K62nv6 : Unymz6[3]);
assign N4k7v6 = (M61jy6 ? Bk6iw6 : Unymz6[8]);
assign G4k7v6 = (U61jy6 ? Z0iov6 : Ojymz6[9]);
assign Z3k7v6 = (U61jy6 ? R62nv6 : Ojymz6[4]);
assign S3k7v6 = (U61jy6 ? Emhov6 : Ojymz6[6]);
assign L3k7v6 = (U61jy6 ? Guhov6 : Ojymz6[7]);
assign E3k7v6 = (U61jy6 ? U42nv6 : Ojymz6[0]);
assign X2k7v6 = (U61jy6 ? B52nv6 : Ojymz6[1]);
assign Q2k7v6 = (U61jy6 ? D62nv6 : Ojymz6[2]);
assign J2k7v6 = (U61jy6 ? K62nv6 : Ojymz6[3]);
assign C2k7v6 = (U61jy6 ? Bk6iw6 : Ojymz6[8]);
assign V1k7v6 = (C71jy6 ? B52nv6 : Kmymz6[1]);
assign O1k7v6 = (C71jy6 ? P52nv6 : Kmymz6[3]);
assign H1k7v6 = (C71jy6 ? Gr5iw6 : Blymz6[1]);
assign A1k7v6 = (C71jy6 ? Jp5iw6 : Blymz6[2]);
assign T0k7v6 = (C71jy6 ? Mn5iw6 : Blymz6[3]);
assign M0k7v6 = (C71jy6 ? U42nv6 : Kmymz6[0]);
assign F0k7v6 = (K71jy6 ? U42nv6 : At67v6);
assign K71jy6 = (S71jy6 & Xid8x6);
assign S71jy6 = (A81jy6 & L9pyx6);
assign L9pyx6 = (~(I81jy6 | Opniy6));
assign Opniy6 = (~(Q81jy6 & Xfymz6[9]));
assign Q81jy6 = (Xfymz6[11] & Xfymz6[10]);
assign Yzj7v6 = (Y81jy6 ? B52nv6 : Wd77z6);
assign Rzj7v6 = (Y81jy6 ? P52nv6 : Cf77z6);
assign Kzj7v6 = (Y81jy6 ? W52nv6 : Kf77z6);
assign Dzj7v6 = (Y81jy6 ? D62nv6 : Sf77z6);
assign Wyj7v6 = (Y81jy6 ? K62nv6 : Ag77z6);
assign Pyj7v6 = (Y81jy6 ? U42nv6 : Gh77z6);
assign Iyj7v6 = (G91jy6 ? B52nv6 : Biymz6[1]);
assign Byj7v6 = (G91jy6 ? P52nv6 : Biymz6[3]);
assign Uxj7v6 = (G91jy6 ? W52nv6 : Biymz6[4]);
assign Nxj7v6 = (G91jy6 ? D62nv6 : Biymz6[5]);
assign Gxj7v6 = (G91jy6 ? K62nv6 : Biymz6[6]);
assign Zwj7v6 = (G91jy6 ? R62nv6 : Biymz6[7]);
assign Swj7v6 = (G91jy6 ? J27iw6 : Biymz6[9]);
assign Lwj7v6 = (G91jy6 ? H17iw6 : Biymz6[10]);
assign Ewj7v6 = (G91jy6 ? Dz6iw6 : Biymz6[11]);
assign Xvj7v6 = (G91jy6 ? Emhov6 : Biymz6[12]);
assign Qvj7v6 = (G91jy6 ? Guhov6 : Biymz6[13]);
assign Jvj7v6 = (G91jy6 ? Bk6iw6 : Biymz6[14]);
assign Cvj7v6 = (G91jy6 ? Z0iov6 : Biymz6[15]);
assign Vuj7v6 = (G91jy6 ? U42nv6 : Biymz6[0]);
assign Ouj7v6 = (O91jy6 ? W52nv6 : Feymz6[0]);
assign Huj7v6 = (O91jy6 ? D62nv6 : Feymz6[1]);
assign Auj7v6 = (O91jy6 ? K62nv6 : Feymz6[2]);
assign Ttj7v6 = (O91jy6 ? Ej5iw6 : Feymz6[3]);
assign Mtj7v6 = (O91jy6 ? Gr5iw6 : Bfymz6[1]);
assign Ftj7v6 = (O91jy6 ? Guhov6 : Bfymz6[2]);
assign Ysj7v6 = (O91jy6 ? Dz6iw6 : Ue77z6);
assign Rsj7v6 = (O91jy6 ? H17iw6 : C477v6);
assign Ksj7v6 = (O91jy6 ? J27iw6 : W177v6);
assign Dsj7v6 = (O91jy6 ? R62nv6 : Vv67v6);
assign Wrj7v6 = (O91jy6 ? U42nv6 : Wy67v6);
assign Prj7v6 = (Lhliw6 ? Tjr7z6[6] : ETMINTNUM[4]);
assign Irj7v6 = (Lhliw6 ? Tjr7z6[10] : ETMINTNUM[8]);
assign Brj7v6 = (O91jy6 ? W14iw6 : Xz67v6);
assign Uqj7v6 = (R1snv6 ? Gnzmz6[0] : TSVALUEB[0]);
assign Nqj7v6 = (R1snv6 ? Ync7v6 : TSVALUEB[47]);
assign Gqj7v6 = (R1snv6 ? Emc7v6 : TSVALUEB[46]);
assign Zpj7v6 = (R1snv6 ? Kkc7v6 : TSVALUEB[45]);
assign Spj7v6 = (R1snv6 ? Qic7v6 : TSVALUEB[44]);
assign Lpj7v6 = (R1snv6 ? Wgc7v6 : TSVALUEB[43]);
assign Epj7v6 = (R1snv6 ? Cfc7v6 : TSVALUEB[42]);
assign Xoj7v6 = (R1snv6 ? Gnzmz6[46] : TSVALUEB[41]);
assign Qoj7v6 = (R1snv6 ? Gnzmz6[45] : TSVALUEB[40]);
assign Joj7v6 = (R1snv6 ? Gnzmz6[44] : TSVALUEB[39]);
assign Coj7v6 = (R1snv6 ? Gnzmz6[43] : TSVALUEB[38]);
assign Vnj7v6 = (R1snv6 ? Gnzmz6[42] : TSVALUEB[37]);
assign Onj7v6 = (R1snv6 ? Gnzmz6[41] : TSVALUEB[36]);
assign Hnj7v6 = (R1snv6 ? Gnzmz6[40] : TSVALUEB[35]);
assign Anj7v6 = (R1snv6 ? Gnzmz6[38] : TSVALUEB[34]);
assign Tmj7v6 = (R1snv6 ? Gnzmz6[37] : TSVALUEB[33]);
assign Mmj7v6 = (R1snv6 ? Gnzmz6[36] : TSVALUEB[32]);
assign Fmj7v6 = (R1snv6 ? Gnzmz6[35] : TSVALUEB[31]);
assign Ylj7v6 = (R1snv6 ? Gnzmz6[34] : TSVALUEB[30]);
assign Rlj7v6 = (R1snv6 ? Gnzmz6[33] : TSVALUEB[29]);
assign Klj7v6 = (R1snv6 ? Gnzmz6[32] : TSVALUEB[28]);
assign Dlj7v6 = (R1snv6 ? Gnzmz6[30] : TSVALUEB[27]);
assign Wkj7v6 = (R1snv6 ? Gnzmz6[29] : TSVALUEB[26]);
assign Pkj7v6 = (R1snv6 ? Gnzmz6[28] : TSVALUEB[25]);
assign Ikj7v6 = (R1snv6 ? Gnzmz6[27] : TSVALUEB[24]);
assign Bkj7v6 = (R1snv6 ? Gnzmz6[26] : TSVALUEB[23]);
assign Ujj7v6 = (R1snv6 ? Gnzmz6[25] : TSVALUEB[22]);
assign Njj7v6 = (R1snv6 ? Gnzmz6[24] : TSVALUEB[21]);
assign Gjj7v6 = (R1snv6 ? Gnzmz6[22] : TSVALUEB[20]);
assign Zij7v6 = (R1snv6 ? Gnzmz6[21] : TSVALUEB[19]);
assign Sij7v6 = (R1snv6 ? Gnzmz6[20] : TSVALUEB[18]);
assign Lij7v6 = (R1snv6 ? Gnzmz6[19] : TSVALUEB[17]);
assign Eij7v6 = (R1snv6 ? Gnzmz6[18] : TSVALUEB[16]);
assign Xhj7v6 = (R1snv6 ? Gnzmz6[17] : TSVALUEB[15]);
assign Qhj7v6 = (R1snv6 ? Gnzmz6[16] : TSVALUEB[14]);
assign Jhj7v6 = (R1snv6 ? Gnzmz6[14] : TSVALUEB[13]);
assign Chj7v6 = (R1snv6 ? Gnzmz6[13] : TSVALUEB[12]);
assign Vgj7v6 = (R1snv6 ? Gnzmz6[12] : TSVALUEB[11]);
assign Ogj7v6 = (R1snv6 ? Gnzmz6[11] : TSVALUEB[10]);
assign Hgj7v6 = (R1snv6 ? Gnzmz6[10] : TSVALUEB[9]);
assign Agj7v6 = (R1snv6 ? Gnzmz6[9] : TSVALUEB[8]);
assign Tfj7v6 = (R1snv6 ? Gnzmz6[8] : TSVALUEB[7]);
assign Mfj7v6 = (R1snv6 ? Gnzmz6[6] : TSVALUEB[6]);
assign Ffj7v6 = (R1snv6 ? Gnzmz6[5] : TSVALUEB[5]);
assign Yej7v6 = (R1snv6 ? Gnzmz6[4] : TSVALUEB[4]);
assign Rej7v6 = (R1snv6 ? Gnzmz6[3] : TSVALUEB[3]);
assign Kej7v6 = (R1snv6 ? Gnzmz6[2] : TSVALUEB[2]);
assign R1snv6 = (!W91jy6);
assign Dej7v6 = (W91jy6 ? TSVALUEB[1] : Gnzmz6[1]);
assign W91jy6 = (Ea1jy6 & Ma1jy6);
assign Ma1jy6 = (Fgzmz6[0] & Xz67v6);
assign Ea1jy6 = (Hqb7v6 & G197z6);
assign Wdj7v6 = (Ua1jy6 ? Z0iov6 : Sgymz6[9]);
assign Pdj7v6 = (Ua1jy6 ? R62nv6 : Sgymz6[4]);
assign Idj7v6 = (Ua1jy6 ? Emhov6 : Sgymz6[6]);
assign Bdj7v6 = (Ua1jy6 ? Guhov6 : Sgymz6[7]);
assign Ucj7v6 = (Ua1jy6 ? U42nv6 : Sgymz6[0]);
assign Ncj7v6 = (Ua1jy6 ? B52nv6 : Sgymz6[1]);
assign Gcj7v6 = (Ua1jy6 ? D62nv6 : Sgymz6[2]);
assign Zbj7v6 = (Ua1jy6 ? K62nv6 : Sgymz6[3]);
assign Sbj7v6 = (Ua1jy6 ? Bk6iw6 : Sgymz6[8]);
assign Lbj7v6 = (Cb1jy6 ? Iklov6 : Ok77v6);
assign Cb1jy6 = (Sz8iy6 & Xid8x6);
assign Sz8iy6 = (Kb1jy6 & J2xyx6);
assign J2xyx6 = (Sb1jy6 & Xfymz6[2]);
assign Sb1jy6 = (Eyyhy6 & J6yyx6);
assign Ebj7v6 = (Qgnhy6 ? J02nz6[2] : Pjb7z6[2]);
assign Qgnhy6 = (!Kniiw6);
assign Kniiw6 = (Ac1jy6 & G51jy6);
assign G51jy6 = (Ic1jy6 & Qc1jy6);
assign Qc1jy6 = (Yc1jy6 & Crhiw6);
assign Crhiw6 = (!Pjb7z6[16]);
assign Yc1jy6 = (~(Pjb7z6[17] | Pjb7z6[19]));
assign Ic1jy6 = (~(Pjb7z6[14] | Pjb7z6[15]));
assign Ac1jy6 = (Gd1jy6 & Od1jy6);
assign Od1jy6 = (~(Pjb7z6[12] | Pjb7z6[13]));
assign Gd1jy6 = (Pjb7z6[18] & Wd1jy6);
assign Xaj7v6 = (Cjliy6 ? Pjb7z6[2] : Ti2nz6[0]);
assign Cjliy6 = (!Maziy6);
assign Maziy6 = (Oduhy6 | W2adt6);
assign Oduhy6 = (~(Ee1jy6 & Me1jy6));
assign Me1jy6 = (Ue1jy6 & Cf1jy6);
assign Cf1jy6 = (Kf1jy6 & Pjb7z6[13]);
assign Kf1jy6 = (Pjb7z6[12] & Wd1jy6);
assign Wd1jy6 = (!E61jy6);
assign E61jy6 = (~(D16ft6 | K2adt6));
assign Ue1jy6 = (Pjb7z6[15] & Pjb7z6[14]);
assign Ee1jy6 = (Sf1jy6 & Ag1jy6);
assign Ag1jy6 = (Pjb7z6[17] & Pjb7z6[16]);
assign Sf1jy6 = (Pjb7z6[19] & Pjb7z6[18]);
assign Qaj7v6 = (Ig1jy6 ? Eshiw6 : L1syx6);
assign Ig1jy6 = (Qg1jy6 & Yg1jy6);
assign Yg1jy6 = (Gh1jy6 & Oh1jy6);
assign Oh1jy6 = (~(Vpd7x6 | C397z6));
assign Vpd7x6 = (!Ihs7z6[0]);
assign Gh1jy6 = (Ihs7z6[2] & Ihs7z6[1]);
assign Qg1jy6 = (Wh1jy6 & Ei1jy6);
assign Wh1jy6 = (Llryx6 & Ihs7z6[3]);
assign Eshiw6 = (~(Mi1jy6 & Ui1jy6));
assign Ui1jy6 = (Cj1jy6 & Kj1jy6);
assign Kj1jy6 = (Sj1jy6 & Ak1jy6);
assign Ak1jy6 = (Ik1jy6 & W52nv6);
assign Ik1jy6 = (H17iw6 & Dz6iw6);
assign Sj1jy6 = (X0hov6 & Jp5iw6);
assign Cj1jy6 = (Qk1jy6 & Yk1jy6);
assign Yk1jy6 = (J27iw6 & K62nv6);
assign Qk1jy6 = (Z0iov6 & Ro3iw6);
assign Mi1jy6 = (Gl1jy6 & Ol1jy6);
assign Ol1jy6 = (Wl1jy6 & Em1jy6);
assign Em1jy6 = (Mm1jy6 & Kxfiw6);
assign Mm1jy6 = (Gofiw6 & Bk6iw6);
assign Wl1jy6 = (Nhfiw6 & Oyhov6);
assign Gl1jy6 = (Um1jy6 & Cn1jy6);
assign Cn1jy6 = (N5m7x6 & Umhiw6);
assign N5m7x6 = (Kn1jy6 & Sn1jy6);
assign Sn1jy6 = (Ao1jy6 & Io1jy6);
assign Io1jy6 = (Qo1jy6 & Wf4iw6);
assign Qo1jy6 = (Cx4iw6 & Ej5iw6);
assign Ao1jy6 = (Mn5iw6 & E64iw6);
assign Kn1jy6 = (Yo1jy6 & Gp1jy6);
assign Yo1jy6 = (N9giw6 & Hsfiw6);
assign Um1jy6 = (Ucdiw6 & Nbeiw6);
assign Nbeiw6 = (Op1jy6 & Tdfiw6);
assign Op1jy6 = (Egfiw6 & Pohov6);
assign Ucdiw6 = (Wp1jy6 & L19iw6);
assign L19iw6 = (!B52nv6);
assign Wp1jy6 = (U42nv6 & I52nv6);
assign Jaj7v6 = (Eq1jy6 ? U42nv6 : Ig27v6);
assign Eq1jy6 = (Foryx6 & Mq1jy6);
assign Foryx6 = (Uq1jy6 & Cr1jy6);
assign Cr1jy6 = (Tt4yx6 & Pfryx6);
assign Uq1jy6 = (Ei1jy6 & Xruyx6);
assign Ei1jy6 = (Kr1jy6 & Zfs7z6[8]);
assign Kr1jy6 = (P7wyx6 & D1syx6);
assign Caj7v6 = (Sr1jy6 ? U42nv6 : Ln6ft6);
assign Sr1jy6 = (As1jy6 & Is1jy6);
assign Is1jy6 = (Qs1jy6 & Mq1jy6);
assign Qs1jy6 = (L51zx6 & Fgryx6);
assign L51zx6 = (!Or27v6);
assign As1jy6 = (Ys1jy6 & Llryx6);
assign Llryx6 = (Gt1jy6 & Ap27v6);
assign Gt1jy6 = (Tn27v6 & Zfs7z6[7]);
assign Ys1jy6 = (~(Pruyx6 | D1syx6));
assign D1syx6 = (!Mm27v6);
assign Pruyx6 = (~(Ot1jy6 & Wt1jy6));
assign Wt1jy6 = (Zfs7z6[11] & Zfs7z6[10]);
assign Ot1jy6 = (Hq27v6 & Zfs7z6[9]);
assign V9j7v6 = (Hr4yx6 ? Gr5iw6 : Mqb7z6[1]);
assign O9j7v6 = (Hr4yx6 ? Jp5iw6 : Mqb7z6[2]);
assign H9j7v6 = (Hr4yx6 ? Mn5iw6 : Mqb7z6[3]);
assign A9j7v6 = (Hr4yx6 ? Bl5iw6 : Mqb7z6[4]);
assign T8j7v6 = (Hr4yx6 ? Ej5iw6 : Mqb7z6[5]);
assign M8j7v6 = (Hr4yx6 ? D85iw6 : Mqb7z6[6]);
assign F8j7v6 = (Hr4yx6 ? U42nv6 : Rj27v6);
assign Y7j7v6 = (Hr4yx6 ? B52nv6 : Ci6ft6);
assign R7j7v6 = (Hr4yx6 ? P52nv6 : D86ft6);
assign K7j7v6 = (Hr4yx6 ? W52nv6 : Og6ft6);
assign D7j7v6 = (Hr4yx6 ? J27iw6 : Zm37v6);
assign W6j7v6 = (Hr4yx6 ? H17iw6 : R8s7z6[0]);
assign P6j7v6 = (Hr4yx6 ? Dz6iw6 : R8s7z6[1]);
assign I6j7v6 = (Eu1jy6 ? B52nv6 : Scs7z6[1]);
assign B6j7v6 = (Eu1jy6 ? P52nv6 : Scs7z6[3]);
assign U5j7v6 = (Eu1jy6 ? U42nv6 : Scs7z6[0]);
assign N5j7v6 = (Mu1jy6 ? Wf4iw6 : Ies7z6[24]);
assign G5j7v6 = (Mu1jy6 ? X0hov6 : Ies7z6[31]);
assign Z4j7v6 = (Mu1jy6 ? Ro3iw6 : Ies7z6[30]);
assign S4j7v6 = (Mu1jy6 ? Zz3iw6 : Ies7z6[29]);
assign L4j7v6 = (Mu1jy6 ? W14iw6 : Ies7z6[28]);
assign E4j7v6 = (Mu1jy6 ? H44iw6 : Ies7z6[27]);
assign X3j7v6 = (Mu1jy6 ? E64iw6 : Ies7z6[26]);
assign Q3j7v6 = (Mu1jy6 ? Iklov6 : Ies7z6[25]);
assign Mu1jy6 = (Uu1jy6 & Cv1jy6);
assign Uu1jy6 = (Ihs7z6[3] & Kv1jy6);
assign Kv1jy6 = (~(C397z6 & Scs7z6[3]));
assign J3j7v6 = (Sv1jy6 ? Z0iov6 : Ies7z6[15]);
assign C3j7v6 = (Sv1jy6 ? Bk6iw6 : Ies7z6[14]);
assign V2j7v6 = (Sv1jy6 ? Guhov6 : Ies7z6[13]);
assign O2j7v6 = (Sv1jy6 ? Emhov6 : Ies7z6[12]);
assign H2j7v6 = (Sv1jy6 ? Dz6iw6 : Ies7z6[11]);
assign A2j7v6 = (Sv1jy6 ? H17iw6 : Ies7z6[10]);
assign T1j7v6 = (Sv1jy6 ? J27iw6 : Ies7z6[9]);
assign M1j7v6 = (Aw1jy6 ? U42nv6 : Ies7z6[0]);
assign F1j7v6 = (Aw1jy6 ? R62nv6 : Ies7z6[7]);
assign Y0j7v6 = (Aw1jy6 ? K62nv6 : Ies7z6[6]);
assign R0j7v6 = (Aw1jy6 ? D62nv6 : Ies7z6[5]);
assign K0j7v6 = (Aw1jy6 ? W52nv6 : Ies7z6[4]);
assign D0j7v6 = (Aw1jy6 ? P52nv6 : Ies7z6[3]);
assign Wzi7v6 = (Aw1jy6 ? B52nv6 : Ies7z6[1]);
assign Pzi7v6 = (Etgiw6 ? I52nv6 : Y7q7z6[1]);
assign Etgiw6 = (Jsgiw6 & B6qyx6);
assign B6qyx6 = (Iw1jy6 & Z6tyx6);
assign Izi7v6 = (E21jy6 ? I52nv6 : Bqp7z6[2]);
assign E21jy6 = (Jsgiw6 & D5qyx6);
assign D5qyx6 = (~(Qw1jy6 | Ghlhy6));
assign Bzi7v6 = (K31jy6 ? I52nv6 : Gop7z6[2]);
assign K31jy6 = (Jsgiw6 & Z6qyx6);
assign Z6qyx6 = (~(Qw1jy6 | Yglhy6));
assign Uyi7v6 = (Y01jy6 ? Rip7z6[2] : I52nv6);
assign Y01jy6 = (~(Jsgiw6 & H7qyx6));
assign H7qyx6 = (Yw1jy6 & Qcjhy6);
assign Yw1jy6 = (!Qw1jy6);
assign Nyi7v6 = (M21jy6 ? I52nv6 : Hmp7z6[2]);
assign M21jy6 = (Jsgiw6 & P3a8x6);
assign P3a8x6 = (Gx1jy6 & Ox1jy6);
assign Ox1jy6 = (Z6tyx6 & Xueiw6);
assign Gx1jy6 = (Nmq7z6[6] & Hbvyx6);
assign Gyi7v6 = (S31jy6 ? I52nv6 : Sgp7z6[2]);
assign S31jy6 = (Jsgiw6 & Ua9ov6);
assign Ua9ov6 = (Wx1jy6 & Ey1jy6);
assign Ey1jy6 = (Hbvyx6 & Xueiw6);
assign Hbvyx6 = (Nmq7z6[3] & My1jy6);
assign Wx1jy6 = (Nmq7z6[6] & B2qyx6);
assign Zxi7v6 = (W11jy6 ? I52nv6 : E6p7z6[2]);
assign W11jy6 = (Jsgiw6 & L9qyx6);
assign L9qyx6 = (~(Uy1jy6 | Ghlhy6));
assign Ghlhy6 = (!Z6tyx6);
assign Sxi7v6 = (C31jy6 ? Q8p7z6[2] : I52nv6);
assign C31jy6 = (~(Jsgiw6 & Xbqyx6));
assign Xbqyx6 = (Cz1jy6 & Vcyyx6);
assign Cz1jy6 = (!Uy1jy6);
assign Lxi7v6 = (A41jy6 ? I52nv6 : B2q7z6[2]);
assign A41jy6 = (Jsgiw6 & Fcqyx6);
assign Fcqyx6 = (~(Uy1jy6 | Wdlhy6));
assign Exi7v6 = (G11jy6 ? I52nv6 : G0q7z6[2]);
assign G11jy6 = (Jsgiw6 & Zaqyx6);
assign Zaqyx6 = (~(Uy1jy6 | Kflhy6));
assign Kflhy6 = (!Qcjhy6);
assign Qcjhy6 = (~(Kz1jy6 | E297z6));
assign Uy1jy6 = (~(Gllhy6 & Gpeiy6));
assign Gllhy6 = (Nmq7z6[5] & Sz1jy6);
assign Xwi7v6 = (O11jy6 ? I52nv6 : I7p7z6[2]);
assign O11jy6 = (Jsgiw6 & Nao7x6);
assign Nao7x6 = (A02jy6 & Z6tyx6);
assign Z6tyx6 = (~(Bxeiw6 | Nmq7z6[4]));
assign A02jy6 = (!I02jy6);
assign Qwi7v6 = (Q41jy6 ? I52nv6 : Hyp7z6[2]);
assign Q41jy6 = (Jsgiw6 & Q0a8x6);
assign Q0a8x6 = (~(I02jy6 | Wdlhy6));
assign I02jy6 = (~(Q02jy6 & Gpeiy6));
assign Q02jy6 = (Nmq7z6[5] & Nmq7z6[3]);
assign Jwi7v6 = (I41jy6 ? I52nv6 : Mkp7z6[2]);
assign I41jy6 = (Jsgiw6 & Tdqyx6);
assign Tdqyx6 = (~(Qw1jy6 | Wdlhy6));
assign Wdlhy6 = (!B2qyx6);
assign B2qyx6 = (~(Bxeiw6 | Kz1jy6));
assign Kz1jy6 = (!Nmq7z6[4]);
assign Bxeiw6 = (!E297z6);
assign Qw1jy6 = (~(Y02jy6 & G12jy6));
assign G12jy6 = (My1jy6 & Xueiw6);
assign Y02jy6 = (Nmq7z6[6] & Sz1jy6);
assign Cwi7v6 = (Zhg7x6 ? I52nv6 : Ayeet6);
assign Zhg7x6 = (O12jy6 & W12jy6);
assign W12jy6 = (E22jy6 & M22jy6);
assign M22jy6 = (U22jy6 & Gr5iw6);
assign U22jy6 = (Jp5iw6 & Is5iw6);
assign E22jy6 = (X0hov6 & Bl5iw6);
assign O12jy6 = (C32jy6 & K32jy6);
assign K32jy6 = (S32jy6 & N42nv6);
assign N42nv6 = (A42jy6 & I42jy6);
assign A42jy6 = (~(G92iw6 | Ej5iw6));
assign G92iw6 = (~(Pb8iw6 & Wnaiw6));
assign S32jy6 = (Q42jy6 & Mn5iw6);
assign C32jy6 = (Hq3iw6 & Zy4iw6);
assign Zy4iw6 = (~(Ie5iw6 | C0giw6));
assign Hq3iw6 = (~(Dv3iw6 | N9giw6));
assign Dv3iw6 = (!Bqi7z6[3]);
assign Vvi7v6 = (Knniy6 ? I52nv6 : Qij7z6[2]);
assign Knniy6 = (Y42jy6 & G52jy6);
assign G52jy6 = (O52jy6 & W52jy6);
assign W52jy6 = (F02nv6 & Wnaiw6);
assign F02nv6 = (!Ldo7v6);
assign O52jy6 = (Kdadt6 & Q42jy6);
assign Q42jy6 = (E62jy6 & Bqi7z6[1]);
assign E62jy6 = (~(Twaiw6 | N92iw6));
assign Y42jy6 = (M62jy6 & Bqi7z6[3]);
assign M62jy6 = (Bqi7z6[2] & Toi7z6[2]);
assign Ovi7v6 = (M20jy6 ? U3cet6 : I52nv6);
assign M20jy6 = (~(Hvjiw6 & Zh18x6));
assign Hvjiw6 = (U62jy6 & Pi8iw6);
assign U62jy6 = (G42nv6 & Pb8iw6);
assign Hvi7v6 = (I01jy6 ? I52nv6 : Dpadt6);
assign I01jy6 = (C72jy6 & Doaiw6);
assign C72jy6 = (T68iw6 & Bqi7z6[0]);
assign T68iw6 = (~(Wnaiw6 | Toi7z6[4]));
assign Wnaiw6 = (!Toi7z6[3]);
assign Avi7v6 = (U20jy6 ? K72jy6 : I52nv6);
assign U20jy6 = (~(Doaiw6 & Zh18x6));
assign Doaiw6 = (~(S72jy6 | Toi7z6[2]));
assign Tui7v6 = (I82jy6 ? A82jy6 : STCLK);
assign Mui7v6 = (I82jy6 ? Q82jy6 : A82jy6);
assign A82jy6 = (!Qg67z6);
assign Fui7v6 = (I82jy6 ? Cndet6 : Q82jy6);
assign I82jy6 = (~(Axaiw6 & A8cet6));
assign Axaiw6 = (~(K72jy6 | STCALIB[25]));
assign K72jy6 = (!Me77z6);
assign Q82jy6 = (!As67z6);
assign Yti7v6 = (Muziy6 ? I52nv6 : H1j7z6[2]);
assign Muziy6 = (Y82jy6 & Zh18x6);
assign Zh18x6 = (~(P48iw6 | Twaiw6));
assign Twaiw6 = (!Bqi7z6[0]);
assign P48iw6 = (!R58iw6);
assign Rti7v6 = (Hr4yx6 ? I52nv6 : X66ft6);
assign Kti7v6 = (Eu1jy6 ? I52nv6 : Scs7z6[2]);
assign Eu1jy6 = (Zmryx6 & Mq1jy6);
assign Zmryx6 = (G92jy6 & Mm27v6);
assign G92jy6 = (~(O92jy6 | Zfs7z6[7]));
assign Dti7v6 = (W92jy6 ? Cx4iw6 : Ies7z6[23]);
assign Wsi7v6 = (W92jy6 ? D85iw6 : Ies7z6[22]);
assign Psi7v6 = (W92jy6 ? Ej5iw6 : Ies7z6[21]);
assign Isi7v6 = (W92jy6 ? Bl5iw6 : Ies7z6[20]);
assign Bsi7v6 = (W92jy6 ? Mn5iw6 : Ies7z6[19]);
assign Uri7v6 = (W92jy6 ? Jp5iw6 : Ies7z6[18]);
assign Nri7v6 = (W92jy6 ? Gr5iw6 : Ies7z6[17]);
assign Gri7v6 = (Aw1jy6 ? I52nv6 : Ies7z6[2]);
assign Aw1jy6 = (Ea2jy6 & Cv1jy6);
assign Ea2jy6 = (Ihs7z6[0] & Ma2jy6);
assign Ma2jy6 = (~(C397z6 & Scs7z6[0]));
assign Zqi7v6 = (Y81jy6 ? I52nv6 : Ee77z6);
assign Y81jy6 = (Xid8x6 & Vcpyx6);
assign Vcpyx6 = (Ua2jy6 & Cb2jy6);
assign Cb2jy6 = (Kb2jy6 & Sb2jy6);
assign Kb2jy6 = (~(Xfymz6[11] | Xfymz6[8]));
assign Ua2jy6 = (A81jy6 & Xfymz6[9]);
assign A81jy6 = (Ac2jy6 & B6pyx6);
assign B6pyx6 = (Aslhy6 & Ic2jy6);
assign Ac2jy6 = (D9pyx6 & R6pyx6);
assign Sqi7v6 = (C71jy6 ? I52nv6 : Kmymz6[2]);
assign Lqi7v6 = (G91jy6 ? I52nv6 : Biymz6[2]);
assign Eqi7v6 = (Hn5yx6 ? Aw77z6 : Rzr7z6[1]);
assign Xpi7v6 = (Hn5yx6 ? Sv77z6 : Rzr7z6[2]);
assign Qpi7v6 = (Hn5yx6 ? Kv77z6 : Rzr7z6[3]);
assign Jpi7v6 = (Hn5yx6 ? Cv77z6 : Rzr7z6[4]);
assign Cpi7v6 = (Hn5yx6 ? Uu77z6 : Rzr7z6[5]);
assign Voi7v6 = (Hn5yx6 ? Mu77z6 : Rzr7z6[6]);
assign Ooi7v6 = (Hn5yx6 ? Eu77z6 : Rzr7z6[7]);
assign Hoi7v6 = (Hn5yx6 ? Wt77z6 : Rzr7z6[8]);
assign Aoi7v6 = (Hn5yx6 ? Ot77z6 : Rzr7z6[9]);
assign Tni7v6 = (Hn5yx6 ? Gt77z6 : Rzr7z6[10]);
assign Mni7v6 = (Hn5yx6 ? Ys77z6 : Rzr7z6[11]);
assign Fni7v6 = (Hn5yx6 ? Qs77z6 : Rzr7z6[12]);
assign Ymi7v6 = (Hn5yx6 ? Is77z6 : Rzr7z6[13]);
assign Rmi7v6 = (Hn5yx6 ? As77z6 : Rzr7z6[14]);
assign Kmi7v6 = (Hn5yx6 ? Sr77z6 : Rzr7z6[15]);
assign Dmi7v6 = (Hn5yx6 ? Kr77z6 : Rzr7z6[16]);
assign Wli7v6 = (Hn5yx6 ? Cr77z6 : Rzr7z6[17]);
assign Pli7v6 = (Hn5yx6 ? Uq77z6 : Rzr7z6[18]);
assign Ili7v6 = (Hn5yx6 ? Mq77z6 : Rzr7z6[19]);
assign Bli7v6 = (Hn5yx6 ? Eq77z6 : Rzr7z6[20]);
assign Uki7v6 = (Hn5yx6 ? Wp77z6 : Rzr7z6[21]);
assign Nki7v6 = (Hn5yx6 ? Op77z6 : Rzr7z6[22]);
assign Gki7v6 = (Hn5yx6 ? Gp77z6 : Rzr7z6[23]);
assign Zji7v6 = (Hn5yx6 ? Yo77z6 : Rzr7z6[24]);
assign Sji7v6 = (Hn5yx6 ? Qo77z6 : Rzr7z6[25]);
assign Lji7v6 = (Hn5yx6 ? Io77z6 : Rzr7z6[26]);
assign Eji7v6 = (Hn5yx6 ? Ao77z6 : Rzr7z6[27]);
assign Xii7v6 = (Hn5yx6 ? Sn77z6 : Rzr7z6[28]);
assign Qii7v6 = (Hn5yx6 ? Kn77z6 : Rzr7z6[29]);
assign Jii7v6 = (Hn5yx6 ? Cn77z6 : Rzr7z6[30]);
assign Cii7v6 = (Hn5yx6 ? Um77z6 : Rzr7z6[31]);
assign Hn5yx6 = (~(Kygnv6 | Wfo7v6));
assign Vhi7v6 = (P9get6 ? E6a7z6 : Jqj7z6[3]);
assign E6a7z6 = (~(Qc2jy6 & Yc2jy6));
assign Yc2jy6 = (~(Gd2jy6 & Ykliy6));
assign Ykliy6 = (~(Od2jy6 & Wd2jy6));
assign Wd2jy6 = (~(Ee2jy6 & Me2jy6));
assign Me2jy6 = (~(Ue2jy6 | Cvniy6));
assign Ue2jy6 = (Lh18x6 | Q0oiy6);
assign Ee2jy6 = (Cf2jy6 & W9ziy6);
assign Cf2jy6 = (!Gd2jy6);
assign Od2jy6 = (~(Kf2jy6 & Sf2jy6));
assign Sf2jy6 = (Ag2jy6 & Ig2jy6);
assign Ig2jy6 = (~(Qg2jy6 & Eqwiy6));
assign Eqwiy6 = (Yg2jy6 & Ccr7x6);
assign Ccr7x6 = (~(Gh2jy6 & Jm98x6));
assign Yg2jy6 = (Ui2nv6 & Xg2nv6);
assign Xg2nv6 = (!X7get6);
assign Ui2nv6 = (Xsinv6 | Rdmov6);
assign Rdmov6 = (~(Oh2jy6 & Za2nv6));
assign Oh2jy6 = (~(Xxjov6 & Wh2jy6));
assign Wh2jy6 = (~(Ei2jy6 & Mi2jy6));
assign Mi2jy6 = (~(Ui2jy6 & Cj2jy6));
assign Cj2jy6 = (Kj2jy6 & Pqliw6);
assign Kj2jy6 = (~(Sj2jy6 & Ak2jy6));
assign Ak2jy6 = (Xnliw6 ? Qk2jy6 : Ik2jy6);
assign Qk2jy6 = (~(Nob7z6[4] & Yk2jy6));
assign Yk2jy6 = (~(Gl2jy6 & Ol2jy6));
assign Ol2jy6 = (Wl2jy6 & Em2jy6);
assign Em2jy6 = (Mm2jy6 & Um2jy6);
assign Um2jy6 = (~(Cn2jy6 & G5j7z6[3]));
assign Mm2jy6 = (Kn2jy6 & Sn2jy6);
assign Sn2jy6 = (~(Ao2jy6 & G5j7z6[0]));
assign Kn2jy6 = (~(Jfmiw6 & G5j7z6[2]));
assign Wl2jy6 = (Io2jy6 & Qo2jy6);
assign Qo2jy6 = (~(Cshov6 & G5j7z6[4]));
assign Io2jy6 = (~(I2oiw6 & G5j7z6[5]));
assign Gl2jy6 = (Yo2jy6 & Gp2jy6);
assign Gp2jy6 = (Op2jy6 & Wp2jy6);
assign Wp2jy6 = (~(G5j7z6[12] & L1i7x6));
assign Op2jy6 = (Eq2jy6 & Mq2jy6);
assign Mq2jy6 = (~(G5j7z6[6] & Rphov6));
assign Eq2jy6 = (~(G5j7z6[11] & Hzh7x6));
assign Yo2jy6 = (Uq2jy6 & Cr2jy6);
assign Cr2jy6 = (~(G5j7z6[14] & P3i7x6));
assign Uq2jy6 = (~(G5j7z6[15] & V6i7x6));
assign Ik2jy6 = (Nob7z6[4] ? Sr2jy6 : Kr2jy6);
assign Sr2jy6 = (As2jy6 & Is2jy6);
assign Is2jy6 = (Qs2jy6 & Ys2jy6);
assign Ys2jy6 = (Gt2jy6 & Ot2jy6);
assign Ot2jy6 = (Wt2jy6 & Eu2jy6);
assign Eu2jy6 = (~(G5j7z6[32] & Ao2jy6));
assign Wt2jy6 = (~(G5j7z6[33] & Nuniw6));
assign Gt2jy6 = (Mu2jy6 & Uu2jy6);
assign Uu2jy6 = (~(G5j7z6[34] & Jfmiw6));
assign Mu2jy6 = (~(G5j7z6[35] & Cn2jy6));
assign Qs2jy6 = (Cv2jy6 & Kv2jy6);
assign Kv2jy6 = (Sv2jy6 & Aw2jy6);
assign Aw2jy6 = (~(Cshov6 & G5j7z6[36]));
assign Sv2jy6 = (~(I2oiw6 & G5j7z6[37]));
assign Cv2jy6 = (Iw2jy6 & Qw2jy6);
assign Qw2jy6 = (~(G5j7z6[38] & Rphov6));
assign Iw2jy6 = (~(J6oiw6 & G5j7z6[39]));
assign As2jy6 = (Yw2jy6 & Gx2jy6);
assign Gx2jy6 = (Ox2jy6 & Wx2jy6);
assign Wx2jy6 = (Ey2jy6 & My2jy6);
assign My2jy6 = (~(Uy2jy6 & G5j7z6[40]));
assign Ey2jy6 = (~(Mbj7x6 & G5j7z6[41]));
assign Ox2jy6 = (Cz2jy6 & Kz2jy6);
assign Kz2jy6 = (~(Nfj7x6 & G5j7z6[42]));
assign Cz2jy6 = (~(G5j7z6[43] & Hzh7x6));
assign Yw2jy6 = (Sz2jy6 & A03jy6);
assign A03jy6 = (I03jy6 & Q03jy6);
assign Q03jy6 = (~(G5j7z6[44] & L1i7x6));
assign I03jy6 = (~(Jrj7x6 & G5j7z6[45]));
assign Sz2jy6 = (Y03jy6 & G13jy6);
assign G13jy6 = (~(G5j7z6[46] & P3i7x6));
assign Y03jy6 = (~(G5j7z6[47] & V6i7x6));
assign Kr2jy6 = (O13jy6 & W13jy6);
assign W13jy6 = (E23jy6 & M23jy6);
assign M23jy6 = (U23jy6 & C33jy6);
assign C33jy6 = (~(G5j7z6[19] & Cn2jy6));
assign U23jy6 = (K33jy6 & S33jy6);
assign S33jy6 = (~(Ao2jy6 & G5j7z6[16]));
assign K33jy6 = (~(G5j7z6[18] & Jfmiw6));
assign E23jy6 = (A43jy6 & I43jy6);
assign I43jy6 = (~(Cshov6 & G5j7z6[20]));
assign A43jy6 = (~(I2oiw6 & G5j7z6[21]));
assign O13jy6 = (Q43jy6 & Y43jy6);
assign Y43jy6 = (G53jy6 & O53jy6);
assign O53jy6 = (~(G5j7z6[28] & L1i7x6));
assign G53jy6 = (W53jy6 & E63jy6);
assign E63jy6 = (~(G5j7z6[22] & Rphov6));
assign W53jy6 = (~(G5j7z6[27] & Hzh7x6));
assign Q43jy6 = (M63jy6 & U63jy6);
assign U63jy6 = (~(G5j7z6[30] & P3i7x6));
assign M63jy6 = (~(G5j7z6[31] & V6i7x6));
assign Sj2jy6 = (C73jy6 & K73jy6);
assign K73jy6 = (~(S73jy6 & A83jy6));
assign A83jy6 = (~(I83jy6 & Q83jy6));
assign Q83jy6 = (Y83jy6 & G93jy6);
assign G93jy6 = (O93jy6 & W93jy6);
assign W93jy6 = (~(Ea3jy6 & Omliw6));
assign Ea3jy6 = (~(Ma3jy6 & Ua3jy6));
assign Ua3jy6 = (Cb3jy6 & Kb3jy6);
assign Kb3jy6 = (~(Nob7z6[0] & Sb3jy6));
assign Sb3jy6 = (~(Ac3jy6 & Ic3jy6));
assign Ic3jy6 = (~(Qc3jy6 & X3get6));
assign Ac3jy6 = (~(Z3j7z6[11] & Yc3jy6));
assign Cb3jy6 = (~(Nob7z6[1] & Gd3jy6));
assign Gd3jy6 = (~(Od3jy6 & Wd3jy6));
assign Wd3jy6 = (~(Z3j7z6[3] & Ee3jy6));
assign Od3jy6 = (~(Fjadt6 & Me3jy6));
assign Ma3jy6 = (Ue3jy6 & Cf3jy6);
assign Cf3jy6 = (~(Z3j7z6[1] & Kf3jy6));
assign Ue3jy6 = (~(Nob7z6[3] & Sf3jy6));
assign Sf3jy6 = (~(Ag3jy6 & Ig3jy6));
assign Ig3jy6 = (~(Z3j7z6[7] & Wjliw6));
assign Ag3jy6 = (Qg3jy6 & Yg3jy6);
assign Yg3jy6 = (~(Z3j7z6[10] & Gh3jy6));
assign Qg3jy6 = (~(Z3j7z6[8] & Giliw6));
assign O93jy6 = (~(Nuniw6 & G5j7z6[1]));
assign Y83jy6 = (Oh3jy6 & Wh3jy6);
assign Wh3jy6 = (~(J6oiw6 & G5j7z6[7]));
assign Oh3jy6 = (~(G5j7z6[8] & Uy2jy6));
assign I83jy6 = (Ei3jy6 & Mi3jy6);
assign Mi3jy6 = (~(Jrj7x6 & G5j7z6[13]));
assign Ei3jy6 = (Ui3jy6 & Cj3jy6);
assign Cj3jy6 = (~(G5j7z6[9] & Mbj7x6));
assign Ui3jy6 = (~(G5j7z6[10] & Nfj7x6));
assign C73jy6 = (Nob7z6[6] ? Sj3jy6 : Kj3jy6);
assign Sj3jy6 = (Ak3jy6 & Ik3jy6);
assign Ik3jy6 = (Qk3jy6 & Yk3jy6);
assign Yk3jy6 = (Gl3jy6 & Ol3jy6);
assign Ol3jy6 = (Wl3jy6 & Em3jy6);
assign Em3jy6 = (~(G5j7z6[48] & Ao2jy6));
assign Wl3jy6 = (~(G5j7z6[49] & Nuniw6));
assign Gl3jy6 = (Mm3jy6 & Um3jy6);
assign Um3jy6 = (~(G5j7z6[50] & Jfmiw6));
assign Mm3jy6 = (~(G5j7z6[51] & Cn2jy6));
assign Qk3jy6 = (Cn3jy6 & Kn3jy6);
assign Kn3jy6 = (Sn3jy6 & Ao3jy6);
assign Ao3jy6 = (~(Cshov6 & G5j7z6[52]));
assign Sn3jy6 = (~(I2oiw6 & G5j7z6[53]));
assign Cn3jy6 = (Io3jy6 & Qo3jy6);
assign Qo3jy6 = (~(G5j7z6[54] & Rphov6));
assign Io3jy6 = (~(J6oiw6 & G5j7z6[55]));
assign Ak3jy6 = (Yo3jy6 & Gp3jy6);
assign Gp3jy6 = (Op3jy6 & Wp3jy6);
assign Wp3jy6 = (Eq3jy6 & Mq3jy6);
assign Mq3jy6 = (~(G5j7z6[56] & Uy2jy6));
assign Eq3jy6 = (~(G5j7z6[57] & Mbj7x6));
assign Op3jy6 = (Uq3jy6 & Cr3jy6);
assign Cr3jy6 = (~(G5j7z6[58] & Nfj7x6));
assign Uq3jy6 = (~(G5j7z6[59] & Hzh7x6));
assign Yo3jy6 = (Kr3jy6 & Sr3jy6);
assign Sr3jy6 = (As3jy6 & Is3jy6);
assign Is3jy6 = (~(G5j7z6[60] & L1i7x6));
assign As3jy6 = (~(Jrj7x6 & G5j7z6[61]));
assign Kr3jy6 = (Qs3jy6 & Ys3jy6);
assign Ys3jy6 = (~(G5j7z6[62] & P3i7x6));
assign Qs3jy6 = (~(G5j7z6[63] & V6i7x6));
assign Kj3jy6 = (~(Gt3jy6 & Omliw6));
assign Gt3jy6 = (~(Ot3jy6 & Wt3jy6));
assign Wt3jy6 = (Eu3jy6 & Mu3jy6);
assign Mu3jy6 = (~(Uy2jy6 & G5j7z6[24]));
assign Eu3jy6 = (Uu3jy6 & Cv3jy6);
assign Cv3jy6 = (~(G5j7z6[17] & Nuniw6));
assign Uu3jy6 = (~(J6oiw6 & G5j7z6[23]));
assign Ot3jy6 = (Kv3jy6 & Sv3jy6);
assign Sv3jy6 = (~(Jrj7x6 & G5j7z6[29]));
assign Kv3jy6 = (Aw3jy6 & Iw3jy6);
assign Iw3jy6 = (~(Mbj7x6 & G5j7z6[25]));
assign Aw3jy6 = (~(Nfj7x6 & G5j7z6[26]));
assign Ui2jy6 = (Qw3jy6 & Yw3jy6);
assign Yw3jy6 = (~(Nob7z6[6] & Gx3jy6));
assign Gx3jy6 = (~(Xnliw6 & Omliw6));
assign Qw3jy6 = (~(Ox3jy6 & Wx3jy6));
assign Wx3jy6 = (~(Ey3jy6 & My3jy6));
assign My3jy6 = (~(Kf3jy6 & Uy3jy6));
assign Uy3jy6 = (!Ee3jy6);
assign Ey3jy6 = (~(J6oiw6 | Cz3jy6));
assign Ei2jy6 = (~(Kz3jy6 & Cshov6));
assign Kz3jy6 = (Z3j7z6[0] & Sz3jy6);
assign Qg2jy6 = (A04jy6 & I04jy6);
assign I04jy6 = (~(Q04jy6 & Y04jy6));
assign Y04jy6 = (~(G14jy6 & Ldr7x6));
assign A04jy6 = (Ldr7x6 | G14jy6);
assign G14jy6 = (O14jy6 & W14jy6);
assign W14jy6 = (~(E24jy6 & Ger7x6));
assign O14jy6 = (~(M24jy6 & U24jy6));
assign M24jy6 = (C34jy6 & CURRPRI[5]);
assign C34jy6 = (~(K34jy6 & Bfr7x6));
assign Bfr7x6 = (!Ger7x6);
assign Ger7x6 = (Zyl8v6 & CURRPRI[6]);
assign Ldr7x6 = (~(H1m8v6 & CURRPRI[7]));
assign Ag2jy6 = (S34jy6 & Hs98x6);
assign Hs98x6 = (!Nmadt6);
assign Kf2jy6 = (A44jy6 & I44jy6);
assign I44jy6 = (~(Q44jy6 & Snwiy6));
assign Snwiy6 = (~(Y44jy6 & G54jy6));
assign G54jy6 = (O54jy6 & W54jy6);
assign O54jy6 = (~(E64jy6 | M64jy6));
assign Y44jy6 = (U64jy6 & C74jy6);
assign U64jy6 = (~(K74jy6 | S74jy6));
assign Q44jy6 = (~(A84jy6 & I84jy6));
assign I84jy6 = (~(Q84jy6 & Y84jy6));
assign Q84jy6 = (G94jy6 | O94jy6);
assign A84jy6 = (~(O94jy6 & G94jy6));
assign G94jy6 = (!Y0t7x6);
assign Y0t7x6 = (W94jy6 & H1m8v6);
assign W94jy6 = (Ua4jy6 ? Ma4jy6 : Ea4jy6);
assign Ea4jy6 = (!Cb4jy6);
assign O94jy6 = (Kb4jy6 & Sb4jy6);
assign Sb4jy6 = (~(E24jy6 & I6t7x6));
assign I6t7x6 = (!B6t7x6);
assign Kb4jy6 = (~(Ac4jy6 & U24jy6));
assign Ac4jy6 = (N5t7x6 & Ic4jy6);
assign Ic4jy6 = (~(K34jy6 & B6t7x6));
assign B6t7x6 = (Qc4jy6 | Yc4jy6);
assign Yc4jy6 = (!Zyl8v6);
assign Qc4jy6 = (Ua4jy6 ? Od4jy6 : Gd4jy6);
assign Ua4jy6 = (!Wd4jy6);
assign N5t7x6 = (!Ee4jy6);
assign Ee4jy6 = (Wd4jy6 ? Ue4jy6 : Me4jy6);
assign Wd4jy6 = (Cf4jy6 & E64jy6);
assign E64jy6 = (Kf4jy6 | Sf4jy6);
assign Kf4jy6 = (Ag4jy6 | Ig4jy6);
assign Cf4jy6 = (~(Qg4jy6 & Yg4jy6));
assign Yg4jy6 = (~(Cb4jy6 & Gh4jy6));
assign Gh4jy6 = (~(Oh4jy6 & Wh4jy6));
assign Oh4jy6 = (Ei4jy6 & Mi4jy6);
assign Mi4jy6 = (Me4jy6 | Ui4jy6);
assign Ui4jy6 = (Cj4jy6 & Od4jy6);
assign Ei4jy6 = (~(Kj4jy6 & Sj4jy6));
assign Cb4jy6 = (Qk4jy6 ? Ik4jy6 : Ak4jy6);
assign Qg4jy6 = (Yk4jy6 & Gl4jy6);
assign Gl4jy6 = (~(Ol4jy6 & Ma4jy6));
assign Ma4jy6 = (Kj4jy6 & Sj4jy6);
assign Sj4jy6 = (Wl4jy6 | Em4jy6);
assign Kj4jy6 = (~(Mm4jy6 & Wl4jy6));
assign Ol4jy6 = (Um4jy6 & Cn4jy6);
assign Cn4jy6 = (~(Me4jy6 & Wh4jy6));
assign Wh4jy6 = (~(Kn4jy6 & Gd4jy6));
assign Kn4jy6 = (!Od4jy6);
assign Um4jy6 = (~(Cj4jy6 & Od4jy6));
assign Od4jy6 = (Io4jy6 ? Ao4jy6 : Sn4jy6);
assign Cj4jy6 = (!Gd4jy6);
assign Gd4jy6 = (Qk4jy6 ? Yo4jy6 : Qo4jy6);
assign Yk4jy6 = (~(Gp4jy6 & Op4jy6));
assign Gp4jy6 = (Wl4jy6 & Wp4jy6);
assign Wl4jy6 = (!Io4jy6);
assign Ue4jy6 = (Qk4jy6 ? Mq4jy6 : Eq4jy6);
assign Qk4jy6 = (~(Uq4jy6 & Cr4jy6));
assign Cr4jy6 = (~(Kr4jy6 & Ig4jy6));
assign Ig4jy6 = (~(Sr4jy6 & As4jy6));
assign As4jy6 = (Is4jy6 & Mpoiw6);
assign Is4jy6 = (~(Baniw6 | Ntoiw6));
assign Sr4jy6 = (Qs4jy6 & Ys4jy6);
assign Qs4jy6 = (Gt4jy6 & Ot4jy6);
assign Kr4jy6 = (~(Wt4jy6 & Eu4jy6));
assign Eu4jy6 = (~(Ik4jy6 & Mu4jy6));
assign Mu4jy6 = (~(Ak4jy6 & Uu4jy6));
assign Ik4jy6 = (Sv4jy6 ? Kv4jy6 : Cv4jy6);
assign Wt4jy6 = (Uu4jy6 | Ak4jy6);
assign Ak4jy6 = (Qw4jy6 ? Iw4jy6 : Aw4jy6);
assign Uu4jy6 = (~(Yw4jy6 & Gx4jy6));
assign Gx4jy6 = (~(Eq4jy6 & Ox4jy6));
assign Ox4jy6 = (~(Yo4jy6 & Wx4jy6));
assign Yw4jy6 = (Wx4jy6 | Yo4jy6);
assign Yo4jy6 = (Sv4jy6 ? My4jy6 : Ey4jy6);
assign Wx4jy6 = (!Qo4jy6);
assign Qo4jy6 = (Qw4jy6 ? Cz4jy6 : Uy4jy6);
assign Uq4jy6 = (Sf4jy6 | Ag4jy6);
assign Sf4jy6 = (~(Kz4jy6 & Sz4jy6));
assign Kz4jy6 = (~(A05jy6 | I05jy6));
assign Mq4jy6 = (Sv4jy6 ? Y05jy6 : Q05jy6);
assign Sv4jy6 = (G15jy6 & O15jy6);
assign O15jy6 = (~(W15jy6 & E25jy6));
assign E25jy6 = (~(Kv4jy6 & M25jy6));
assign W15jy6 = (U25jy6 & C35jy6);
assign C35jy6 = (~(K35jy6 & S35jy6));
assign S35jy6 = (M25jy6 | Kv4jy6);
assign Kv4jy6 = (Q45jy6 ? I45jy6 : A45jy6);
assign M25jy6 = (!Cv4jy6);
assign Cv4jy6 = (O55jy6 ? G55jy6 : Y45jy6);
assign K35jy6 = (W55jy6 & E65jy6);
assign E65jy6 = (My4jy6 | M65jy6);
assign M65jy6 = (~(Q05jy6 | Ey4jy6));
assign My4jy6 = (Q45jy6 ? C75jy6 : U65jy6);
assign C75jy6 = (!K75jy6);
assign W55jy6 = (~(Ey4jy6 & Q05jy6));
assign Ey4jy6 = (O55jy6 ? A85jy6 : S75jy6);
assign A85jy6 = (!I85jy6);
assign U25jy6 = (~(Q85jy6 & O55jy6));
assign Q85jy6 = (Ot4jy6 & Mpoiw6);
assign G15jy6 = (~(Ys4jy6 & Gt4jy6));
assign Gt4jy6 = (!Y85jy6);
assign Y05jy6 = (Q45jy6 ? O95jy6 : G95jy6);
assign Q45jy6 = (W95jy6 | Ys4jy6);
assign Ys4jy6 = (Ea5jy6 & Ma5jy6);
assign Ma5jy6 = (~(G5j7z6[55] & Ua5jy6));
assign Ea5jy6 = (Cb5jy6 & Kb5jy6);
assign Kb5jy6 = (Px2nv6 | Sb5jy6);
assign Px2nv6 = (Fnl7x6 & Sjl7x6);
assign Sjl7x6 = (!G5j7z6[54]);
assign Fnl7x6 = (!G5j7z6[55]);
assign Cb5jy6 = (~(G5j7z6[54] & Ac5jy6));
assign W95jy6 = (Ic5jy6 & Qc5jy6);
assign Qc5jy6 = (Yc5jy6 & Y85jy6);
assign Y85jy6 = (~(Gd5jy6 & Od5jy6));
assign Od5jy6 = (~(G5j7z6[53] & Wd5jy6));
assign Gd5jy6 = (Ee5jy6 & Me5jy6);
assign Me5jy6 = (~(Wx2nv6 & Ytl7x6));
assign Wx2nv6 = (~(Fgl7x6 & Scl7x6));
assign Scl7x6 = (!G5j7z6[52]);
assign Fgl7x6 = (!G5j7z6[53]);
assign Ee5jy6 = (~(G5j7z6[52] & Ue5jy6));
assign Yc5jy6 = (~(Cf5jy6 & G95jy6));
assign Cf5jy6 = (Kf5jy6 & Sf5jy6);
assign Sf5jy6 = (U65jy6 | K75jy6);
assign Ic5jy6 = (Ag5jy6 & Ig5jy6);
assign Ig5jy6 = (~(Qg5jy6 & K75jy6));
assign K75jy6 = (Yg5jy6 ? Lgj7z6[160] : Lgj7z6[157]);
assign Qg5jy6 = (U65jy6 & Kf5jy6);
assign Kf5jy6 = (A45jy6 | Gh5jy6);
assign U65jy6 = (Oh5jy6 ? C2u7x6 : J2u7x6);
assign Ag5jy6 = (~(Gh5jy6 & A45jy6));
assign A45jy6 = (Oh5jy6 ? Wh5jy6 : Am88x6);
assign Wh5jy6 = (!Lgj7z6[164]);
assign Gh5jy6 = (!I45jy6);
assign I45jy6 = (Yg5jy6 ? V1u7x6 : O1u7x6);
assign O95jy6 = (Yg5jy6 ? M0u7x6 : F0u7x6);
assign Yg5jy6 = (Ei5jy6 & G5j7z6[53]);
assign Ei5jy6 = (Mi5jy6 & Ui5jy6);
assign Ui5jy6 = (Cj5jy6 | U4u7x6);
assign U4u7x6 = (~(Kj5jy6 & Sj5jy6));
assign Sj5jy6 = (~(Lgj7z6[158] & V1u7x6));
assign V1u7x6 = (!Lgj7z6[161]);
assign Kj5jy6 = (Ak5jy6 & Ik5jy6);
assign Ik5jy6 = (~(Qk5jy6 & Yk5jy6));
assign Yk5jy6 = (Gl5jy6 & M0u7x6);
assign Gl5jy6 = (~(Lgj7z6[160] & H888x6));
assign H888x6 = (!Lgj7z6[157]);
assign Qk5jy6 = (Lgj7z6[156] & Ol5jy6);
assign Ol5jy6 = (~(Lgj7z6[161] & O1u7x6));
assign Ak5jy6 = (~(Wl5jy6 & Lgj7z6[157]));
assign Wl5jy6 = (~(Em5jy6 | Lgj7z6[160]));
assign Em5jy6 = (Lgj7z6[161] & O1u7x6);
assign O1u7x6 = (!Lgj7z6[158]);
assign Cj5jy6 = (~(G5j7z6[52] & Mm5jy6));
assign Mm5jy6 = (~(Cshov6 & Sb5jy6));
assign Mi5jy6 = (~(I2oiw6 & Sb5jy6));
assign M0u7x6 = (!Lgj7z6[159]);
assign F0u7x6 = (!Lgj7z6[156]);
assign G95jy6 = (Oh5jy6 ? Cg88x6 : Rk88x6);
assign Oh5jy6 = (~(Um5jy6 & G5j7z6[55]));
assign Um5jy6 = (Cn5jy6 & Kn5jy6);
assign Kn5jy6 = (~(Sn5jy6 & L3u7x6));
assign L3u7x6 = (Ao5jy6 & Io5jy6);
assign Io5jy6 = (~(Lgj7z6[164] & Am88x6));
assign Ao5jy6 = (Qo5jy6 & Yo5jy6);
assign Yo5jy6 = (~(Gp5jy6 & Op5jy6));
assign Op5jy6 = (Wp5jy6 & Rk88x6);
assign Gp5jy6 = (Lgj7z6[162] & Eq5jy6);
assign Eq5jy6 = (~(Lgj7z6[166] & C2u7x6));
assign C2u7x6 = (!Lgj7z6[163]);
assign Qo5jy6 = (~(Mq5jy6 & Lgj7z6[163]));
assign Mq5jy6 = (Wp5jy6 & J2u7x6);
assign J2u7x6 = (!Lgj7z6[166]);
assign Wp5jy6 = (Am88x6 | Lgj7z6[164]);
assign Am88x6 = (!Lgj7z6[167]);
assign Sn5jy6 = (G5j7z6[54] & Uq5jy6);
assign Uq5jy6 = (~(Sb5jy6 & Rphov6));
assign Cn5jy6 = (~(J6oiw6 & Sb5jy6));
assign Cg88x6 = (!Lgj7z6[162]);
assign Rk88x6 = (!Lgj7z6[165]);
assign Q05jy6 = (O55jy6 ? Kr5jy6 : Cr5jy6);
assign O55jy6 = (~(Sr5jy6 & As5jy6));
assign As5jy6 = (Baniw6 | Ntoiw6);
assign Sr5jy6 = (~(Is5jy6 & Qs5jy6));
assign Qs5jy6 = (Ys5jy6 & Gt5jy6);
assign Gt5jy6 = (~(Ot5jy6 & Cr5jy6));
assign Ot5jy6 = (Wt5jy6 & Eu5jy6);
assign Wt5jy6 = (S75jy6 | I85jy6);
assign Ys5jy6 = (~(Mu5jy6 & I85jy6));
assign I85jy6 = (Uu5jy6 ? Lgj7z6[148] : Lgj7z6[145]);
assign Mu5jy6 = (S75jy6 & Eu5jy6);
assign Eu5jy6 = (Y45jy6 | Cv5jy6);
assign S75jy6 = (Kv5jy6 ? Gbu7x6 : Zau7x6);
assign Kv5jy6 = (!Sv5jy6);
assign Is5jy6 = (Aw5jy6 & Iw5jy6);
assign Iw5jy6 = (~(Cv5jy6 & Y45jy6));
assign Y45jy6 = (Sv5jy6 ? S388x6 : Qw5jy6);
assign Cv5jy6 = (!G55jy6);
assign G55jy6 = (Uu5jy6 ? Vu78x6 : Yw5jy6);
assign Aw5jy6 = (~(Ot4jy6 & Mpoiw6));
assign Ot4jy6 = (!F5niw6);
assign Kr5jy6 = (Uu5jy6 ? Qvt7x6 : Xvt7x6);
assign Uu5jy6 = (~(Mpoiw6 | Gx5jy6));
assign Gx5jy6 = (Feu7x6 & F5niw6);
assign F5niw6 = (G5j7z6[48] & Ox5jy6);
assign Ox5jy6 = (~(Sb5jy6 & Ao2jy6));
assign Feu7x6 = (Wx5jy6 & Ey5jy6);
assign Ey5jy6 = (~(My5jy6 & Lgj7z6[145]));
assign My5jy6 = (Uy5jy6 & Ddu7x6);
assign Ddu7x6 = (!Lgj7z6[148]);
assign Wx5jy6 = (Cz5jy6 & Kz5jy6);
assign Kz5jy6 = (~(Sz5jy6 & A06jy6));
assign A06jy6 = (I06jy6 & Qvt7x6);
assign I06jy6 = (~(Lgj7z6[148] & Wcu7x6));
assign Wcu7x6 = (!Lgj7z6[145]);
assign Sz5jy6 = (Lgj7z6[144] & Uy5jy6);
assign Uy5jy6 = (~(Lgj7z6[149] & Yw5jy6));
assign Yw5jy6 = (!Lgj7z6[146]);
assign Cz5jy6 = (~(Lgj7z6[146] & Vu78x6));
assign Vu78x6 = (!Lgj7z6[149]);
assign Mpoiw6 = (~(G5j7z6[49] & Q06jy6));
assign Q06jy6 = (~(Sb5jy6 & Nuniw6));
assign Qvt7x6 = (!Lgj7z6[147]);
assign Xvt7x6 = (!Lgj7z6[144]);
assign Cr5jy6 = (Sv5jy6 ? C9u7x6 : J9u7x6);
assign Sv5jy6 = (Ntoiw6 & Y06jy6);
assign Y06jy6 = (~(Baniw6 & Icu7x6));
assign Icu7x6 = (G16jy6 & O16jy6);
assign O16jy6 = (~(Lgj7z6[152] & S388x6));
assign S388x6 = (!Lgj7z6[155]);
assign G16jy6 = (W16jy6 & E26jy6);
assign E26jy6 = (~(M26jy6 & U26jy6));
assign U26jy6 = (C36jy6 & C9u7x6);
assign C36jy6 = (~(Lgj7z6[154] & Gbu7x6));
assign Gbu7x6 = (!Lgj7z6[151]);
assign M26jy6 = (Lgj7z6[150] & K36jy6);
assign W16jy6 = (~(S36jy6 & Lgj7z6[151]));
assign S36jy6 = (K36jy6 & Zau7x6);
assign Zau7x6 = (!Lgj7z6[154]);
assign K36jy6 = (~(Lgj7z6[155] & Qw5jy6));
assign Qw5jy6 = (!Lgj7z6[152]);
assign Baniw6 = (G5j7z6[50] & A46jy6);
assign A46jy6 = (~(Sb5jy6 & Jfmiw6));
assign Ntoiw6 = (G5j7z6[51] & I46jy6);
assign I46jy6 = (~(Sb5jy6 & Cn2jy6));
assign C9u7x6 = (!Lgj7z6[153]);
assign J9u7x6 = (!Lgj7z6[150]);
assign Eq4jy6 = (Qw4jy6 ? Y46jy6 : Q46jy6);
assign Qw4jy6 = (G56jy6 & O56jy6);
assign O56jy6 = (~(W56jy6 & E66jy6));
assign E66jy6 = (~(Sz4jy6 & M66jy6));
assign Sz4jy6 = (U66jy6 & C76jy6);
assign W56jy6 = (K76jy6 & S76jy6);
assign S76jy6 = (~(Iw4jy6 & A86jy6));
assign A86jy6 = (~(Aw4jy6 & I86jy6));
assign Iw4jy6 = (G96jy6 ? Y86jy6 : Q86jy6);
assign Y86jy6 = (!O96jy6);
assign K76jy6 = (I86jy6 | Aw4jy6);
assign Aw4jy6 = (M66jy6 ? Ea6jy6 : W96jy6);
assign I86jy6 = (Ma6jy6 | Ua6jy6);
assign Ua6jy6 = (Uy4jy6 & Q46jy6);
assign Ma6jy6 = (~(Cz4jy6 | Cb6jy6));
assign Cb6jy6 = (~(Q46jy6 | Uy4jy6));
assign Uy4jy6 = (M66jy6 ? Sb6jy6 : Kb6jy6);
assign Sb6jy6 = (!Ac6jy6);
assign Cz4jy6 = (G96jy6 ? Qc6jy6 : Ic6jy6);
assign Qc6jy6 = (!Yc6jy6);
assign G56jy6 = (A05jy6 | I05jy6);
assign Y46jy6 = (G96jy6 ? Od6jy6 : Gd6jy6);
assign G96jy6 = (~(Wd6jy6 & A05jy6));
assign A05jy6 = (~(Ee6jy6 & Me6jy6));
assign Me6jy6 = (~(G5j7z6[63] & Ue6jy6));
assign Ee6jy6 = (Cf6jy6 & Kf6jy6);
assign Kf6jy6 = (~(Yy2nv6 & Ytl7x6));
assign Yy2nv6 = (~(Y4hov6 & Zbm7x6));
assign Zbm7x6 = (!G5j7z6[62]);
assign Y4hov6 = (!G5j7z6[63]);
assign Cf6jy6 = (~(G5j7z6[62] & Erk7x6));
assign Wd6jy6 = (~(Sf6jy6 & Ag6jy6));
assign Ag6jy6 = (Ig6jy6 & I05jy6);
assign I05jy6 = (~(Qg6jy6 & Yg6jy6));
assign Yg6jy6 = (~(G5j7z6[61] & Ktl7x6));
assign Qg6jy6 = (Gh6jy6 & Oh6jy6);
assign Oh6jy6 = (~(Fz2nv6 & Ytl7x6));
assign Ytl7x6 = (!Sb5jy6);
assign Fz2nv6 = (~(Vvl7x6 & Grl7x6));
assign Grl7x6 = (!G5j7z6[60]);
assign Vvl7x6 = (!G5j7z6[61]);
assign Gh6jy6 = (~(G5j7z6[60] & Qpl7x6));
assign Ig6jy6 = (~(Wh6jy6 & Gd6jy6));
assign Wh6jy6 = (Ei6jy6 & Mi6jy6);
assign Mi6jy6 = (Ic6jy6 | Yc6jy6);
assign Sf6jy6 = (Ui6jy6 & Cj6jy6);
assign Cj6jy6 = (~(Kj6jy6 & Yc6jy6));
assign Yc6jy6 = (Sj6jy6 ? Lgj7z6[181] : Lgj7z6[184]);
assign Sj6jy6 = (!Ak6jy6);
assign Kj6jy6 = (Ic6jy6 & Ei6jy6);
assign Ei6jy6 = (Q86jy6 | O96jy6);
assign Ic6jy6 = (Qk6jy6 ? Ik6jy6 : Zg98x6);
assign Ui6jy6 = (~(O96jy6 & Q86jy6));
assign Q86jy6 = (Qk6jy6 ? En98x6 : Dj98x6);
assign O96jy6 = (Ak6jy6 ? Lgj7z6[185] : Lgj7z6[182]);
assign Od6jy6 = (Ak6jy6 ? Dc98x6 : H798x6);
assign Ak6jy6 = (Yk6jy6 & G5j7z6[61]);
assign Yk6jy6 = (Gl6jy6 & Ol6jy6);
assign Ol6jy6 = (~(Wl6jy6 & Evu7x6));
assign Evu7x6 = (Em6jy6 & Mm6jy6);
assign Mm6jy6 = (~(Lgj7z6[182] & Ae98x6));
assign Em6jy6 = (Um6jy6 & Cn6jy6);
assign Cn6jy6 = (~(Kn6jy6 & Sn6jy6));
assign Sn6jy6 = (~(Ao6jy6 | Lgj7z6[183]));
assign Kn6jy6 = (Lgj7z6[180] & Io6jy6);
assign Io6jy6 = (~(Lgj7z6[184] & Q898x6));
assign Q898x6 = (!Lgj7z6[181]);
assign Um6jy6 = (~(Qo6jy6 & Lgj7z6[181]));
assign Qo6jy6 = (~(Ao6jy6 | Lgj7z6[184]));
assign Ao6jy6 = (~(Ae98x6 | Lgj7z6[182]));
assign Ae98x6 = (!Lgj7z6[185]);
assign Wl6jy6 = (G5j7z6[60] & Yo6jy6);
assign Yo6jy6 = (~(Sb5jy6 & L1i7x6));
assign Gl6jy6 = (~(Jrj7x6 & Sb5jy6));
assign Dc98x6 = (!Lgj7z6[183]);
assign H798x6 = (!Lgj7z6[180]);
assign Gd6jy6 = (Qk6jy6 ? Rru7x6 : Yru7x6);
assign Qk6jy6 = (Gp6jy6 & G5j7z6[63]);
assign Gp6jy6 = (Op6jy6 & Wp6jy6);
assign Wp6jy6 = (~(Eq6jy6 & Vtu7x6));
assign Vtu7x6 = (Mq6jy6 & Uq6jy6);
assign Uq6jy6 = (~(Lgj7z6[188] & En98x6));
assign En98x6 = (!Lgj7z6[191]);
assign Mq6jy6 = (Cr6jy6 & Kr6jy6);
assign Kr6jy6 = (~(Sr6jy6 & As6jy6));
assign As6jy6 = (Is6jy6 & Rru7x6);
assign Is6jy6 = (~(Lgj7z6[190] & Zg98x6));
assign Zg98x6 = (!Lgj7z6[187]);
assign Sr6jy6 = (Lgj7z6[186] & Qs6jy6);
assign Cr6jy6 = (~(Ys6jy6 & Lgj7z6[187]));
assign Ys6jy6 = (Qs6jy6 & Ik6jy6);
assign Ik6jy6 = (!Lgj7z6[190]);
assign Qs6jy6 = (~(Lgj7z6[191] & Dj98x6));
assign Dj98x6 = (!Lgj7z6[188]);
assign Eq6jy6 = (G5j7z6[62] & Gt6jy6);
assign Gt6jy6 = (~(Sb5jy6 & P3i7x6));
assign Op6jy6 = (~(Sb5jy6 & V6i7x6));
assign Rru7x6 = (!Lgj7z6[189]);
assign Yru7x6 = (!Lgj7z6[186]);
assign Q46jy6 = (M66jy6 ? Wt6jy6 : Ot6jy6);
assign M66jy6 = (~(Ag4jy6 & Eu6jy6));
assign Eu6jy6 = (~(Mu6jy6 & Uu6jy6));
assign Uu6jy6 = (Cv6jy6 & Kv6jy6);
assign Kv6jy6 = (~(Sv6jy6 & Ot6jy6));
assign Sv6jy6 = (Aw6jy6 & Iw6jy6);
assign Iw6jy6 = (Kb6jy6 | Ac6jy6);
assign Cv6jy6 = (~(Qw6jy6 & W96jy6));
assign Qw6jy6 = (!Ea6jy6);
assign Mu6jy6 = (Yw6jy6 & Gx6jy6);
assign Gx6jy6 = (~(Ox6jy6 & Ac6jy6));
assign Ac6jy6 = (Wx6jy6 ? Lgj7z6[169] : Lgj7z6[172]);
assign Wx6jy6 = (!Ey6jy6);
assign Ox6jy6 = (Kb6jy6 & Aw6jy6);
assign Aw6jy6 = (~(My6jy6 & Ea6jy6));
assign Ea6jy6 = (Ey6jy6 ? J1v7x6 : C1v7x6);
assign My6jy6 = (!W96jy6);
assign W96jy6 = (Uy6jy6 ? V0v7x6 : O0v7x6);
assign Kb6jy6 = (Uy6jy6 ? Mz88x6 : Cz6jy6);
assign Yw6jy6 = (~(C76jy6 & U66jy6));
assign U66jy6 = (!Gzk7x6);
assign Ag4jy6 = (~(Kz6jy6 & B7l7x6));
assign Kz6jy6 = (~(Sz6jy6 & A07jy6));
assign A07jy6 = (~(I07jy6 & Iq2nv6));
assign Iq2nv6 = (!G5j7z6[58]);
assign Wt6jy6 = (Ey6jy6 ? Vmu7x6 : Cnu7x6);
assign Ey6jy6 = (Gzk7x6 & Q07jy6);
assign Q07jy6 = (C76jy6 | U3v7x6);
assign U3v7x6 = (~(Y07jy6 & G17jy6));
assign G17jy6 = (~(Lgj7z6[170] & J1v7x6));
assign J1v7x6 = (!Lgj7z6[173]);
assign Y07jy6 = (O17jy6 & W17jy6);
assign W17jy6 = (~(E27jy6 & M27jy6));
assign M27jy6 = (~(U27jy6 | Lgj7z6[171]));
assign E27jy6 = (Lgj7z6[168] & C37jy6);
assign C37jy6 = (~(Lgj7z6[172] & Pq88x6));
assign Pq88x6 = (!Lgj7z6[169]);
assign O17jy6 = (~(K37jy6 & Lgj7z6[169]));
assign K37jy6 = (~(U27jy6 | Lgj7z6[172]));
assign U27jy6 = (Lgj7z6[173] & C1v7x6);
assign C1v7x6 = (!Lgj7z6[170]);
assign C76jy6 = (!Fvk7x6);
assign Fvk7x6 = (G5j7z6[56] & S37jy6);
assign S37jy6 = (~(Uy2jy6 & Sb5jy6));
assign Gzk7x6 = (G5j7z6[57] & A47jy6);
assign A47jy6 = (~(Mbj7x6 & Sb5jy6));
assign Vmu7x6 = (!Lgj7z6[171]);
assign Cnu7x6 = (!Lgj7z6[168]);
assign Ot6jy6 = (Uy6jy6 ? A0v7x6 : H0v7x6);
assign Uy6jy6 = (~(I47jy6 & Q47jy6));
assign Q47jy6 = (~(Y47jy6 & G5j7z6[58]));
assign Y47jy6 = (L2v7x6 & Sz6jy6);
assign Sz6jy6 = (~(Nfj7x6 & Sb5jy6));
assign L2v7x6 = (G57jy6 & O57jy6);
assign O57jy6 = (~(W57jy6 & Lgj7z6[175]));
assign W57jy6 = (E67jy6 & Cz6jy6);
assign Cz6jy6 = (!Lgj7z6[178]);
assign G57jy6 = (M67jy6 & U67jy6);
assign U67jy6 = (~(C77jy6 & K77jy6));
assign K77jy6 = (S77jy6 & H0v7x6);
assign S77jy6 = (~(Lgj7z6[178] & Mz88x6));
assign Mz88x6 = (!Lgj7z6[175]);
assign C77jy6 = (Lgj7z6[174] & E67jy6);
assign E67jy6 = (~(Lgj7z6[179] & V0v7x6));
assign V0v7x6 = (!Lgj7z6[176]);
assign M67jy6 = (~(Lgj7z6[176] & O0v7x6));
assign O0v7x6 = (!Lgj7z6[179]);
assign I47jy6 = (~(B7l7x6 & I07jy6));
assign I07jy6 = (So2nv6 | Sb5jy6);
assign Sb5jy6 = (A87jy6 & Xxjov6);
assign So2nv6 = (!G5j7z6[59]);
assign B7l7x6 = (~(G5j7z6[59] & Pfk7x6));
assign A0v7x6 = (!Lgj7z6[174]);
assign H0v7x6 = (!Lgj7z6[177]);
assign Me4jy6 = (Io4jy6 ? Q87jy6 : I87jy6);
assign Io4jy6 = (~(Y87jy6 | W54jy6));
assign W54jy6 = (~(G97jy6 | O97jy6));
assign G97jy6 = (W97jy6 | Ea7jy6);
assign Y87jy6 = (Ma7jy6 & Ua7jy6);
assign Ua7jy6 = (Cb7jy6 & Kb7jy6);
assign Kb7jy6 = (~(Sb7jy6 & Q87jy6));
assign Sb7jy6 = (Ac7jy6 & Ic7jy6);
assign Ac7jy6 = (Ao4jy6 | Qc7jy6);
assign Qc7jy6 = (!Sn4jy6);
assign Cb7jy6 = (Yc7jy6 | Sn4jy6);
assign Sn4jy6 = (Wd7jy6 ? Od7jy6 : Gd7jy6);
assign Yc7jy6 = (~(Ao4jy6 & Ic7jy6));
assign Ic7jy6 = (~(Mm4jy6 & Em4jy6));
assign Ao4jy6 = (Ue7jy6 ? Me7jy6 : Ee7jy6);
assign Ma7jy6 = (Cf7jy6 & Kf7jy6);
assign Kf7jy6 = (~(Op4jy6 & Wp4jy6));
assign Cf7jy6 = (Em4jy6 | Mm4jy6);
assign Mm4jy6 = (Wd7jy6 ? Ag7jy6 : Sf7jy6);
assign Wd7jy6 = (!Wp4jy6);
assign Em4jy6 = (!Ig7jy6);
assign Ig7jy6 = (Ue7jy6 ? Yg7jy6 : Qg7jy6);
assign Q87jy6 = (Ue7jy6 ? Oh7jy6 : Gh7jy6);
assign Ue7jy6 = (W97jy6 & Wh7jy6);
assign Wh7jy6 = (~(Ei7jy6 & Mi7jy6));
assign Mi7jy6 = (Ui7jy6 | Qg7jy6);
assign Ei7jy6 = (Cj7jy6 & Kj7jy6);
assign Kj7jy6 = (~(Yg7jy6 & Sj7jy6));
assign Sj7jy6 = (~(Qg7jy6 & Ui7jy6));
assign Ui7jy6 = (~(Ak7jy6 & Ik7jy6));
assign Ik7jy6 = (~(Ee7jy6 & Qk7jy6));
assign Qk7jy6 = (Yk7jy6 | Gh7jy6);
assign Ee7jy6 = (Wl7jy6 ? Ol7jy6 : Gl7jy6);
assign Ak7jy6 = (~(Gh7jy6 & Yk7jy6));
assign Yk7jy6 = (!Me7jy6);
assign Me7jy6 = (Um7jy6 ? Mm7jy6 : Em7jy6);
assign Qg7jy6 = (Wl7jy6 ? Kn7jy6 : Cn7jy6);
assign Cn7jy6 = (!Sn7jy6);
assign Yg7jy6 = (Um7jy6 ? Io7jy6 : Ao7jy6);
assign Cj7jy6 = (O97jy6 | Wl7jy6);
assign W97jy6 = (~(Qo7jy6 & Yo7jy6));
assign Yo7jy6 = (Gp7jy6 & Op7jy6);
assign Gp7jy6 = (~(Wp7jy6 | Eq7jy6));
assign Oh7jy6 = (Mq7jy6 | Uq7jy6);
assign Uq7jy6 = (Cr7jy6 & Kr7jy6);
assign Kr7jy6 = (Is7jy6 ? As7jy6 : Sr7jy6);
assign As7jy6 = (Qs7jy6 ? Myv7x6 : Q88iw6);
assign Myv7x6 = (!Lgj7z6[111]);
assign Q88iw6 = (!Lgj7z6[108]);
assign Cr7jy6 = (~(Ys7jy6 | Um7jy6));
assign Mq7jy6 = (Um7jy6 ? Ot7jy6 : Gt7jy6);
assign Um7jy6 = (Wt7jy6 & Eq7jy6);
assign Eq7jy6 = (~(Eu7jy6 & Mu7jy6));
assign Eu7jy6 = (~(Uu7jy6 | Cv7jy6));
assign Wt7jy6 = (~(Kv7jy6 & Sv7jy6));
assign Sv7jy6 = (~(Io7jy6 & Aw7jy6));
assign Kv7jy6 = (Iw7jy6 & Qw7jy6);
assign Qw7jy6 = (~(Qo7jy6 & Yw7jy6));
assign Yw7jy6 = (Op7jy6 & Gx7jy6);
assign Qo7jy6 = (~(Ox7jy6 | Wx7jy6));
assign Iw7jy6 = (Ao7jy6 | Ey7jy6);
assign Ey7jy6 = (~(Aw7jy6 | Io7jy6));
assign Io7jy6 = (Cz7jy6 ? Uy7jy6 : My7jy6);
assign Uy7jy6 = (!Kz7jy6);
assign Aw7jy6 = (~(Sz7jy6 & A08jy6));
assign A08jy6 = (~(Mm7jy6 & I08jy6));
assign I08jy6 = (Ot7jy6 | Q08jy6);
assign Mm7jy6 = (Cz7jy6 ? G18jy6 : Y08jy6);
assign Sz7jy6 = (~(Q08jy6 & Ot7jy6));
assign Q08jy6 = (!Em7jy6);
assign Em7jy6 = (Ys7jy6 ? W18jy6 : O18jy6);
assign Ao7jy6 = (Ys7jy6 ? M28jy6 : E28jy6);
assign M28jy6 = (!U28jy6);
assign Ot7jy6 = (Cz7jy6 ? K38jy6 : C38jy6);
assign Cz7jy6 = (S38jy6 & Cv7jy6);
assign Cv7jy6 = (A48jy6 | I48jy6);
assign S38jy6 = (~(Q48jy6 & Y48jy6));
assign Y48jy6 = (~(Mu7jy6 & G58jy6));
assign Q48jy6 = (O58jy6 & W58jy6);
assign W58jy6 = (~(E68jy6 & M68jy6));
assign M68jy6 = (~(My7jy6 & Kz7jy6));
assign E68jy6 = (U68jy6 & C78jy6);
assign C78jy6 = (G18jy6 | K78jy6);
assign K78jy6 = (~(Y08jy6 | C38jy6));
assign G18jy6 = (I88jy6 ? A88jy6 : S78jy6);
assign A88jy6 = (!Q88jy6);
assign U68jy6 = (~(C38jy6 & Y08jy6));
assign Y08jy6 = (G58jy6 ? G98jy6 : Y88jy6);
assign O58jy6 = (Kz7jy6 | My7jy6);
assign My7jy6 = (G58jy6 ? W98jy6 : O98jy6);
assign Kz7jy6 = (Ua8jy6 ? Ma8jy6 : Ea8jy6);
assign Ea8jy6 = (!Cb8jy6);
assign K38jy6 = (!Kb8jy6);
assign Kb8jy6 = (I88jy6 ? Ac8jy6 : Sb8jy6);
assign I88jy6 = (!Ua8jy6);
assign Ua8jy6 = (Ic8jy6 & I48jy6);
assign I48jy6 = (~(Qc8jy6 & Yc8jy6));
assign Yc8jy6 = (~(G5j7z6[47] & Ue6jy6));
assign Qc8jy6 = (Gd8jy6 & Od8jy6);
assign Od8jy6 = (X13nv6 | Qjk7x6);
assign X13nv6 = (H5iov6 & Itk7x6);
assign Itk7x6 = (!G5j7z6[46]);
assign H5iov6 = (!G5j7z6[47]);
assign Gd8jy6 = (~(G5j7z6[46] & Erk7x6));
assign Ic8jy6 = (~(Wd8jy6 & Ee8jy6));
assign Ee8jy6 = (Me8jy6 & A48jy6);
assign A48jy6 = (~(Ue8jy6 & Cf8jy6));
assign Cf8jy6 = (~(G5j7z6[45] & Ktl7x6));
assign Ue8jy6 = (Kf8jy6 & Sf8jy6);
assign Sf8jy6 = (Q13nv6 | Qjk7x6);
assign Q13nv6 = (Apk7x6 & Glk7x6);
assign Glk7x6 = (!G5j7z6[44]);
assign Apk7x6 = (!G5j7z6[45]);
assign Kf8jy6 = (~(G5j7z6[44] & Qpl7x6));
assign Me8jy6 = (~(Ag8jy6 & Ig8jy6));
assign Ig8jy6 = (Qg8jy6 ? Guw7x6 : Nuw7x6);
assign Guw7x6 = (!Lgj7z6[138]);
assign Ag8jy6 = (Yg8jy6 & Gh8jy6);
assign Gh8jy6 = (S78jy6 | Q88jy6);
assign Wd8jy6 = (Oh8jy6 & Wh8jy6);
assign Wh8jy6 = (~(Ei8jy6 & Q88jy6));
assign Q88jy6 = (Mi8jy6 ? Lgj7z6[136] : Lgj7z6[133]);
assign Ei8jy6 = (S78jy6 & Yg8jy6);
assign Yg8jy6 = (~(Ma8jy6 & Cb8jy6));
assign S78jy6 = (Qg8jy6 ? Dww7x6 : Wvw7x6);
assign Oh8jy6 = (Cb8jy6 | Ma8jy6);
assign Ma8jy6 = (Qg8jy6 ? Lgj7z6[140] : Lgj7z6[143]);
assign Cb8jy6 = (Mi8jy6 ? Pvw7x6 : Ub7iw6);
assign Ub7iw6 = (!Lgj7z6[134]);
assign Ac8jy6 = (Mi8jy6 ? Lgj7z6[135] : Lgj7z6[132]);
assign Mi8jy6 = (Ui8jy6 & G5j7z6[45]);
assign Ui8jy6 = (Cj8jy6 & Kj8jy6);
assign Kj8jy6 = (~(Sj8jy6 & Vyw7x6));
assign Vyw7x6 = (Ak8jy6 & Ik8jy6);
assign Ik8jy6 = (~(Lgj7z6[134] & Pvw7x6));
assign Ak8jy6 = (Qk8jy6 & Yk8jy6);
assign Yk8jy6 = (~(Gl8jy6 & Ol8jy6));
assign Ol8jy6 = (Wl8jy6 & Ltw7x6);
assign Ltw7x6 = (!Lgj7z6[135]);
assign Gl8jy6 = (Lgj7z6[132] & Em8jy6);
assign Em8jy6 = (~(Lgj7z6[136] & Yr7iw6));
assign Yr7iw6 = (!Lgj7z6[133]);
assign Qk8jy6 = (~(Mm8jy6 & Lgj7z6[133]));
assign Mm8jy6 = (Wl8jy6 & Txw7x6);
assign Txw7x6 = (!Lgj7z6[136]);
assign Wl8jy6 = (Pvw7x6 | Lgj7z6[134]);
assign Pvw7x6 = (!Lgj7z6[137]);
assign Sj8jy6 = (G5j7z6[44] & Um8jy6);
assign Um8jy6 = (~(Qjk7x6 & L1i7x6));
assign Cj8jy6 = (~(Qjk7x6 & Jrj7x6));
assign Sb8jy6 = (Qg8jy6 ? Lgj7z6[138] : Lgj7z6[141]);
assign Qg8jy6 = (~(Cn8jy6 & G5j7z6[47]));
assign Cn8jy6 = (Kn8jy6 & Sn8jy6);
assign Sn8jy6 = (~(Ao8jy6 & Fxw7x6));
assign Fxw7x6 = (Io8jy6 & Qo8jy6);
assign Qo8jy6 = (~(Lgj7z6[140] & Uuw7x6));
assign Uuw7x6 = (!Lgj7z6[143]);
assign Io8jy6 = (Yo8jy6 & Gp8jy6);
assign Gp8jy6 = (~(Op8jy6 & Wp8jy6));
assign Wp8jy6 = (Eq8jy6 & Nuw7x6);
assign Nuw7x6 = (!Lgj7z6[141]);
assign Eq8jy6 = (~(Lgj7z6[142] & Dww7x6));
assign Dww7x6 = (!Lgj7z6[139]);
assign Op8jy6 = (Lgj7z6[138] & Mq8jy6);
assign Yo8jy6 = (~(Uq8jy6 & Lgj7z6[139]));
assign Uq8jy6 = (Mq8jy6 & Wvw7x6);
assign Wvw7x6 = (!Lgj7z6[142]);
assign Mq8jy6 = (~(Lgj7z6[143] & Bvw7x6));
assign Bvw7x6 = (!Lgj7z6[140]);
assign Ao8jy6 = (G5j7z6[46] & Cr8jy6);
assign Cr8jy6 = (~(Qjk7x6 & P3i7x6));
assign Kn8jy6 = (~(Qjk7x6 & V6i7x6));
assign C38jy6 = (G58jy6 ? Sr8jy6 : Kr8jy6);
assign G58jy6 = (~(As8jy6 & Uu7jy6));
assign Uu7jy6 = (~(Is8jy6 & Qs8jy6));
assign Qs8jy6 = (~(G5j7z6[43] & Pfk7x6));
assign Is8jy6 = (Ys8jy6 & Gt8jy6);
assign Gt8jy6 = (J13nv6 | Qjk7x6);
assign J13nv6 = (Fhk7x6 & Edk7x6);
assign Edk7x6 = (!G5j7z6[42]);
assign Fhk7x6 = (!G5j7z6[43]);
assign Ys8jy6 = (~(G5j7z6[42] & O3l7x6));
assign As8jy6 = (~(Ot8jy6 & Wt8jy6));
assign Wt8jy6 = (~(Eu8jy6 | Mu7jy6));
assign Mu7jy6 = (Mu8jy6 & Uu8jy6);
assign Uu8jy6 = (~(G5j7z6[41] & U7k7x6));
assign Mu8jy6 = (Cv8jy6 & Kv8jy6);
assign Kv8jy6 = (B43nv6 | Qjk7x6);
assign B43nv6 = (K9k7x6 & Q5k7x6);
assign Q5k7x6 = (!G5j7z6[40]);
assign K9k7x6 = (!G5j7z6[41]);
assign Cv8jy6 = (~(G5j7z6[40] & T3k7x6));
assign Eu8jy6 = (Sv8jy6 & Kr8jy6);
assign Sv8jy6 = (Aw8jy6 & Iw8jy6);
assign Iw8jy6 = (~(Qw8jy6 & G98jy6));
assign Ot8jy6 = (Yw8jy6 & Gx8jy6);
assign Gx8jy6 = (Ox8jy6 | G98jy6);
assign G98jy6 = (Wx8jy6 ? M4x7x6 : Ts7iw6);
assign Ox8jy6 = (~(Y88jy6 & Aw8jy6));
assign Aw8jy6 = (O98jy6 | Ey8jy6);
assign Y88jy6 = (!Qw8jy6);
assign Qw8jy6 = (My8jy6 ? Lgj7z6[127] : Lgj7z6[130]);
assign Yw8jy6 = (~(Ey8jy6 & O98jy6));
assign O98jy6 = (My8jy6 ? Uy8jy6 : S478x6);
assign Ey8jy6 = (!W98jy6);
assign W98jy6 = (Wx8jy6 ? Vv68x6 : Wc7iw6);
assign Wc7iw6 = (!Lgj7z6[122]);
assign Sr8jy6 = (Wx8jy6 ? Rpw7x6 : O78iw6);
assign Wx8jy6 = (Cz8jy6 & G5j7z6[41]);
assign Cz8jy6 = (Kz8jy6 & Sz8jy6);
assign Sz8jy6 = (~(A09jy6 & O5x7x6));
assign O5x7x6 = (I09jy6 & Q09jy6);
assign Q09jy6 = (~(Lgj7z6[122] & Vv68x6));
assign I09jy6 = (Y09jy6 & G19jy6);
assign G19jy6 = (~(O19jy6 & W19jy6));
assign W19jy6 = (E29jy6 & Rpw7x6);
assign O19jy6 = (Lgj7z6[120] & M29jy6);
assign M29jy6 = (~(Lgj7z6[124] & Ts7iw6));
assign Ts7iw6 = (!Lgj7z6[121]);
assign Y09jy6 = (~(U29jy6 & Lgj7z6[121]));
assign U29jy6 = (E29jy6 & M4x7x6);
assign M4x7x6 = (!Lgj7z6[124]);
assign E29jy6 = (Vv68x6 | Lgj7z6[122]);
assign Vv68x6 = (!Lgj7z6[125]);
assign A09jy6 = (G5j7z6[40] & C39jy6);
assign C39jy6 = (~(Qjk7x6 & Uy2jy6));
assign Kz8jy6 = (~(Qjk7x6 & Mbj7x6));
assign Rpw7x6 = (!Lgj7z6[123]);
assign O78iw6 = (!Lgj7z6[120]);
assign Kr8jy6 = (My8jy6 ? Y3x7x6 : R3x7x6);
assign My8jy6 = (~(K39jy6 & G5j7z6[43]));
assign K39jy6 = (S39jy6 & A49jy6);
assign A49jy6 = (~(I49jy6 & L7x7x6));
assign L7x7x6 = (Q49jy6 & Y49jy6);
assign Y49jy6 = (~(G59jy6 & Lgj7z6[127]));
assign G59jy6 = (O59jy6 & C6x7x6);
assign C6x7x6 = (!Lgj7z6[130]);
assign Q49jy6 = (W59jy6 & E69jy6);
assign E69jy6 = (~(M69jy6 & U69jy6));
assign U69jy6 = (C79jy6 & R3x7x6);
assign C79jy6 = (~(Lgj7z6[130] & J6x7x6));
assign J6x7x6 = (!Lgj7z6[127]);
assign M69jy6 = (Lgj7z6[126] & O59jy6);
assign O59jy6 = (~(Lgj7z6[131] & Uy8jy6));
assign Uy8jy6 = (!Lgj7z6[128]);
assign W59jy6 = (~(Lgj7z6[128] & S478x6));
assign S478x6 = (!Lgj7z6[131]);
assign I49jy6 = (G5j7z6[42] & K79jy6);
assign K79jy6 = (~(Qjk7x6 & Nfj7x6));
assign S39jy6 = (~(Qjk7x6 & Hzh7x6));
assign Y3x7x6 = (!Lgj7z6[126]);
assign R3x7x6 = (!Lgj7z6[129]);
assign Gt7jy6 = (S79jy6 & Ys7jy6);
assign Ys7jy6 = (~(A89jy6 & I89jy6));
assign I89jy6 = (~(Q89jy6 & Y89jy6));
assign Y89jy6 = (Wx7jy6 | G99jy6);
assign Q89jy6 = (O99jy6 & W99jy6);
assign W99jy6 = (~(Ea9jy6 & Ma9jy6));
assign Ma9jy6 = (U28jy6 | E28jy6);
assign Ea9jy6 = (Ua9jy6 & Cb9jy6);
assign Cb9jy6 = (O18jy6 | Kb9jy6);
assign Kb9jy6 = (!Sb9jy6);
assign Sb9jy6 = (S79jy6 | W18jy6);
assign O18jy6 = (Is7jy6 ? Ic9jy6 : Ac9jy6);
assign Ic9jy6 = (!Qc9jy6);
assign Ua9jy6 = (~(W18jy6 & S79jy6));
assign W18jy6 = (G99jy6 ? Gd9jy6 : Yc9jy6);
assign O99jy6 = (~(E28jy6 & U28jy6));
assign U28jy6 = (G99jy6 ? Wd9jy6 : Od9jy6);
assign E28jy6 = (Is7jy6 ? Me9jy6 : Ee9jy6);
assign Is7jy6 = (~(Ue9jy6 & Wp7jy6));
assign Wp7jy6 = (!Gx7jy6);
assign Ue9jy6 = (~(Cf9jy6 & Kf9jy6));
assign Kf9jy6 = (~(Sf9jy6 | Op7jy6));
assign Sf9jy6 = (Ag9jy6 & Sr7jy6);
assign Sr7jy6 = (Ig9jy6 ? A6w7x6 : T5w7x6);
assign T5w7x6 = (!Lgj7z6[114]);
assign Ag9jy6 = (Qg9jy6 & Yg9jy6);
assign Yg9jy6 = (Ac9jy6 | Qc9jy6);
assign Cf9jy6 = (Gh9jy6 & Oh9jy6);
assign Oh9jy6 = (~(Wh9jy6 & Qc9jy6));
assign Qc9jy6 = (Qs7jy6 ? Lgj7z6[112] : Lgj7z6[109]);
assign Wh9jy6 = (Ac9jy6 & Qg9jy6);
assign Qg9jy6 = (~(Ei9jy6 & Me9jy6));
assign Ac9jy6 = (Ig9jy6 ? Mi9jy6 : Qi68x6);
assign Gh9jy6 = (Me9jy6 | Ei9jy6);
assign Ei9jy6 = (!Ee9jy6);
assign Me9jy6 = (Qs7jy6 ? V6w7x6 : Yd7iw6);
assign Qs7jy6 = (Ui9jy6 & G5j7z6[37]);
assign Ui9jy6 = (Cj9jy6 & Kj9jy6);
assign Kj9jy6 = (~(Sj9jy6 & E8w7x6));
assign E8w7x6 = (Ak9jy6 & Ik9jy6);
assign Ik9jy6 = (~(Lgj7z6[110] & V6w7x6));
assign Ak9jy6 = (Qk9jy6 & Yk9jy6);
assign Yk9jy6 = (~(Gl9jy6 & Ol9jy6));
assign Ol9jy6 = (~(Wl9jy6 | Lgj7z6[111]));
assign Gl9jy6 = (Lgj7z6[108] & Em9jy6);
assign Em9jy6 = (~(Lgj7z6[112] & Ot7iw6));
assign Ot7iw6 = (!Lgj7z6[109]);
assign Qk9jy6 = (~(Mm9jy6 & Lgj7z6[109]));
assign Mm9jy6 = (~(Wl9jy6 | Lgj7z6[112]));
assign Wl9jy6 = (Lgj7z6[113] & Yd7iw6);
assign Sj9jy6 = (G5j7z6[36] & Um9jy6);
assign Um9jy6 = (~(Qjk7x6 & Cshov6));
assign Cj9jy6 = (~(Qjk7x6 & I2oiw6));
assign V6w7x6 = (!Lgj7z6[113]);
assign Yd7iw6 = (!Lgj7z6[110]);
assign Ee9jy6 = (Ig9jy6 ? O6w7x6 : H6w7x6);
assign Ig9jy6 = (Cn9jy6 & G5j7z6[39]);
assign Cn9jy6 = (Kn9jy6 & Sn9jy6);
assign Sn9jy6 = (~(Ao9jy6 & G9w7x6));
assign G9w7x6 = (Io9jy6 & Qo9jy6);
assign Qo9jy6 = (~(Yo9jy6 & Lgj7z6[115]));
assign Yo9jy6 = (Gp9jy6 & Mi9jy6);
assign Mi9jy6 = (!Lgj7z6[118]);
assign Io9jy6 = (Op9jy6 & Wp9jy6);
assign Wp9jy6 = (~(Eq9jy6 & Mq9jy6));
assign Mq9jy6 = (Uq9jy6 & A6w7x6);
assign A6w7x6 = (!Lgj7z6[117]);
assign Uq9jy6 = (~(Lgj7z6[118] & Qi68x6));
assign Qi68x6 = (!Lgj7z6[115]);
assign Eq9jy6 = (Lgj7z6[114] & Gp9jy6);
assign Gp9jy6 = (~(Lgj7z6[119] & H6w7x6));
assign Op9jy6 = (~(Lgj7z6[116] & O6w7x6));
assign Ao9jy6 = (G5j7z6[38] & Cr9jy6);
assign Cr9jy6 = (~(Qjk7x6 & Rphov6));
assign Kn9jy6 = (~(Qjk7x6 & J6oiw6));
assign O6w7x6 = (!Lgj7z6[119]);
assign H6w7x6 = (!Lgj7z6[116]);
assign A89jy6 = (~(Op7jy6 & Gx7jy6));
assign Gx7jy6 = (Kr9jy6 & Sr9jy6);
assign Sr9jy6 = (~(G5j7z6[39] & Ua5jy6));
assign Kr9jy6 = (As9jy6 & Is9jy6);
assign Is9jy6 = (U33nv6 | Qjk7x6);
assign U33nv6 = (Bnoiw6 & I3niw6);
assign I3niw6 = (!G5j7z6[38]);
assign Bnoiw6 = (!G5j7z6[39]);
assign As9jy6 = (~(G5j7z6[38] & Ac5jy6));
assign Op7jy6 = (Qs9jy6 & Ys9jy6);
assign Ys9jy6 = (~(G5j7z6[37] & Wd5jy6));
assign Qs9jy6 = (Gt9jy6 & Ot9jy6);
assign Ot9jy6 = (N33nv6 | Qjk7x6);
assign N33nv6 = (Ajoiw6 & Vzmiw6);
assign Vzmiw6 = (!G5j7z6[36]);
assign Ajoiw6 = (!G5j7z6[37]);
assign Gt9jy6 = (~(G5j7z6[36] & Ue5jy6));
assign S79jy6 = (G99jy6 ? Eu9jy6 : Wt9jy6);
assign G99jy6 = (Mu9jy6 & Ox7jy6);
assign Ox7jy6 = (~(Uu9jy6 & Cv9jy6));
assign Cv9jy6 = (~(G5j7z6[35] & Xdoiw6));
assign Uu9jy6 = (Kv9jy6 & Sv9jy6);
assign Sv9jy6 = (W43nv6 | Qjk7x6);
assign W43nv6 = (Nfoiw6 & Aw9jy6);
assign Aw9jy6 = (!G5j7z6[34]);
assign Nfoiw6 = (!G5j7z6[35]);
assign Kv9jy6 = (~(G5j7z6[34] & Zumiw6));
assign Mu9jy6 = (~(Iw9jy6 & Qw9jy6));
assign Qw9jy6 = (Yw9jy6 & Wx7jy6);
assign Wx7jy6 = (~(Gx9jy6 & Ox9jy6));
assign Ox9jy6 = (~(G5j7z6[33] & Daoiw6));
assign Gx9jy6 = (Wx9jy6 & Ey9jy6);
assign Ey9jy6 = (D53nv6 | Qjk7x6);
assign D53nv6 = (Tboiw6 & Hsmiw6);
assign Hsmiw6 = (!G5j7z6[32]);
assign Tboiw6 = (!G5j7z6[33]);
assign Wx9jy6 = (~(G5j7z6[32] & Rqmiw6));
assign Yw9jy6 = (~(My9jy6 & Eu9jy6));
assign My9jy6 = (Uy9jy6 & Cz9jy6);
assign Cz9jy6 = (~(Kz9jy6 & Yc9jy6));
assign Iw9jy6 = (Sz9jy6 & A0ajy6);
assign A0ajy6 = (I0ajy6 | Yc9jy6);
assign Yc9jy6 = (Q0ajy6 ? Efw7x6 : Ju7iw6);
assign I0ajy6 = (~(Gd9jy6 & Uy9jy6));
assign Uy9jy6 = (Y0ajy6 | Od9jy6);
assign Gd9jy6 = (!Kz9jy6);
assign Kz9jy6 = (G1ajy6 ? Lgj7z6[103] : Lgj7z6[106]);
assign Sz9jy6 = (~(Od9jy6 & Y0ajy6));
assign Y0ajy6 = (!Wd9jy6);
assign Wd9jy6 = (G1ajy6 ? Lgj7z6[104] : Lgj7z6[107]);
assign Od9jy6 = (Q0ajy6 ? Lgj7z6[101] : Lgj7z6[98]);
assign Eu9jy6 = (G1ajy6 ? Qew7x6 : Jew7x6);
assign G1ajy6 = (~(O1ajy6 & G5j7z6[35]));
assign O1ajy6 = (W1ajy6 & E2ajy6);
assign E2ajy6 = (~(M2ajy6 & Diw7x6));
assign Diw7x6 = (U2ajy6 & C3ajy6);
assign C3ajy6 = (~(K3ajy6 & Lgj7z6[103]));
assign K3ajy6 = (S3ajy6 & Ugw7x6);
assign Ugw7x6 = (!Lgj7z6[106]);
assign U2ajy6 = (A4ajy6 & I4ajy6);
assign I4ajy6 = (~(Q4ajy6 & Y4ajy6));
assign Y4ajy6 = (G5ajy6 & Jew7x6);
assign G5ajy6 = (~(Lgj7z6[106] & Bhw7x6));
assign Bhw7x6 = (!Lgj7z6[103]);
assign Q4ajy6 = (Lgj7z6[102] & S3ajy6);
assign S3ajy6 = (~(Lgj7z6[107] & O5ajy6));
assign O5ajy6 = (!Lgj7z6[104]);
assign A4ajy6 = (~(Lgj7z6[104] & L568x6));
assign L568x6 = (!Lgj7z6[107]);
assign M2ajy6 = (G5j7z6[34] & W5ajy6);
assign W5ajy6 = (~(Qjk7x6 & Jfmiw6));
assign W1ajy6 = (~(Qjk7x6 & Cn2jy6));
assign Qew7x6 = (!Lgj7z6[102]);
assign Jew7x6 = (!Lgj7z6[105]);
assign Wt9jy6 = (Q0ajy6 ? J0w7x6 : Ua8iw6);
assign Q0ajy6 = (E6ajy6 & G5j7z6[33]);
assign E6ajy6 = (M6ajy6 & U6ajy6);
assign U6ajy6 = (~(C7ajy6 & Ggw7x6));
assign Ggw7x6 = (K7ajy6 & S7ajy6);
assign S7ajy6 = (~(Lgj7z6[98] & Ow58x6));
assign K7ajy6 = (A8ajy6 & I8ajy6);
assign I8ajy6 = (~(Q8ajy6 & Y8ajy6));
assign Y8ajy6 = (G9ajy6 & J0w7x6);
assign Q8ajy6 = (Lgj7z6[96] & O9ajy6);
assign O9ajy6 = (~(Lgj7z6[100] & Ju7iw6));
assign Ju7iw6 = (!Lgj7z6[97]);
assign A8ajy6 = (~(W9ajy6 & Lgj7z6[97]));
assign W9ajy6 = (G9ajy6 & Efw7x6);
assign Efw7x6 = (!Lgj7z6[100]);
assign G9ajy6 = (Ow58x6 | Lgj7z6[98]);
assign Ow58x6 = (!Lgj7z6[101]);
assign C7ajy6 = (G5j7z6[32] & Eaajy6);
assign Eaajy6 = (~(Qjk7x6 & Ao2jy6));
assign M6ajy6 = (~(Qjk7x6 & Nuniw6));
assign Qjk7x6 = (Maajy6 & Xxjov6);
assign J0w7x6 = (!Lgj7z6[99]);
assign Ua8iw6 = (!Lgj7z6[96]);
assign Gh7jy6 = (~(Uaajy6 | Cbajy6));
assign Cbajy6 = (~(Kbajy6 | Wl7jy6));
assign Kbajy6 = (Icajy6 ? Acajy6 : Sbajy6);
assign Acajy6 = (~(Qcajy6 & Ycajy6));
assign Ycajy6 = (Gdajy6 ? Lgj7z6[66] : Lgj7z6[69]);
assign Uaajy6 = (Wl7jy6 ? Wdajy6 : Odajy6);
assign Wl7jy6 = (Eeajy6 & Ea7jy6);
assign Ea7jy6 = (~(Meajy6 & Ueajy6));
assign Ueajy6 = (~(Cfajy6 | Kfajy6));
assign Meajy6 = (~(Sfajy6 | Agajy6));
assign Eeajy6 = (~(Igajy6 & Qgajy6));
assign Qgajy6 = (Ygajy6 & O97jy6);
assign O97jy6 = (~(Ghajy6 & Ohajy6));
assign Ohajy6 = (Whajy6 & Eiajy6);
assign Whajy6 = (Miajy6 & Uiajy6);
assign Ghajy6 = (~(Cjajy6 | Kjajy6));
assign Ygajy6 = (~(Ol7jy6 & Sjajy6));
assign Sjajy6 = (~(Akajy6 & Ikajy6));
assign Ikajy6 = (Wdajy6 | Qkajy6);
assign Ol7jy6 = (Olajy6 ? Glajy6 : Ykajy6);
assign Ykajy6 = (!Wlajy6);
assign Igajy6 = (Emajy6 & Mmajy6);
assign Mmajy6 = (Akajy6 | Wdajy6);
assign Akajy6 = (Gl7jy6 | Qkajy6);
assign Qkajy6 = (~(Sn7jy6 | Kn7jy6));
assign Gl7jy6 = (Icajy6 ? Cnajy6 : Umajy6);
assign Emajy6 = (~(Kn7jy6 & Sn7jy6));
assign Sn7jy6 = (Icajy6 ? Snajy6 : Knajy6);
assign Kn7jy6 = (Olajy6 ? Ioajy6 : Aoajy6);
assign Wdajy6 = (Olajy6 ? Yoajy6 : Qoajy6);
assign Olajy6 = (Gpajy6 & Opajy6);
assign Opajy6 = (~(Wpajy6 & Eqajy6));
assign Eqajy6 = (Sfajy6 | Mqajy6);
assign Wpajy6 = (Uqajy6 & Crajy6);
assign Crajy6 = (~(Ioajy6 & Krajy6));
assign Krajy6 = (Srajy6 | Asajy6);
assign Ioajy6 = (Ysajy6 ? Qsajy6 : Isajy6);
assign Uqajy6 = (~(Asajy6 & Srajy6));
assign Srajy6 = (!Aoajy6);
assign Aoajy6 = (Mqajy6 ? Otajy6 : Gtajy6);
assign Asajy6 = (Wtajy6 & Euajy6);
assign Euajy6 = (~(Muajy6 & Uuajy6));
assign Uuajy6 = (~(Wlajy6 & Glajy6));
assign Wtajy6 = (Glajy6 | Wlajy6);
assign Wlajy6 = (Mqajy6 ? Kvajy6 : Cvajy6);
assign Kvajy6 = (!Svajy6);
assign Glajy6 = (Ysajy6 ? Iwajy6 : Awajy6);
assign Awajy6 = (!Qwajy6);
assign Gpajy6 = (Cfajy6 | Kfajy6);
assign Yoajy6 = (Ysajy6 ? Gxajy6 : Ywajy6);
assign Ysajy6 = (Oxajy6 & Kfajy6);
assign Kfajy6 = (~(Wxajy6 & Eyajy6));
assign Eyajy6 = (~(G5j7z6[31] & Ue6jy6));
assign Wxajy6 = (Myajy6 & Uyajy6);
assign Uyajy6 = (Ry2nv6 | Czajy6);
assign Ry2nv6 = (B1k7x6 & Twj7x6);
assign Twj7x6 = (!G5j7z6[30]);
assign B1k7x6 = (!G5j7z6[31]);
assign Myajy6 = (~(G5j7z6[30] & Erk7x6));
assign Oxajy6 = (~(Kzajy6 & Szajy6));
assign Szajy6 = (A0bjy6 & Cfajy6);
assign Cfajy6 = (~(I0bjy6 & Q0bjy6));
assign Q0bjy6 = (~(G5j7z6[29] & Ktl7x6));
assign I0bjy6 = (Y0bjy6 & G1bjy6);
assign G1bjy6 = (~(V03nv6 & Inj7x6));
assign V03nv6 = (~(Zsj7x6 & Yoj7x6));
assign Yoj7x6 = (!G5j7z6[28]);
assign Zsj7x6 = (!G5j7z6[29]);
assign Y0bjy6 = (~(G5j7z6[28] & Qpl7x6));
assign A0bjy6 = (~(O1bjy6 & W1bjy6));
assign W1bjy6 = (E2bjy6 ? Xrx7x6 : Esx7x6);
assign Xrx7x6 = (!Lgj7z6[90]);
assign O1bjy6 = (M2bjy6 & U2bjy6);
assign U2bjy6 = (Iwajy6 | Qwajy6);
assign Kzajy6 = (C3bjy6 & K3bjy6);
assign K3bjy6 = (~(S3bjy6 & Qwajy6));
assign Qwajy6 = (A4bjy6 ? Lgj7z6[88] : Lgj7z6[85]);
assign S3bjy6 = (Iwajy6 & M2bjy6);
assign M2bjy6 = (~(I4bjy6 & Isajy6));
assign Iwajy6 = (E2bjy6 ? Cj58x6 : Q4bjy6);
assign C3bjy6 = (Isajy6 | I4bjy6);
assign I4bjy6 = (!Qsajy6);
assign Qsajy6 = (E2bjy6 ? Y4bjy6 : Rn58x6);
assign Isajy6 = (A4bjy6 ? T16iw6 : G5bjy6);
assign G5bjy6 = (!Lgj7z6[86]);
assign Gxajy6 = (E2bjy6 ? Lgj7z6[90] : Lgj7z6[93]);
assign E2bjy6 = (~(O5bjy6 & G5j7z6[31]));
assign O5bjy6 = (W5bjy6 & E6bjy6);
assign E6bjy6 = (~(M6bjy6 & Wux7x6));
assign Wux7x6 = (U6bjy6 & C7bjy6);
assign C7bjy6 = (~(K7bjy6 & Lgj7z6[91]));
assign K7bjy6 = (S7bjy6 & Q4bjy6);
assign Q4bjy6 = (!Lgj7z6[94]);
assign U6bjy6 = (A8bjy6 & I8bjy6);
assign I8bjy6 = (~(Q8bjy6 & Y8bjy6));
assign Y8bjy6 = (G9bjy6 & Esx7x6);
assign Esx7x6 = (!Lgj7z6[93]);
assign G9bjy6 = (~(Lgj7z6[94] & Cj58x6));
assign Cj58x6 = (!Lgj7z6[91]);
assign Q8bjy6 = (Lgj7z6[90] & S7bjy6);
assign S7bjy6 = (~(Lgj7z6[95] & Y4bjy6));
assign Y4bjy6 = (!Lgj7z6[92]);
assign A8bjy6 = (~(Lgj7z6[92] & Rn58x6));
assign Rn58x6 = (!Lgj7z6[95]);
assign M6bjy6 = (G5j7z6[30] & O9bjy6);
assign O9bjy6 = (~(Czajy6 & P3i7x6));
assign W5bjy6 = (~(Czajy6 & V6i7x6));
assign Ywajy6 = (A4bjy6 ? Lgj7z6[87] : Lgj7z6[84]);
assign A4bjy6 = (W9bjy6 & G5j7z6[29]);
assign W9bjy6 = (Eabjy6 & Mabjy6);
assign Mabjy6 = (~(Uabjy6 & Ntx7x6));
assign Ntx7x6 = (Cbbjy6 & Kbbjy6);
assign Kbbjy6 = (~(Lgj7z6[86] & T16iw6));
assign Cbbjy6 = (Sbbjy6 & Acbjy6);
assign Acbjy6 = (~(Icbjy6 & Qcbjy6));
assign Qcbjy6 = (Ycbjy6 & Gq6iw6);
assign Gq6iw6 = (!Lgj7z6[87]);
assign Icbjy6 = (Lgj7z6[84] & Gdbjy6);
assign Gdbjy6 = (~(Lgj7z6[88] & Fa58x6));
assign Fa58x6 = (!Lgj7z6[85]);
assign Sbbjy6 = (~(Odbjy6 & Lgj7z6[85]));
assign Odbjy6 = (Ycbjy6 & Ff6iw6);
assign Ff6iw6 = (!Lgj7z6[88]);
assign Ycbjy6 = (T16iw6 | Lgj7z6[86]);
assign T16iw6 = (!Lgj7z6[89]);
assign Uabjy6 = (G5j7z6[28] & Wdbjy6);
assign Wdbjy6 = (~(Czajy6 & L1i7x6));
assign Eabjy6 = (~(Jrj7x6 & Czajy6));
assign Qoajy6 = (!Muajy6);
assign Muajy6 = (Mqajy6 ? Mebjy6 : Eebjy6);
assign Mqajy6 = (Uebjy6 & Agajy6);
assign Agajy6 = (~(Cfbjy6 & Kfbjy6));
assign Kfbjy6 = (~(G5j7z6[27] & Pfk7x6));
assign Cfbjy6 = (Sfbjy6 & Agbjy6);
assign Agbjy6 = (~(O03nv6 & Inj7x6));
assign O03nv6 = (~(Xkj7x6 & Dhj7x6));
assign Dhj7x6 = (!G5j7z6[26]);
assign Xkj7x6 = (!G5j7z6[27]);
assign Sfbjy6 = (~(G5j7z6[26] & O3l7x6));
assign O3l7x6 = (!Nfj7x6);
assign Uebjy6 = (~(Igbjy6 & Qgbjy6));
assign Qgbjy6 = (Ygbjy6 & Sfajy6);
assign Sfajy6 = (~(Ghbjy6 & Ohbjy6));
assign Ohbjy6 = (~(G5j7z6[25] & U7k7x6));
assign Ghbjy6 = (Whbjy6 & Eibjy6);
assign Eibjy6 = (H03nv6 | Czajy6);
assign H03nv6 = (Cdj7x6 & N8j7x6);
assign N8j7x6 = (!G5j7z6[24]);
assign Cdj7x6 = (!G5j7z6[25]);
assign Whbjy6 = (~(G5j7z6[24] & T3k7x6));
assign T3k7x6 = (!Uy2jy6);
assign Ygbjy6 = (~(Mibjy6 & Mebjy6));
assign Mibjy6 = (Uibjy6 & Cjbjy6);
assign Cjbjy6 = (Svajy6 | Cvajy6);
assign Igbjy6 = (Kjbjy6 & Sjbjy6);
assign Sjbjy6 = (~(Akbjy6 & Cvajy6));
assign Cvajy6 = (Ikbjy6 ? Lgj7z6[73] : Lgj7z6[76]);
assign Ikbjy6 = (!Qkbjy6);
assign Akbjy6 = (Svajy6 & Uibjy6);
assign Uibjy6 = (Otajy6 | Ykbjy6);
assign Svajy6 = (Glbjy6 ? R2y7x6 : K2y7x6);
assign Kjbjy6 = (~(Ykbjy6 & Otajy6));
assign Otajy6 = (Glbjy6 ? Olbjy6 : Q558x6);
assign Ykbjy6 = (!Gtajy6);
assign Gtajy6 = (Qkbjy6 ? Tw48x6 : Wlbjy6);
assign Wlbjy6 = (!Lgj7z6[74]);
assign Mebjy6 = (Glbjy6 ? Zzx7x6 : Szx7x6);
assign Glbjy6 = (~(Embjy6 & G5j7z6[27]));
assign Embjy6 = (Mmbjy6 & Umbjy6);
assign Umbjy6 = (~(Cnbjy6 & T3y7x6));
assign T3y7x6 = (Knbjy6 & Snbjy6);
assign Snbjy6 = (~(Lgj7z6[80] & Q558x6));
assign Q558x6 = (!Lgj7z6[83]);
assign Knbjy6 = (Aobjy6 & Iobjy6);
assign Iobjy6 = (~(Qobjy6 & Yobjy6));
assign Yobjy6 = (Gpbjy6 & Szx7x6);
assign Gpbjy6 = (~(Lgj7z6[82] & R2y7x6));
assign R2y7x6 = (!Lgj7z6[79]);
assign Qobjy6 = (Lgj7z6[78] & Opbjy6);
assign Aobjy6 = (~(Wpbjy6 & Lgj7z6[79]));
assign Wpbjy6 = (Opbjy6 & K2y7x6);
assign K2y7x6 = (!Lgj7z6[82]);
assign Opbjy6 = (~(Lgj7z6[83] & Olbjy6));
assign Olbjy6 = (!Lgj7z6[80]);
assign Cnbjy6 = (G5j7z6[26] & Eqbjy6);
assign Eqbjy6 = (~(Nfj7x6 & Czajy6));
assign Mmbjy6 = (~(Czajy6 & Hzh7x6));
assign Zzx7x6 = (!Lgj7z6[78]);
assign Szx7x6 = (!Lgj7z6[81]);
assign Eebjy6 = (Qkbjy6 ? Inx7x6 : Bnx7x6);
assign Qkbjy6 = (Mqbjy6 & G5j7z6[25]);
assign Mqbjy6 = (Uqbjy6 & Crbjy6);
assign Crbjy6 = (~(Krbjy6 & W1y7x6));
assign W1y7x6 = (Srbjy6 & Asbjy6);
assign Asbjy6 = (~(Lgj7z6[74] & Tw48x6));
assign Srbjy6 = (Isbjy6 & Qsbjy6);
assign Qsbjy6 = (~(Ysbjy6 & Gtbjy6));
assign Gtbjy6 = (Otbjy6 & Inx7x6);
assign Ysbjy6 = (Lgj7z6[72] & Wtbjy6);
assign Wtbjy6 = (~(Lgj7z6[76] & N0y7x6));
assign N0y7x6 = (!Lgj7z6[73]);
assign Isbjy6 = (~(Eubjy6 & Lgj7z6[73]));
assign Eubjy6 = (Otbjy6 & U0y7x6);
assign U0y7x6 = (!Lgj7z6[76]);
assign Otbjy6 = (Tw48x6 | Lgj7z6[74]);
assign Tw48x6 = (!Lgj7z6[77]);
assign Krbjy6 = (G5j7z6[24] & Mubjy6);
assign Mubjy6 = (~(Uy2jy6 & Czajy6));
assign Uqbjy6 = (~(Mbj7x6 & Czajy6));
assign Inx7x6 = (!Lgj7z6[75]);
assign Bnx7x6 = (!Lgj7z6[72]);
assign Odajy6 = (Uubjy6 & Icajy6);
assign Icajy6 = (Cvbjy6 & Kvbjy6);
assign Kvbjy6 = (~(Svbjy6 & Awbjy6));
assign Awbjy6 = (~(Miajy6 & Iwbjy6));
assign Miajy6 = (!Qwbjy6);
assign Svbjy6 = (Ywbjy6 & Gxbjy6);
assign Gxbjy6 = (Snajy6 | Oxbjy6);
assign Oxbjy6 = (~(Knajy6 | Wxbjy6));
assign Snajy6 = (Qcajy6 ? Mybjy6 : Eybjy6);
assign Qcajy6 = (!Uybjy6);
assign Mybjy6 = (!Czbjy6);
assign Ywbjy6 = (~(Wxbjy6 & Knajy6));
assign Knajy6 = (Iwbjy6 ? Szbjy6 : Kzbjy6);
assign Wxbjy6 = (~(A0cjy6 | I0cjy6));
assign I0cjy6 = (Umajy6 & Sbajy6);
assign A0cjy6 = (~(Cnajy6 | Q0cjy6));
assign Q0cjy6 = (~(Sbajy6 | Umajy6));
assign Umajy6 = (Iwbjy6 ? G1cjy6 : Y0cjy6);
assign G1cjy6 = (!O1cjy6);
assign Sbajy6 = (Iwbjy6 ? E2cjy6 : W1cjy6);
assign Iwbjy6 = (~(M2cjy6 & U2cjy6));
assign U2cjy6 = (~(C3cjy6 & K3cjy6));
assign K3cjy6 = (S3cjy6 & A4cjy6);
assign A4cjy6 = (~(I4cjy6 & W1cjy6));
assign I4cjy6 = (Q4cjy6 & Y4cjy6);
assign Q4cjy6 = (Y0cjy6 | O1cjy6);
assign S3cjy6 = (~(G5cjy6 & O1cjy6));
assign O1cjy6 = (O5cjy6 ? Lgj7z6[49] : Lgj7z6[52]);
assign O5cjy6 = (!W5cjy6);
assign G5cjy6 = (Y0cjy6 & Y4cjy6);
assign Y4cjy6 = (~(Kzbjy6 & E6cjy6));
assign Y0cjy6 = (M6cjy6 ? Oiy7x6 : Viy7x6);
assign C3cjy6 = (Qwbjy6 & U6cjy6);
assign U6cjy6 = (E6cjy6 | Kzbjy6);
assign Kzbjy6 = (M6cjy6 ? Lgj7z6[59] : Lgj7z6[56]);
assign E6cjy6 = (!Szbjy6);
assign Szbjy6 = (W5cjy6 ? Lgj7z6[53] : Lgj7z6[50]);
assign Qwbjy6 = (C7cjy6 & K7cjy6);
assign K7cjy6 = (~(S7cjy6 & Namiw6));
assign Namiw6 = (~(G5j7z6[16] & Rqmiw6));
assign C7cjy6 = (A8cjy6 | G5j7z6[17]);
assign M2cjy6 = (~(Uiajy6 & Eiajy6));
assign Uiajy6 = (!Txniw6);
assign E2cjy6 = (W5cjy6 ? Ccy7x6 : Jcy7x6);
assign W5cjy6 = (I8cjy6 & G5j7z6[17]);
assign I8cjy6 = (~(Q8cjy6 | S7cjy6));
assign S7cjy6 = (Nuniw6 & Czajy6);
assign Q8cjy6 = (Uly7x6 & A8cjy6);
assign A8cjy6 = (G5j7z6[16] & Y8cjy6);
assign Y8cjy6 = (~(Ao2jy6 & Czajy6));
assign Uly7x6 = (G9cjy6 & O9cjy6);
assign O9cjy6 = (~(Lgj7z6[50] & Mx38x6));
assign G9cjy6 = (W9cjy6 & Eacjy6);
assign Eacjy6 = (~(Macjy6 & Uacjy6));
assign Uacjy6 = (Cbcjy6 & Ccy7x6);
assign Macjy6 = (Lgj7z6[48] & Kbcjy6);
assign Kbcjy6 = (~(Lgj7z6[52] & Lky7x6));
assign Lky7x6 = (!Lgj7z6[49]);
assign W9cjy6 = (~(Sbcjy6 & Lgj7z6[49]));
assign Sbcjy6 = (Cbcjy6 & Sky7x6);
assign Sky7x6 = (!Lgj7z6[52]);
assign Cbcjy6 = (Mx38x6 | Lgj7z6[50]);
assign Mx38x6 = (!Lgj7z6[53]);
assign Ccy7x6 = (!Lgj7z6[51]);
assign Jcy7x6 = (!Lgj7z6[48]);
assign W1cjy6 = (M6cjy6 ? Ygy7x6 : Fhy7x6);
assign M6cjy6 = (Txniw6 & Accjy6);
assign Accjy6 = (Xjy7x6 | Eiajy6);
assign Eiajy6 = (~(G5j7z6[18] & Iccjy6));
assign Iccjy6 = (~(Jfmiw6 & Czajy6));
assign Xjy7x6 = (~(Qccjy6 & Yccjy6));
assign Yccjy6 = (~(Lgj7z6[56] & J648x6));
assign Qccjy6 = (Gdcjy6 & Odcjy6);
assign Odcjy6 = (~(Wdcjy6 & Eecjy6));
assign Eecjy6 = (Mecjy6 & Ygy7x6);
assign Wdcjy6 = (Lgj7z6[54] & Uecjy6);
assign Uecjy6 = (~(Lgj7z6[58] & Viy7x6));
assign Viy7x6 = (!Lgj7z6[55]);
assign Gdcjy6 = (~(Cfcjy6 & Lgj7z6[55]));
assign Cfcjy6 = (Mecjy6 & Oiy7x6);
assign Oiy7x6 = (!Lgj7z6[58]);
assign Mecjy6 = (J648x6 | Lgj7z6[56]);
assign J648x6 = (!Lgj7z6[59]);
assign Txniw6 = (G5j7z6[19] & Kfcjy6);
assign Kfcjy6 = (~(Czajy6 & Cn2jy6));
assign Ygy7x6 = (!Lgj7z6[57]);
assign Fhy7x6 = (!Lgj7z6[54]);
assign Cnajy6 = (Uybjy6 ? Agcjy6 : Sfcjy6);
assign Agcjy6 = (!Igcjy6);
assign Cvbjy6 = (Cjajy6 | Kjajy6);
assign Uubjy6 = (Qgcjy6 & Uybjy6);
assign Uybjy6 = (~(Ygcjy6 & Kjajy6));
assign Kjajy6 = (~(Ghcjy6 & Ohcjy6));
assign Ohcjy6 = (~(G5j7z6[23] & Ua5jy6));
assign Ghcjy6 = (Whcjy6 & Eicjy6);
assign Eicjy6 = (P43nv6 | Czajy6);
assign P43nv6 = (Z7oiw6 & Gomiw6);
assign Gomiw6 = (!G5j7z6[22]);
assign Z7oiw6 = (!G5j7z6[23]);
assign Whcjy6 = (~(G5j7z6[22] & Ac5jy6));
assign Ygcjy6 = (~(Micjy6 & Uicjy6));
assign Uicjy6 = (Cjcjy6 & Cjajy6);
assign Cjajy6 = (~(Kjcjy6 & Sjcjy6));
assign Sjcjy6 = (~(G5j7z6[21] & Wd5jy6));
assign Kjcjy6 = (Akcjy6 & Ikcjy6);
assign Ikcjy6 = (~(T63nv6 & Inj7x6));
assign Inj7x6 = (!Czajy6);
assign T63nv6 = (~(Y3oiw6 & Mkmiw6));
assign Mkmiw6 = (!G5j7z6[20]);
assign Y3oiw6 = (!G5j7z6[21]);
assign Akcjy6 = (~(G5j7z6[20] & Ue5jy6));
assign Cjcjy6 = (~(Qkcjy6 & Ykcjy6));
assign Ykcjy6 = (Gdajy6 ? May7x6 : Tay7x6);
assign May7x6 = (!Lgj7z6[66]);
assign Qkcjy6 = (Glcjy6 & Olcjy6);
assign Olcjy6 = (Sfcjy6 | Igcjy6);
assign Micjy6 = (Wlcjy6 & Emcjy6);
assign Emcjy6 = (~(Mmcjy6 & Igcjy6));
assign Igcjy6 = (Umcjy6 ? Lgj7z6[64] : Lgj7z6[61]);
assign Mmcjy6 = (Sfcjy6 & Glcjy6);
assign Glcjy6 = (Czbjy6 | Eybjy6);
assign Sfcjy6 = (Gdajy6 ? Oj48x6 : Cncjy6);
assign Wlcjy6 = (~(Eybjy6 & Czbjy6));
assign Czbjy6 = (Gdajy6 ? Ery7x6 : Xqy7x6);
assign Gdajy6 = (~(Kncjy6 & G5j7z6[23]));
assign Kncjy6 = (Sncjy6 & Aocjy6);
assign Aocjy6 = (~(Iocjy6 & Nsy7x6));
assign Nsy7x6 = (Qocjy6 & Yocjy6);
assign Yocjy6 = (~(Lgj7z6[68] & Xqy7x6));
assign Qocjy6 = (Gpcjy6 & Opcjy6);
assign Opcjy6 = (~(Wpcjy6 & Eqcjy6));
assign Eqcjy6 = (Mqcjy6 & Tay7x6);
assign Tay7x6 = (!Lgj7z6[69]);
assign Mqcjy6 = (~(Lgj7z6[70] & Oj48x6));
assign Oj48x6 = (!Lgj7z6[67]);
assign Wpcjy6 = (Lgj7z6[66] & Uqcjy6);
assign Gpcjy6 = (~(Crcjy6 & Lgj7z6[67]));
assign Crcjy6 = (Uqcjy6 & Cncjy6);
assign Cncjy6 = (!Lgj7z6[70]);
assign Uqcjy6 = (~(Lgj7z6[71] & Ery7x6));
assign Iocjy6 = (G5j7z6[22] & Krcjy6);
assign Krcjy6 = (~(Czajy6 & Rphov6));
assign Sncjy6 = (~(J6oiw6 & Czajy6));
assign Ery7x6 = (!Lgj7z6[68]);
assign Xqy7x6 = (!Lgj7z6[71]);
assign Eybjy6 = (Umcjy6 ? Lgj7z6[65] : Lgj7z6[62]);
assign Qgcjy6 = (Umcjy6 ? Lgj7z6[63] : Lgj7z6[60]);
assign Umcjy6 = (Srcjy6 & G5j7z6[21]);
assign Srcjy6 = (Ascjy6 & Iscjy6);
assign Iscjy6 = (~(Qscjy6 & Duy7x6));
assign Duy7x6 = (Yscjy6 & Gtcjy6);
assign Gtcjy6 = (~(Lgj7z6[62] & Lry7x6));
assign Lry7x6 = (!Lgj7z6[65]);
assign Yscjy6 = (Otcjy6 & Wtcjy6);
assign Wtcjy6 = (~(Eucjy6 & Mucjy6));
assign Mucjy6 = (~(Uucjy6 | Lgj7z6[63]));
assign Eucjy6 = (Lgj7z6[60] & Cvcjy6);
assign Cvcjy6 = (~(Lgj7z6[64] & Gw7iw6));
assign Gw7iw6 = (!Lgj7z6[61]);
assign Otcjy6 = (~(Kvcjy6 & Lgj7z6[61]));
assign Kvcjy6 = (~(Uucjy6 | Lgj7z6[64]));
assign Uucjy6 = (Lgj7z6[65] & Sh7iw6);
assign Sh7iw6 = (!Lgj7z6[62]);
assign Qscjy6 = (G5j7z6[20] & Svcjy6);
assign Svcjy6 = (~(Cshov6 & Czajy6));
assign Ascjy6 = (~(I2oiw6 & Czajy6));
assign Czajy6 = (Awcjy6 & Xxjov6);
assign I87jy6 = (Wp4jy6 ? Qwcjy6 : Iwcjy6);
assign Wp4jy6 = (~(Ywcjy6 & Gxcjy6));
assign Gxcjy6 = (~(Oxcjy6 & Wxcjy6));
assign Wxcjy6 = (~(Eycjy6 | Op4jy6));
assign Op4jy6 = (Mycjy6 & Gh2jy6);
assign Mycjy6 = (C74jy6 & Uycjy6);
assign C74jy6 = (Czcjy6 & Kzcjy6);
assign Kzcjy6 = (~(Szcjy6 | A0djy6));
assign Czcjy6 = (~(I0djy6 | Q0djy6));
assign Eycjy6 = (Od7jy6 & Y0djy6);
assign Y0djy6 = (~(G1djy6 & O1djy6));
assign O1djy6 = (Qwcjy6 | W1djy6);
assign Od7jy6 = (U2djy6 ? M2djy6 : E2djy6);
assign M2djy6 = (!C3djy6);
assign Oxcjy6 = (K3djy6 & S3djy6);
assign S3djy6 = (G1djy6 | Qwcjy6);
assign G1djy6 = (Gd7jy6 | W1djy6);
assign W1djy6 = (~(A4djy6 | Ag7jy6));
assign Gd7jy6 = (Y4djy6 ? Q4djy6 : I4djy6);
assign I4djy6 = (!G5djy6);
assign K3djy6 = (~(Ag7jy6 & A4djy6));
assign A4djy6 = (!Sf7jy6);
assign Sf7jy6 = (E6djy6 ? W5djy6 : O5djy6);
assign W5djy6 = (M6djy6 & U6djy6);
assign Ag7jy6 = (U2djy6 ? K7djy6 : C7djy6);
assign C7djy6 = (!S7djy6);
assign Ywcjy6 = (K74jy6 | M64jy6);
assign Qwcjy6 = (Y4djy6 ? I8djy6 : A8djy6);
assign Y4djy6 = (!E6djy6);
assign E6djy6 = (Q8djy6 & Y8djy6);
assign Y8djy6 = (~(G9djy6 & O9djy6));
assign O9djy6 = (O5djy6 | W9djy6);
assign G9djy6 = (Eadjy6 & Madjy6);
assign Madjy6 = (~(Uadjy6 & M6djy6));
assign M6djy6 = (Cbdjy6 | Kbdjy6);
assign Uadjy6 = (Sbdjy6 & U6djy6);
assign U6djy6 = (~(Gaj7z6[2] & Cbdjy6));
assign Sbdjy6 = (~(W9djy6 & O5djy6));
assign O5djy6 = (Qcdjy6 ? Icdjy6 : Acdjy6);
assign Acdjy6 = (~(Uycjy6 & Gx08x6));
assign W9djy6 = (~(Ycdjy6 | Gddjy6));
assign Gddjy6 = (~(G5djy6 | Q4djy6));
assign Ycdjy6 = (~(I8djy6 | Oddjy6));
assign Oddjy6 = (Q4djy6 & G5djy6);
assign G5djy6 = (Eedjy6 ? Wddjy6 : Gaj7z6[1]);
assign Q4djy6 = (Qcdjy6 ? Uedjy6 : Medjy6);
assign Uedjy6 = (!Cfdjy6);
assign Eadjy6 = (~(Kfdjy6 & Gh2jy6));
assign Kfdjy6 = (Uycjy6 & Sfdjy6);
assign Q8djy6 = (Q0djy6 | Szcjy6);
assign I8djy6 = (Qcdjy6 ? Igdjy6 : Agdjy6);
assign Qcdjy6 = (!Sfdjy6);
assign Sfdjy6 = (~(Qgdjy6 & Ygdjy6));
assign Ygdjy6 = (~(Ghdjy6 & Ohdjy6));
assign Ohdjy6 = (~(Uycjy6 & Whdjy6));
assign Whdjy6 = (~(Za2nv6 & Eidjy6));
assign Eidjy6 = (~(Midjy6 & Gx08x6));
assign Midjy6 = (~(Uidjy6 & Cjdjy6));
assign Cjdjy6 = (Cfdjy6 | Xg18x6);
assign Za2nv6 = (!Gh2jy6);
assign Gh2jy6 = (Kjdjy6 & Giliw6);
assign Kjdjy6 = (!Vs98x6);
assign Ghdjy6 = (~(Icdjy6 & Sjdjy6));
assign Sjdjy6 = (~(Akdjy6 & Uidjy6));
assign Uidjy6 = (~(Igdjy6 & Ikdjy6));
assign Ikdjy6 = (~(Cfdjy6 & Medjy6));
assign Medjy6 = (S74jy6 | Xg18x6);
assign S74jy6 = (!Uycjy6);
assign Akdjy6 = (~(Uycjy6 & Qkdjy6));
assign Qkdjy6 = (~(Ykdjy6 & Cfdjy6));
assign Cfdjy6 = (Oldjy6 ? Tcj7z6[1] : Gldjy6);
assign Ykdjy6 = (!Gx08x6);
assign Icdjy6 = (Oldjy6 ? Zw08x6 : Wldjy6);
assign Zw08x6 = (!Tcj7z6[2]);
assign Qgdjy6 = (I0djy6 | A0djy6);
assign Igdjy6 = (Oldjy6 ? F018x6 : Emdjy6);
assign Oldjy6 = (A0djy6 & Mmdjy6);
assign Mmdjy6 = (~(I0djy6 & Umdjy6));
assign Umdjy6 = (~(Cndjy6 & Kndjy6));
assign Kndjy6 = (~(Tcj7z6[2] & Wldjy6));
assign Cndjy6 = (~(Sndjy6 & Aodjy6));
assign Aodjy6 = (~(Gldjy6 & Ub18x6));
assign Sndjy6 = (Iodjy6 & Qodjy6);
assign Qodjy6 = (~(Yodjy6 & Gpdjy6));
assign Gpdjy6 = (Ub18x6 | Gldjy6);
assign Gldjy6 = (Opdjy6 ? Ffj7z6[1] : Zdj7z6[1]);
assign Ub18x6 = (!Tcj7z6[1]);
assign Iodjy6 = (Wldjy6 | Tcj7z6[2]);
assign Wldjy6 = (Opdjy6 ? Eqdjy6 : Wpdjy6);
assign I0djy6 = (~(Mqdjy6 & Uqdjy6));
assign Uqdjy6 = (~(Z3j7z6[1] & Wd5jy6));
assign Mqdjy6 = (Crdjy6 & Krdjy6);
assign Krdjy6 = (H73nv6 | H2m7x6);
assign H73nv6 = (R0m7x6 & Bvhov6);
assign Bvhov6 = (!Z3j7z6[0]);
assign R0m7x6 = (!Z3j7z6[1]);
assign Crdjy6 = (~(Z3j7z6[0] & Ue5jy6));
assign A0djy6 = (Z3j7z6[3] & Srdjy6);
assign Srdjy6 = (Ac5jy6 | Asdjy6);
assign F018x6 = (!Tcj7z6[0]);
assign Emdjy6 = (!Yodjy6);
assign Yodjy6 = (Opdjy6 ? Ffj7z6[0] : Zdj7z6[0]);
assign Opdjy6 = (~(Isdjy6 & Z3j7z6[1]));
assign Isdjy6 = (Qsdjy6 & Ysdjy6);
assign Ysdjy6 = (~(Gtdjy6 & Qg18x6));
assign Qg18x6 = (Otdjy6 & Wtdjy6);
assign Wtdjy6 = (~(Ffj7z6[2] & Wpdjy6));
assign Wpdjy6 = (!Zdj7z6[2]);
assign Otdjy6 = (Eudjy6 & Mudjy6);
assign Mudjy6 = (~(Uudjy6 & Cvdjy6));
assign Cvdjy6 = (~(Kvdjy6 | Zdj7z6[0]));
assign Kvdjy6 = (~(Svdjy6 | Ffj7z6[1]));
assign Uudjy6 = (Ffj7z6[0] & Awdjy6);
assign Eudjy6 = (~(Iwdjy6 & Ffj7z6[1]));
assign Iwdjy6 = (Awdjy6 & Svdjy6);
assign Svdjy6 = (!Zdj7z6[1]);
assign Awdjy6 = (~(Zdj7z6[2] & Eqdjy6));
assign Eqdjy6 = (!Ffj7z6[2]);
assign Gtdjy6 = (Z3j7z6[0] & Qwdjy6);
assign Qwdjy6 = (Ue5jy6 | Asdjy6);
assign Qsdjy6 = (Wd5jy6 | Asdjy6);
assign Agdjy6 = (~(Uycjy6 & M018x6));
assign Uycjy6 = (Ywdjy6 & Gxdjy6);
assign Gxdjy6 = (~(Fjadt6 & Uvgov6));
assign Uvgov6 = (Vs98x6 | Giliw6);
assign Vs98x6 = (~(Oxdjy6 & Me3jy6));
assign Oxdjy6 = (H2m7x6 & Flliw6);
assign Ywdjy6 = (~(X3get6 & N4fov6));
assign N4fov6 = (~(Cn2jy6 & H2m7x6));
assign A8djy6 = (!Wxdjy6);
assign Wxdjy6 = (Eedjy6 ? Eydjy6 : Gaj7z6[0]);
assign Eedjy6 = (!Cbdjy6);
assign Cbdjy6 = (~(Q0djy6 & Mydjy6));
assign Mydjy6 = (~(Uydjy6 & Szcjy6));
assign Szcjy6 = (Z3j7z6[7] & Czdjy6);
assign Czdjy6 = (Pfk7x6 | Asdjy6);
assign Uydjy6 = (Kzdjy6 & Szdjy6);
assign Szdjy6 = (~(Kbdjy6 & A0ejy6));
assign A0ejy6 = (~(I0ejy6 & Q0ejy6));
assign I0ejy6 = (Y0ejy6 & Cv08x6);
assign Cv08x6 = (!Gaj7z6[2]);
assign Kbdjy6 = (O1ejy6 ? G1ejy6 : Z318x6);
assign Z318x6 = (!Nbj7z6[2]);
assign Kzdjy6 = (~(Gaj7z6[2] & W1ejy6));
assign W1ejy6 = (~(Q0ejy6 & Y0ejy6));
assign Y0ejy6 = (Eydjy6 | E2ejy6);
assign E2ejy6 = (Wddjy6 & N418x6);
assign Q0ejy6 = (N418x6 | Wddjy6);
assign Wddjy6 = (O1ejy6 ? M2ejy6 : Nbj7z6[1]);
assign N418x6 = (!Gaj7z6[1]);
assign Q0djy6 = (~(U2ejy6 & C3ejy6));
assign C3ejy6 = (~(Z3j7z6[8] & K3ejy6));
assign Eydjy6 = (O1ejy6 ? S3ejy6 : Nbj7z6[0]);
assign O1ejy6 = (~(A4ejy6 | U2ejy6));
assign U2ejy6 = (~(I4ejy6 | Q4ejy6));
assign A4ejy6 = (Y4ejy6 & G5ejy6);
assign G5ejy6 = (O5ejy6 & W5ejy6);
assign W5ejy6 = (~(Nbj7z6[2] & G1ejy6));
assign O5ejy6 = (E6ejy6 & M6ejy6);
assign M6ejy6 = (U6ejy6 | S3ejy6);
assign U6ejy6 = (~(C7ejy6 & K7ejy6));
assign C7ejy6 = (S7ejy6 | Nbj7z6[1]);
assign E6ejy6 = (~(A8ejy6 & Nbj7z6[1]));
assign A8ejy6 = (S7ejy6 & K7ejy6);
assign K7ejy6 = (G1ejy6 | Nbj7z6[2]);
assign G1ejy6 = (I8ejy6 ? Q918x6 : X918x6);
assign S7ejy6 = (!M2ejy6);
assign M2ejy6 = (I8ejy6 ? Z8j7z6[1] : T7j7z6[1]);
assign Y4ejy6 = (Z3j7z6[8] & K3ejy6);
assign K3ejy6 = (Qpl7x6 | Asdjy6);
assign S3ejy6 = (I8ejy6 ? Z8j7z6[0] : T7j7z6[0]);
assign I8ejy6 = (~(Q4ejy6 & Q8ejy6));
assign Q8ejy6 = (~(Sa18x6 & I4ejy6));
assign I4ejy6 = (Z3j7z6[10] & Y8ejy6);
assign Y8ejy6 = (Erk7x6 | Asdjy6);
assign Sa18x6 = (G9ejy6 & O9ejy6);
assign O9ejy6 = (~(Z8j7z6[2] & X918x6));
assign X918x6 = (!T7j7z6[2]);
assign G9ejy6 = (W9ejy6 & Eaejy6);
assign Eaejy6 = (~(Maejy6 & Z8j7z6[1]));
assign Maejy6 = (Uaejy6 & Cbejy6);
assign W9ejy6 = (~(Kbejy6 & Sbejy6));
assign Sbejy6 = (~(Acejy6 | T7j7z6[0]));
assign Acejy6 = (~(Cbejy6 | Z8j7z6[1]));
assign Cbejy6 = (!T7j7z6[1]);
assign Kbejy6 = (Z8j7z6[0] & Uaejy6);
assign Uaejy6 = (~(T7j7z6[2] & Q918x6));
assign Q918x6 = (!Z8j7z6[2]);
assign Q4ejy6 = (Z3j7z6[11] & Icejy6);
assign Icejy6 = (Ue6jy6 | Asdjy6);
assign Asdjy6 = (!H2m7x6);
assign H2m7x6 = (Sz3jy6 & Xxjov6);
assign Iwcjy6 = (~(Qcejy6 & Ycejy6));
assign Ycejy6 = (~(Gdejy6 & Odejy6));
assign Odejy6 = (Meejy6 ? Eeejy6 : Wdejy6);
assign Eeejy6 = (Ueejy6 ? Bd08x6 : Zg8iw6);
assign Zg8iw6 = (!Lgj7z6[12]);
assign Gdejy6 = (~(Cfejy6 | U2djy6));
assign Qcejy6 = (U2djy6 ? Sfejy6 : Kfejy6);
assign U2djy6 = (Agejy6 & M64jy6);
assign M64jy6 = (~(Igejy6 & Qgejy6));
assign Qgejy6 = (Ygejy6 & Ghejy6);
assign Ygejy6 = (~(Dii7x6 | Emi7x6));
assign Igejy6 = (~(Ohejy6 | Whejy6));
assign Agejy6 = (~(Eiejy6 & Miejy6));
assign Miejy6 = (Uiejy6 & K74jy6);
assign K74jy6 = (~(Cjejy6 & Kjejy6));
assign Kjejy6 = (~(Sjejy6 | Akejy6));
assign Cjejy6 = (~(Ikejy6 | Qkejy6));
assign Uiejy6 = (E2djy6 | Ykejy6);
assign Ykejy6 = (Glejy6 & Olejy6);
assign Olejy6 = (Sfejy6 | Wlejy6);
assign E2djy6 = (Cfejy6 ? Mmejy6 : Emejy6);
assign Emejy6 = (Meejy6 ? Cnejy6 : Umejy6);
assign Eiejy6 = (Knejy6 & Snejy6);
assign Snejy6 = (Glejy6 | Sfejy6);
assign Glejy6 = (C3djy6 | Wlejy6);
assign Wlejy6 = (~(S7djy6 | K7djy6));
assign C3djy6 = (Qoejy6 ? Ioejy6 : Aoejy6);
assign Knejy6 = (~(K7djy6 & S7djy6));
assign S7djy6 = (Cfejy6 ? Gpejy6 : Yoejy6);
assign K7djy6 = (Qoejy6 ? Wpejy6 : Opejy6);
assign Sfejy6 = (Qoejy6 ? Mqejy6 : Eqejy6);
assign Qoejy6 = (Uqejy6 & Crejy6);
assign Crejy6 = (~(Krejy6 & Srejy6));
assign Srejy6 = (Ohejy6 | Asejy6);
assign Krejy6 = (Isejy6 & Qsejy6);
assign Qsejy6 = (~(Wpejy6 & Ysejy6));
assign Ysejy6 = (~(Opejy6 & Gtejy6));
assign Wpejy6 = (Euejy6 ? Wtejy6 : Otejy6);
assign Wtejy6 = (!Muejy6);
assign Isejy6 = (Gtejy6 | Opejy6);
assign Opejy6 = (Asejy6 ? Cvejy6 : Uuejy6);
assign Uuejy6 = (!Kvejy6);
assign Gtejy6 = (Svejy6 | Awejy6);
assign Awejy6 = (~(Aoejy6 | Eqejy6));
assign Svejy6 = (Ioejy6 & Iwejy6);
assign Iwejy6 = (~(Eqejy6 & Aoejy6));
assign Aoejy6 = (Asejy6 ? Ywejy6 : Qwejy6);
assign Ywejy6 = (!Gxejy6);
assign Ioejy6 = (Euejy6 ? Wxejy6 : Oxejy6);
assign Uqejy6 = (~(Eyejy6 & Ghejy6));
assign Eyejy6 = (!Whejy6);
assign Mqejy6 = (Euejy6 ? Uyejy6 : Myejy6);
assign Euejy6 = (Czejy6 | Ghejy6);
assign Ghejy6 = (Kzejy6 & Szejy6);
assign Szejy6 = (~(G5j7z6[15] & Ue6jy6));
assign Ue6jy6 = (!V6i7x6);
assign Kzejy6 = (A0fjy6 & I0fjy6);
assign I0fjy6 = (Xu2nv6 | Q0fjy6);
assign Xu2nv6 = (M4j7x6 & Qzi7x6);
assign Qzi7x6 = (!G5j7z6[14]);
assign M4j7x6 = (!G5j7z6[15]);
assign A0fjy6 = (~(G5j7z6[14] & Erk7x6));
assign Erk7x6 = (!P3i7x6);
assign Czejy6 = (Y0fjy6 & G1fjy6);
assign G1fjy6 = (O1fjy6 & Whejy6);
assign Whejy6 = (~(W1fjy6 & E2fjy6));
assign E2fjy6 = (~(G5j7z6[13] & Ktl7x6));
assign Ktl7x6 = (!Jrj7x6);
assign W1fjy6 = (M2fjy6 & U2fjy6);
assign U2fjy6 = (~(Dy2nv6 & B2j7x6));
assign Dy2nv6 = (~(Dwi7x6 & Csi7x6));
assign Csi7x6 = (!G5j7z6[12]);
assign Dwi7x6 = (!G5j7z6[13]);
assign M2fjy6 = (~(G5j7z6[12] & Qpl7x6));
assign O1fjy6 = (~(C3fjy6 & K3fjy6));
assign K3fjy6 = (S3fjy6 ? Ki38x6 : Gn38x6);
assign Ki38x6 = (!Lgj7z6[42]);
assign C3fjy6 = (A4fjy6 & I4fjy6);
assign I4fjy6 = (Q4fjy6 | Wxejy6);
assign Y0fjy6 = (Y4fjy6 & G5fjy6);
assign G5fjy6 = (~(O5fjy6 & Wxejy6));
assign Wxejy6 = (W5fjy6 ? Lgj7z6[40] : Lgj7z6[37]);
assign O5fjy6 = (Q4fjy6 & A4fjy6);
assign A4fjy6 = (Otejy6 | Muejy6);
assign Q4fjy6 = (!Oxejy6);
assign Oxejy6 = (S3fjy6 ? Lgj7z6[43] : Lgj7z6[46]);
assign Y4fjy6 = (~(Muejy6 & Otejy6));
assign Otejy6 = (S3fjy6 ? Ak38x6 : Po38x6);
assign Muejy6 = (W5fjy6 ? Lgj7z6[41] : Lgj7z6[38]);
assign Uyejy6 = (W5fjy6 ? Lgj7z6[39] : Lgj7z6[36]);
assign W5fjy6 = (E6fjy6 & G5j7z6[13]);
assign E6fjy6 = (M6fjy6 & U6fjy6);
assign U6fjy6 = (~(C7fjy6 & Psz7x6));
assign Psz7x6 = (K7fjy6 & S7fjy6);
assign S7fjy6 = (~(Lgj7z6[38] & Qe38x6));
assign K7fjy6 = (A8fjy6 & I8fjy6);
assign I8fjy6 = (~(Q8fjy6 & Y8fjy6));
assign Y8fjy6 = (G9fjy6 & Hd38x6);
assign Hd38x6 = (!Lgj7z6[39]);
assign Q8fjy6 = (Lgj7z6[36] & O9fjy6);
assign O9fjy6 = (~(Lgj7z6[40] & N938x6));
assign N938x6 = (!Lgj7z6[37]);
assign A8fjy6 = (~(W9fjy6 & Lgj7z6[37]));
assign W9fjy6 = (G9fjy6 & Ef38x6);
assign Ef38x6 = (!Lgj7z6[40]);
assign G9fjy6 = (Qe38x6 | Lgj7z6[38]);
assign Qe38x6 = (!Lgj7z6[41]);
assign C7fjy6 = (G5j7z6[12] & Eafjy6);
assign Eafjy6 = (~(Q0fjy6 & L1i7x6));
assign M6fjy6 = (~(Jrj7x6 & Q0fjy6));
assign Myejy6 = (S3fjy6 ? Lgj7z6[42] : Lgj7z6[45]);
assign S3fjy6 = (~(Mafjy6 & G5j7z6[15]));
assign Mafjy6 = (Uafjy6 & Cbfjy6);
assign Cbfjy6 = (~(Kbfjy6 & Grz7x6));
assign Grz7x6 = (Sbfjy6 & Acfjy6);
assign Acfjy6 = (~(Icfjy6 & Lgj7z6[43]));
assign Icfjy6 = (Qcfjy6 & Qpz7x6);
assign Qpz7x6 = (!Lgj7z6[46]);
assign Sbfjy6 = (Ycfjy6 & Gdfjy6);
assign Gdfjy6 = (~(Odfjy6 & Wdfjy6));
assign Wdfjy6 = (Eefjy6 & Gn38x6);
assign Gn38x6 = (!Lgj7z6[45]);
assign Eefjy6 = (~(Lgj7z6[46] & Xpz7x6));
assign Xpz7x6 = (!Lgj7z6[43]);
assign Odfjy6 = (Lgj7z6[42] & Qcfjy6);
assign Qcfjy6 = (~(Lgj7z6[47] & Ak38x6));
assign Ak38x6 = (!Lgj7z6[44]);
assign Ycfjy6 = (~(Lgj7z6[44] & Po38x6));
assign Po38x6 = (!Lgj7z6[47]);
assign Kbfjy6 = (G5j7z6[14] & Mefjy6);
assign Mefjy6 = (~(Q0fjy6 & P3i7x6));
assign Uafjy6 = (~(Q0fjy6 & V6i7x6));
assign Eqejy6 = (!Uefjy6);
assign Uefjy6 = (Asejy6 ? Kffjy6 : Cffjy6);
assign Asejy6 = (Sffjy6 & Agfjy6);
assign Agfjy6 = (~(Igfjy6 & Qgfjy6));
assign Qgfjy6 = (Ygfjy6 & Ohejy6);
assign Ohejy6 = (~(Ghfjy6 & U9i7x6));
assign Ghfjy6 = (~(G5j7z6[9] & Ohfjy6));
assign Ygfjy6 = (~(Whfjy6 & Kffjy6));
assign Whfjy6 = (Eifjy6 & Mifjy6);
assign Eifjy6 = (Gxejy6 | Qwejy6);
assign Igfjy6 = (Uifjy6 & Cjfjy6);
assign Cjfjy6 = (~(Kjfjy6 & Qwejy6));
assign Qwejy6 = (Sjfjy6 ? Lgj7z6[28] : Lgj7z6[25]);
assign Kjfjy6 = (Gxejy6 & Mifjy6);
assign Mifjy6 = (Cvejy6 | Kvejy6);
assign Gxejy6 = (Akfjy6 ? Wzz7x6 : Pzz7x6);
assign Uifjy6 = (~(Kvejy6 & Cvejy6));
assign Cvejy6 = (Akfjy6 ? Q038x6 : Y438x6);
assign Kvejy6 = (Sjfjy6 ? Lgj7z6[29] : Lgj7z6[26]);
assign Sffjy6 = (Emi7x6 | Dii7x6);
assign Kffjy6 = (Akfjy6 ? Lxz7x6 : Exz7x6);
assign Akfjy6 = (~(Emi7x6 & Ikfjy6));
assign Ikfjy6 = (~(Dii7x6 & Y008x6));
assign Y008x6 = (Qkfjy6 & Ykfjy6);
assign Ykfjy6 = (~(Lgj7z6[32] & Y438x6));
assign Y438x6 = (!Lgj7z6[35]);
assign Qkfjy6 = (Glfjy6 & Olfjy6);
assign Olfjy6 = (~(Wlfjy6 & Emfjy6));
assign Emfjy6 = (Mmfjy6 & Exz7x6);
assign Mmfjy6 = (~(Lgj7z6[34] & Wzz7x6));
assign Wzz7x6 = (!Lgj7z6[31]);
assign Wlfjy6 = (Lgj7z6[30] & Umfjy6);
assign Glfjy6 = (~(Cnfjy6 & Lgj7z6[31]));
assign Cnfjy6 = (Umfjy6 & Pzz7x6);
assign Pzz7x6 = (!Lgj7z6[34]);
assign Umfjy6 = (~(Lgj7z6[35] & Q038x6));
assign Q038x6 = (!Lgj7z6[32]);
assign Dii7x6 = (G5j7z6[10] & Knfjy6);
assign Knfjy6 = (~(Q0fjy6 & Nfj7x6));
assign Emi7x6 = (G5j7z6[11] & Snfjy6);
assign Snfjy6 = (~(Q0fjy6 & Hzh7x6));
assign Lxz7x6 = (!Lgj7z6[30]);
assign Exz7x6 = (!Lgj7z6[33]);
assign Cffjy6 = (Sjfjy6 ? Gkz7x6 : Eg8iw6);
assign Sjfjy6 = (Aofjy6 & G5j7z6[9]);
assign Aofjy6 = (Iofjy6 & Ohfjy6);
assign Ohfjy6 = (B2j7x6 | U7k7x6);
assign Iofjy6 = (U9i7x6 | Bzz7x6);
assign Bzz7x6 = (~(Qofjy6 & Yofjy6));
assign Yofjy6 = (~(Lgj7z6[26] & Uv28x6));
assign Uv28x6 = (!Lgj7z6[29]);
assign Qofjy6 = (Gpfjy6 & Opfjy6);
assign Opfjy6 = (~(Wpfjy6 & Eqfjy6));
assign Eqfjy6 = (Mqfjy6 & Gkz7x6);
assign Mqfjy6 = (~(Lgj7z6[28] & Dy7iw6));
assign Dy7iw6 = (!Lgj7z6[25]);
assign Wpfjy6 = (Lgj7z6[24] & Uqfjy6);
assign Gpfjy6 = (~(Crfjy6 & Lgj7z6[25]));
assign Crfjy6 = (Uqfjy6 & Zxz7x6);
assign Zxz7x6 = (!Lgj7z6[28]);
assign Uqfjy6 = (~(Lgj7z6[29] & Kk7iw6));
assign Kk7iw6 = (!Lgj7z6[26]);
assign U9i7x6 = (~(G5j7z6[8] & Krfjy6));
assign Krfjy6 = (~(Q0fjy6 & Uy2jy6));
assign Gkz7x6 = (!Lgj7z6[27]);
assign Eg8iw6 = (!Lgj7z6[24]);
assign Kfejy6 = (~(Srfjy6 & Cfejy6));
assign Cfejy6 = (~(Asfjy6 & Isfjy6));
assign Isfjy6 = (~(Qsfjy6 & Ysfjy6));
assign Ysfjy6 = (Qkejy6 | Gtfjy6);
assign Qsfjy6 = (Otfjy6 & Wtfjy6);
assign Wtfjy6 = (~(Eufjy6 & Mufjy6));
assign Mufjy6 = (Gpejy6 | Uufjy6);
assign Eufjy6 = (Cvfjy6 & Kvfjy6);
assign Kvfjy6 = (~(Svfjy6 & Awfjy6));
assign Awfjy6 = (Srfjy6 | Mmejy6);
assign Svfjy6 = (Meejy6 ? Qwfjy6 : Iwfjy6);
assign Cvfjy6 = (~(Mmejy6 & Srfjy6));
assign Mmejy6 = (Gtfjy6 ? Gxfjy6 : Ywfjy6);
assign Otfjy6 = (~(Uufjy6 & Gpejy6));
assign Gpejy6 = (Gtfjy6 ? Wxfjy6 : Oxfjy6);
assign Wxfjy6 = (!Eyfjy6);
assign Uufjy6 = (!Yoejy6);
assign Yoejy6 = (Meejy6 ? Uyfjy6 : Myfjy6);
assign Meejy6 = (~(Czfjy6 & Akejy6));
assign Czfjy6 = (~(Kzfjy6 & Szfjy6));
assign Szfjy6 = (A0gjy6 & Sjejy6);
assign A0gjy6 = (~(I0gjy6 & Wdejy6));
assign Wdejy6 = (Q0gjy6 ? Ol28x6 : Sg28x6);
assign Sg28x6 = (!Lgj7z6[18]);
assign I0gjy6 = (Y0gjy6 & G1gjy6);
assign G1gjy6 = (~(Iwfjy6 & Cnejy6));
assign Cnejy6 = (!Qwfjy6);
assign Iwfjy6 = (!Umejy6);
assign Kzfjy6 = (O1gjy6 & W1gjy6);
assign W1gjy6 = (~(E2gjy6 & Qwfjy6));
assign Qwfjy6 = (Ueejy6 ? Lgj7z6[16] : Lgj7z6[13]);
assign E2gjy6 = (Umejy6 & Y0gjy6);
assign Y0gjy6 = (~(Myfjy6 & M2gjy6));
assign Umejy6 = (Q0gjy6 ? En28x6 : Bi28x6);
assign O1gjy6 = (M2gjy6 | Myfjy6);
assign M2gjy6 = (!Uyfjy6);
assign Uyfjy6 = (Ueejy6 ? Lgj7z6[17] : Lgj7z6[14]);
assign Ueejy6 = (U2gjy6 & G5j7z6[5]);
assign U2gjy6 = (C3gjy6 & K3gjy6);
assign K3gjy6 = (~(S3gjy6 & Qh08x6));
assign Qh08x6 = (A4gjy6 & I4gjy6);
assign I4gjy6 = (~(Lgj7z6[14] & Ff08x6));
assign A4gjy6 = (Q4gjy6 & Y4gjy6);
assign Y4gjy6 = (~(G5gjy6 & O5gjy6));
assign O5gjy6 = (W5gjy6 & Bd08x6);
assign Bd08x6 = (!Lgj7z6[15]);
assign G5gjy6 = (Lgj7z6[12] & E6gjy6);
assign E6gjy6 = (~(Lgj7z6[16] & Yy7iw6));
assign Yy7iw6 = (!Lgj7z6[13]);
assign Q4gjy6 = (~(M6gjy6 & Lgj7z6[13]));
assign M6gjy6 = (W5gjy6 & Md28x6);
assign Md28x6 = (!Lgj7z6[16]);
assign W5gjy6 = (Ff08x6 | Lgj7z6[14]);
assign Ff08x6 = (!Lgj7z6[17]);
assign S3gjy6 = (G5j7z6[4] & U6gjy6);
assign U6gjy6 = (~(Cshov6 & Q0fjy6));
assign C3gjy6 = (~(I2oiw6 & Q0fjy6));
assign Myfjy6 = (Q0gjy6 ? Lgj7z6[23] : Lgj7z6[20]);
assign Q0gjy6 = (C7gjy6 & G5j7z6[7]);
assign C7gjy6 = (K7gjy6 & S7gjy6);
assign S7gjy6 = (~(A8gjy6 & Hg08x6));
assign Hg08x6 = (I8gjy6 & Q8gjy6);
assign Q8gjy6 = (~(Lgj7z6[20] & Ke08x6));
assign I8gjy6 = (Y8gjy6 & G9gjy6);
assign G9gjy6 = (~(O9gjy6 & W9gjy6));
assign W9gjy6 = (Eagjy6 & Ol28x6);
assign Ol28x6 = (!Lgj7z6[21]);
assign O9gjy6 = (Lgj7z6[18] & Magjy6);
assign Magjy6 = (~(Lgj7z6[22] & Bi28x6));
assign Bi28x6 = (!Lgj7z6[19]);
assign Y8gjy6 = (~(Uagjy6 & Lgj7z6[19]));
assign Uagjy6 = (Eagjy6 & En28x6);
assign En28x6 = (!Lgj7z6[22]);
assign Eagjy6 = (Ke08x6 | Lgj7z6[20]);
assign Ke08x6 = (!Lgj7z6[23]);
assign A8gjy6 = (G5j7z6[6] & Cbgjy6);
assign Cbgjy6 = (~(Q0fjy6 & Rphov6));
assign K7gjy6 = (~(J6oiw6 & Q0fjy6));
assign Asfjy6 = (Sjejy6 | Akejy6);
assign Akejy6 = (~(Kbgjy6 & Sbgjy6));
assign Sbgjy6 = (~(G5j7z6[7] & Ua5jy6));
assign Ua5jy6 = (!J6oiw6);
assign Kbgjy6 = (Acgjy6 & Icgjy6);
assign Icgjy6 = (~(M63nv6 & B2j7x6));
assign B2j7x6 = (!Q0fjy6);
assign M63nv6 = (~(Vrniw6 & V7miw6));
assign V7miw6 = (!G5j7z6[6]);
assign Vrniw6 = (!G5j7z6[7]);
assign Acgjy6 = (~(G5j7z6[6] & Ac5jy6));
assign Ac5jy6 = (!Rphov6);
assign Sjejy6 = (~(Qcgjy6 & Ycgjy6));
assign Ycgjy6 = (~(G5j7z6[5] & Wd5jy6));
assign Wd5jy6 = (!I2oiw6);
assign Qcgjy6 = (Gdgjy6 & Odgjy6);
assign Odgjy6 = (F63nv6 | Q0fjy6);
assign F63nv6 = (Nnniw6 & B4miw6);
assign B4miw6 = (!G5j7z6[4]);
assign Nnniw6 = (!G5j7z6[5]);
assign Gdgjy6 = (~(G5j7z6[4] & Ue5jy6));
assign Srfjy6 = (Gtfjy6 ? Eegjy6 : Wdgjy6);
assign Gtfjy6 = (Megjy6 & Ikejy6);
assign Ikejy6 = (~(Uegjy6 & Cfgjy6));
assign Cfgjy6 = (~(G5j7z6[3] & Xdoiw6));
assign Uegjy6 = (Kfgjy6 & Sfgjy6);
assign Sfgjy6 = (O73nv6 | Q0fjy6);
assign O73nv6 = (~(G5j7z6[3] | G5j7z6[2]));
assign Kfgjy6 = (~(G5j7z6[2] & Zumiw6));
assign Megjy6 = (~(Aggjy6 & Iggjy6));
assign Iggjy6 = (Qggjy6 & Qkejy6);
assign Qkejy6 = (~(Yggjy6 & Ghgjy6));
assign Ghgjy6 = (~(G5j7z6[1] & Daoiw6));
assign Yggjy6 = (Ohgjy6 & Whgjy6);
assign Whgjy6 = (V73nv6 | Q0fjy6);
assign V73nv6 = (~(G5j7z6[1] | G5j7z6[0]));
assign Ohgjy6 = (~(G5j7z6[0] & Rqmiw6));
assign Qggjy6 = (~(Eigjy6 & Eegjy6));
assign Eigjy6 = (Migjy6 & Uigjy6);
assign Uigjy6 = (Gxfjy6 | Cjgjy6);
assign Aggjy6 = (Kjgjy6 & Sjgjy6);
assign Sjgjy6 = (~(Akgjy6 & Cjgjy6));
assign Cjgjy6 = (!Ywfjy6);
assign Ywfjy6 = (Ikgjy6 ? Co08x6 : Vn08x6);
assign Akgjy6 = (Gxfjy6 & Migjy6);
assign Migjy6 = (Eyfjy6 | Oxfjy6);
assign Gxfjy6 = (Qkgjy6 ? Zp08x6 : Sp08x6);
assign Qkgjy6 = (!Ykgjy6);
assign Kjgjy6 = (~(Oxfjy6 & Eyfjy6));
assign Eyfjy6 = (Ykgjy6 ? I428x6 : A028x6);
assign Oxfjy6 = (Ikgjy6 ? Lgj7z6[5] : Lgj7z6[2]);
assign Eegjy6 = (Ykgjy6 ? Fm08x6 : Mm08x6);
assign Ykgjy6 = (Glgjy6 & G5j7z6[3]);
assign Glgjy6 = (Olgjy6 & Wlgjy6);
assign Wlgjy6 = (~(Emgjy6 & Br08x6));
assign Br08x6 = (Mmgjy6 & Umgjy6);
assign Umgjy6 = (~(Lgj7z6[8] & I428x6));
assign I428x6 = (!Lgj7z6[11]);
assign Mmgjy6 = (Cngjy6 & Kngjy6);
assign Kngjy6 = (~(Sngjy6 & Aogjy6));
assign Aogjy6 = (Iogjy6 & Fm08x6);
assign Iogjy6 = (~(Lgj7z6[10] & Zp08x6));
assign Zp08x6 = (!Lgj7z6[7]);
assign Sngjy6 = (Lgj7z6[6] & Qogjy6);
assign Cngjy6 = (~(Yogjy6 & Lgj7z6[7]));
assign Yogjy6 = (Qogjy6 & Sp08x6);
assign Sp08x6 = (!Lgj7z6[10]);
assign Qogjy6 = (~(Lgj7z6[11] & A028x6));
assign A028x6 = (!Lgj7z6[8]);
assign Emgjy6 = (G5j7z6[2] & Gpgjy6);
assign Gpgjy6 = (~(Q0fjy6 & Jfmiw6));
assign Olgjy6 = (~(Q0fjy6 & Cn2jy6));
assign Fm08x6 = (!Lgj7z6[9]);
assign Mm08x6 = (!Lgj7z6[6]);
assign Wdgjy6 = (Ikgjy6 ? T808x6 : M808x6);
assign Ikgjy6 = (Opgjy6 & G5j7z6[1]);
assign Opgjy6 = (Wpgjy6 & Eqgjy6);
assign Eqgjy6 = (~(Mqgjy6 & Ep08x6));
assign Ep08x6 = (Uqgjy6 & Crgjy6);
assign Crgjy6 = (~(Lgj7z6[2] & On08x6));
assign Uqgjy6 = (Krgjy6 & Srgjy6);
assign Srgjy6 = (~(Asgjy6 & Isgjy6));
assign Isgjy6 = (Qsgjy6 & T808x6);
assign Asgjy6 = (Lgj7z6[0] & Ysgjy6);
assign Ysgjy6 = (~(Lgj7z6[4] & Vn08x6));
assign Vn08x6 = (!Lgj7z6[1]);
assign Krgjy6 = (~(Gtgjy6 & Lgj7z6[1]));
assign Gtgjy6 = (Qsgjy6 & Co08x6);
assign Co08x6 = (!Lgj7z6[4]);
assign Qsgjy6 = (On08x6 | Lgj7z6[2]);
assign On08x6 = (!Lgj7z6[5]);
assign Mqgjy6 = (G5j7z6[0] & Otgjy6);
assign Otgjy6 = (~(Q0fjy6 & Ao2jy6));
assign Wpgjy6 = (~(Q0fjy6 & Nuniw6));
assign Q0fjy6 = (Wtgjy6 & Xxjov6);
assign Xxjov6 = (!Nob7z6[8]);
assign T808x6 = (!Lgj7z6[3]);
assign M808x6 = (!Lgj7z6[0]);
assign A44jy6 = (Eugjy6 & Mugjy6);
assign Mugjy6 = (~(Uugjy6 & Cvgjy6));
assign Cvgjy6 = (~(Q04jy6 & Kvgjy6));
assign Q04jy6 = (!Y84jy6);
assign Uugjy6 = (Svgjy6 & J92nv6);
assign Svgjy6 = (~(Awgjy6 & H1m8v6));
assign Awgjy6 = (Ppb7z6[7] & Iwgjy6);
assign Iwgjy6 = (~(Qwgjy6 & Y84jy6));
assign Y84jy6 = (~(Ywgjy6 & Gxgjy6));
assign Gxgjy6 = (~(H1m8v6 & Oxgjy6));
assign Oxgjy6 = (~(Wxgjy6 & Eygjy6));
assign Eygjy6 = (Mygjy6 & Uygjy6);
assign Uygjy6 = (~(Q0oiy6 & Gaj7z6[2]));
assign Mygjy6 = (~(Tcj7z6[2] & Cvniy6));
assign Wxgjy6 = (Czgjy6 & Kzgjy6);
assign Kzgjy6 = (~(Ffj7z6[2] & Szgjy6));
assign Czgjy6 = (~(Zdj7z6[2] & Gd2jy6));
assign Ywgjy6 = (~(Lh18x6 & Pahov6));
assign Pahov6 = (H1m8v6 & Nbj7z6[2]);
assign Qwgjy6 = (!Kvgjy6);
assign Kvgjy6 = (~(A0hjy6 & I0hjy6));
assign I0hjy6 = (~(Q0hjy6 & E24jy6));
assign E24jy6 = (!K34jy6);
assign Q0hjy6 = (Zyl8v6 & Ppb7z6[6]);
assign A0hjy6 = (~(Y0hjy6 & U24jy6));
assign U24jy6 = (Gpu5z6 & Opu5z6);
assign Opu5z6 = (Wpu5z6 & Equ5z6);
assign Equ5z6 = (~(Tcj7z6[0] & Cvniy6));
assign Wpu5z6 = (Mqu5z6 & Uqu5z6);
assign Uqu5z6 = (~(Lh18x6 & Nbj7z6[0]));
assign Mqu5z6 = (~(Q0oiy6 & Gaj7z6[0]));
assign Gpu5z6 = (Cru5z6 & Rwl8v6);
assign Cru5z6 = (Kru5z6 & Sru5z6);
assign Sru5z6 = (~(Ffj7z6[0] & Szgjy6));
assign Kru5z6 = (~(Zdj7z6[0] & Gd2jy6));
assign Y0hjy6 = (Ppb7z6[5] & Asu5z6);
assign Asu5z6 = (~(K34jy6 & I8oiy6));
assign K34jy6 = (~(Isu5z6 & Qsu5z6));
assign Qsu5z6 = (~(Zyl8v6 & Ysu5z6));
assign Ysu5z6 = (~(Gtu5z6 & Otu5z6));
assign Otu5z6 = (Wtu5z6 & Euu5z6);
assign Euu5z6 = (~(Q0oiy6 & Gaj7z6[1]));
assign Q0oiy6 = (!Q8ziy6);
assign Wtu5z6 = (~(Tcj7z6[1] & Cvniy6));
assign Gtu5z6 = (Muu5z6 & Uuu5z6);
assign Uuu5z6 = (~(Ffj7z6[1] & Szgjy6));
assign Muu5z6 = (~(Zdj7z6[1] & Gd2jy6));
assign Isu5z6 = (~(Lh18x6 & Jehov6));
assign Jehov6 = (Zyl8v6 & Nbj7z6[1]);
assign Eugjy6 = (~(Cvu5z6 & Kvu5z6));
assign Kvu5z6 = (Svu5z6 & Awu5z6);
assign Awu5z6 = (~(Micet6 & Cvniy6));
assign Cvniy6 = (~(Iwu5z6 & Glviy6));
assign Glviy6 = (T5b7x6 & Qwu5z6);
assign Qwu5z6 = (~(Zjb7z6[8] | Zjb7z6[9]));
assign T5b7x6 = (~(Qg77z6 | Ig77z6));
assign Iwu5z6 = (Ywu5z6 & Wlviy6);
assign Wlviy6 = (W3b7x6 & O6b7x6);
assign O6b7x6 = (~(Pxfov6 & Gxu5z6));
assign Gxu5z6 = (~(Oxu5z6 & Mah7v6));
assign Oxu5z6 = (~(F4edt6 & Xsinv6));
assign W3b7x6 = (~(B6edt6 & Pxfov6));
assign Ywu5z6 = (Qc77z6 & Wwgov6);
assign Wwgov6 = (E697z6 & Wxu5z6);
assign Wxu5z6 = (Ftlov6 | Tlmov6);
assign Svu5z6 = (Eyu5z6 & Q8ziy6);
assign Q8ziy6 = (~(Myu5z6 & F4edt6));
assign Myu5z6 = (Etinv6 & Pxfov6);
assign Eyu5z6 = (~(Lh18x6 & E1cet6));
assign Lh18x6 = (Ffadt6 & Amg7x6);
assign Amg7x6 = (~(A0fet6 & Uyu5z6));
assign Uyu5z6 = (Nneet6 | Cwadt6);
assign Cvu5z6 = (Czu5z6 & Kzu5z6);
assign Kzu5z6 = (~(Ykcet6 & Szgjy6));
assign Szgjy6 = (!W9ziy6);
assign W9ziy6 = (Szu5z6 & Uva7x6);
assign Uva7x6 = (~(Wkb7z6[0] | Wkb7z6[2]));
assign Szu5z6 = (Gd77z6 & M697z6);
assign Czu5z6 = (~(Sjcet6 & Gd2jy6));
assign Gd2jy6 = (~(Emviy6 & A0v5z6));
assign A0v5z6 = (~(I0v5z6 & Mlmov6));
assign I0v5z6 = (~(Wwa7x6 & Losiw6));
assign Losiw6 = (!Tlb7z6[4]);
assign Wwa7x6 = (~(Tlb7z6[3] | Tlb7z6[0]));
assign Emviy6 = (~(Tlb7z6[1] & Mlmov6));
assign Mlmov6 = (~(Fuadt6 & Xsinv6));
assign Xsinv6 = (!Etinv6);
assign Qc2jy6 = (Jws7x6 | S8b7x6);
assign S8b7x6 = (Q0v5z6 & Ifo7v6);
assign Q0v5z6 = (~(Y0v5z6 & Sb0jy6));
assign Y0v5z6 = (Ac0jy6 & O1eiw6);
assign O1eiw6 = (G1v5z6 | O1v5z6);
assign O1v5z6 = (Qln7z6[1] ? E2v5z6 : W1v5z6);
assign E2v5z6 = (HREADYS & Y0kiw6);
assign Y0kiw6 = (~(M2v5z6 & U2v5z6));
assign M2v5z6 = (Gazet6 & C3v5z6);
assign C3v5z6 = (Kyn7z6[0] | Kyn7z6[1]);
assign W1v5z6 = (Uvixx6 ? K3v5z6 : HREADYD);
assign Uvixx6 = (~(Xnnyx6 & Hm1ov6));
assign Xnnyx6 = (B2jnv6 & Zgonv6);
assign Zgonv6 = (!Zblov6);
assign K3v5z6 = (S3v5z6 & HREADYS);
assign G1v5z6 = (~(A4v5z6 & Ag0jy6));
assign Ac0jy6 = (~(I4v5z6 & Q4v5z6));
assign Q4v5z6 = (~(HRESPD[0] & Qln7z6[0]));
assign I4v5z6 = (~(HRESPS[0] & Qln7z6[1]));
assign Jws7x6 = (!Sjcet6);
assign Ohi7v6 = (Euziy6 ? U47iw6 : H1j7z6[8]);
assign Euziy6 = (Y4v5z6 & Y82jy6);
assign Y4v5z6 = (R58iw6 & Bqi7z6[1]);
assign Hhi7v6 = (Hr4yx6 ? U47iw6 : H56ft6);
assign Ahi7v6 = (Sv1jy6 ? U47iw6 : Ies7z6[8]);
assign Sv1jy6 = (G5v5z6 & Cv1jy6);
assign G5v5z6 = (Ihs7z6[1] & O5v5z6);
assign O5v5z6 = (~(C397z6 & Scs7z6[1]));
assign Tgi7v6 = (O91jy6 ? U47iw6 : T077v6);
assign Mgi7v6 = (Ua1jy6 ? U47iw6 : Sgymz6[5]);
assign Fgi7v6 = (U61jy6 ? U47iw6 : Ojymz6[5]);
assign Yfi7v6 = (G91jy6 ? U47iw6 : Biymz6[8]);
assign G91jy6 = (Xid8x6 & Ddpyx6);
assign Ddpyx6 = (W5v5z6 & E6v5z6);
assign E6v5z6 = (M6v5z6 & Xfymz6[6]);
assign M6v5z6 = (Xfymz6[8] & R6pyx6);
assign W5v5z6 = (D9pyx6 & U6v5z6);
assign Rfi7v6 = (M61jy6 ? U47iw6 : Unymz6[5]);
assign Kfi7v6 = (W10jy6 ? Ykcet6 : Is5iw6);
assign W10jy6 = (~(Bzl7x6 & Bqi7z6[2]));
assign Bzl7x6 = (C7v5z6 & Eec7x6);
assign Eec7x6 = (~(K7v5z6 | S7v5z6));
assign K7v5z6 = (!G42nv6);
assign G42nv6 = (A8v5z6 & Qkfiy6);
assign A8v5z6 = (Toi7z6[8] & Qgfiy6);
assign C7v5z6 = (Wdm7x6 & Toi7z6[2]);
assign Wdm7x6 = (~(Toi7z6[3] | Toi7z6[4]));
assign Dfi7v6 = (Hyhov6 ? Is5iw6 : E1cet6);
assign Hyhov6 = (~(Uq0jy6 | Ie5iw6));
assign Ie5iw6 = (!Bqi7z6[2]);
assign Uq0jy6 = (!E60jy6);
assign E60jy6 = (I8v5z6 & Toi7z6[3]);
assign I8v5z6 = (~(Pb8iw6 | N92iw6));
assign N92iw6 = (~(Q8v5z6 & Y8v5z6));
assign Y8v5z6 = (~(Ualhy6 | S7v5z6));
assign S7v5z6 = (!S98iw6);
assign S98iw6 = (~(E32nv6 | Toi7z6[9]));
assign E32nv6 = (!Toi7z6[5]);
assign Ualhy6 = (~(G9v5z6 & Toi7z6[7]));
assign G9v5z6 = (Toi7z6[6] & Qgfiy6);
assign Qgfiy6 = (Toi7z6[11] & Toi7z6[10]);
assign Q8v5z6 = (Toi7z6[8] & Toi7z6[4]);
assign Wei7v6 = (Wtziy6 ? Is5iw6 : H1j7z6[16]);
assign Wtziy6 = (O9v5z6 & Y82jy6);
assign Y82jy6 = (~(S72jy6 | Pb8iw6));
assign Pb8iw6 = (!Toi7z6[2]);
assign S72jy6 = (~(W9v5z6 & Z98iw6));
assign Z98iw6 = (Eav5z6 & Qkfiy6);
assign Qkfiy6 = (~(Toi7z6[6] | Toi7z6[7]));
assign Eav5z6 = (~(Toi7z6[11] | Toi7z6[8]));
assign W9v5z6 = (Pi8iw6 & Cvfiy6);
assign Cvfiy6 = (!Toi7z6[10]);
assign Pi8iw6 = (~(Toi7z6[5] | Toi7z6[9]));
assign O9v5z6 = (R58iw6 & Bqi7z6[2]);
assign R58iw6 = (~(X22nv6 | Toi7z6[3]));
assign X22nv6 = (!Toi7z6[4]);
assign Pei7v6 = (P9get6 ? M5bdt6 : Jqj7z6[8]);
assign Iei7v6 = (Hr4yx6 ? Is5iw6 : Mqb7z6[0]);
assign Hr4yx6 = (Mav5z6 & Uav5z6);
assign Uav5z6 = (Cbv5z6 & Ihs7z6[1]);
assign Cbv5z6 = (Mq1jy6 & Hfryx6);
assign Mq1jy6 = (Kbv5z6 & Ihs7z6[0]);
assign Kbv5z6 = (~(L1syx6 | C397z6));
assign L1syx6 = (!Q097z6);
assign Mav5z6 = (Sbv5z6 & Zfs7z6[7]);
assign Sbv5z6 = (Ihs7z6[3] & Ihs7z6[2]);
assign Bei7v6 = (W92jy6 ? Is5iw6 : Ies7z6[16]);
assign W92jy6 = (Acv5z6 & Cv1jy6);
assign Cv1jy6 = (Icv5z6 & Hfryx6);
assign Hfryx6 = (~(O92jy6 | Mm27v6));
assign O92jy6 = (~(Qcv5z6 & Ycv5z6));
assign Ycv5z6 = (Tt4yx6 & Fgryx6);
assign Fgryx6 = (!Zfs7z6[8]);
assign Tt4yx6 = (!Tn27v6);
assign Qcv5z6 = (P7wyx6 & Xruyx6);
assign Xruyx6 = (!Ap27v6);
assign P7wyx6 = (~(Ohkhy6 | Or27v6));
assign Ohkhy6 = (!V0syx6);
assign V0syx6 = (Gdv5z6 & Odv5z6);
assign Odv5z6 = (~(Wdv5z6 | Hq27v6));
assign Wdv5z6 = (!Zfs7z6[10]);
assign Gdv5z6 = (Zfs7z6[9] & Zfs7z6[11]);
assign Icv5z6 = (Q097z6 & Pfryx6);
assign Pfryx6 = (!Zfs7z6[7]);
assign Acv5z6 = (Ihs7z6[2] & Eev5z6);
assign Eev5z6 = (~(C397z6 & Scs7z6[2]));
assign Udi7v6 = (O91jy6 ? Is5iw6 : Bfymz6[0]);
assign O91jy6 = (Xid8x6 & Fgpyx6);
assign Fgpyx6 = (D9pyx6 & P3xyx6);
assign Ndi7v6 = (Ua1jy6 ? Is5iw6 : Sgymz6[10]);
assign Ua1jy6 = (Xid8x6 & Ngpyx6);
assign Ngpyx6 = (Pbpyx6 & W5qhy6);
assign Pbpyx6 = (Mev5z6 & Xfymz6[4]);
assign Mev5z6 = (~(Eyyhy6 | Xfymz6[2]));
assign Gdi7v6 = (U61jy6 ? Is5iw6 : Ojymz6[10]);
assign U61jy6 = (Xid8x6 & Hfpyx6);
assign Hfpyx6 = (Kb1jy6 & D9pyx6);
assign D9pyx6 = (~(Uev5z6 | Xfymz6[2]));
assign Uev5z6 = (~(Eyyhy6 & J6yyx6));
assign Eyyhy6 = (!Xfymz6[3]);
assign Zci7v6 = (C71jy6 ? Is5iw6 : Blymz6[0]);
assign C71jy6 = (Xid8x6 & Lhpyx6);
assign Lhpyx6 = (Gthiw6 & W5qhy6);
assign W5qhy6 = (Cfv5z6 & Kfv5z6);
assign Cfv5z6 = (Mulhy6 & Xfymz6[8]);
assign Mulhy6 = (Sfv5z6 & Xfymz6[7]);
assign Sfv5z6 = (Xfymz6[6] & Xfymz6[5]);
assign Gthiw6 = (Agv5z6 & Xfymz6[4]);
assign Agv5z6 = (~(Xfymz6[2] | Xfymz6[3]));
assign Sci7v6 = (M61jy6 ? Is5iw6 : Unymz6[10]);
assign M61jy6 = (Xid8x6 & Thpyx6);
assign Thpyx6 = (Ied8x6 & P3xyx6);
assign P3xyx6 = (Igv5z6 & R6pyx6);
assign Igv5z6 = (!Qgv5z6);
assign Ied8x6 = (Ygv5z6 & Xfymz6[3]);
assign Ygv5z6 = (~(Xfymz6[2] | Xfymz6[4]));
assign Lci7v6 = (~(Ghv5z6 & Ohv5z6));
assign Ohv5z6 = (~(Whv5z6 & U42nv6));
assign U42nv6 = (~(Eiv5z6 & Miv5z6));
assign Miv5z6 = (~(Uiv5z6 & I8r7x6));
assign Eiv5z6 = (~(Itb7z6[0] & Cjv5z6));
assign Ghv5z6 = (~(Fjd7v6 & Kjv5z6));
assign Eci7v6 = (~(Sjv5z6 & Akv5z6));
assign Akv5z6 = (~(Whv5z6 & B52nv6));
assign B52nv6 = (~(Ikv5z6 & Qkv5z6));
assign Qkv5z6 = (~(Uiv5z6 & L7q7x6));
assign Ikv5z6 = (~(Itb7z6[1] & Cjv5z6));
assign Sjv5z6 = (~(Hcymz6[1] & Kjv5z6));
assign Xbi7v6 = (~(Ykv5z6 & Glv5z6));
assign Glv5z6 = (~(Whv5z6 & I52nv6));
assign I52nv6 = (~(Olv5z6 & Wlv5z6));
assign Wlv5z6 = (~(Uiv5z6 & Vcq7x6));
assign Olv5z6 = (~(Itb7z6[2] & Cjv5z6));
assign Whv5z6 = (Emv5z6 & Mmv5z6);
assign Emv5z6 = (!Kjv5z6);
assign Ykv5z6 = (~(Hcymz6[2] & Kjv5z6));
assign Qbi7v6 = (Kjv5z6 ? Hcymz6[3] : Umv5z6);
assign Umv5z6 = (~(Mmv5z6 & Pohov6));
assign Pohov6 = (!P52nv6);
assign Jbi7v6 = (Lhliw6 ? Tjr7z6[2] : ETMINTNUM[0]);
assign Cbi7v6 = (Lhliw6 ? Tjr7z6[9] : ETMINTNUM[7]);
assign Vai7v6 = (Lhliw6 ? Tjr7z6[8] : ETMINTNUM[6]);
assign Oai7v6 = (Lhliw6 ? Tjr7z6[7] : ETMINTNUM[5]);
assign Hai7v6 = (Lhliw6 ? Tjr7z6[5] : ETMINTNUM[3]);
assign Aai7v6 = (Lhliw6 ? Tjr7z6[3] : ETMINTNUM[1]);
assign T9i7v6 = (Nw5yx6 ? Gy2ft6 : Fw5yx6);
assign Fw5yx6 = (Id4ft6 ? U9p7z6[10] : U9p7z6[6]);
assign M9i7v6 = (O7fiw6 ? Hu2ft6 : Mbhiw6);
assign O7fiw6 = (Cnv5z6 & Q8fiw6);
assign Q8fiw6 = (~(Jsgiw6 & Hfqyx6));
assign Hfqyx6 = (~(Yglhy6 | Odlhy6));
assign Odlhy6 = (!Iw1jy6);
assign Iw1jy6 = (Knv5z6 & Gpeiy6);
assign Gpeiy6 = (Snv5z6 & Xueiw6);
assign Xueiw6 = (!Ah4ft6);
assign Snv5z6 = (!Nmq7z6[6]);
assign Knv5z6 = (Sz1jy6 & My1jy6);
assign My1jy6 = (!Nmq7z6[5]);
assign Sz1jy6 = (!Nmq7z6[3]);
assign Yglhy6 = (!Vcyyx6);
assign Vcyyx6 = (~(Nmq7z6[4] | E297z6));
assign Jsgiw6 = (Aj4ft6 & Cueiw6);
assign Cueiw6 = (!M297z6);
assign Cnv5z6 = (Nw5yx6 | Vw5yx6);
assign Vw5yx6 = (!Qb4ft6);
assign Nw5yx6 = (Kygnv6 | A9i8v6);
assign A9i8v6 = (Aov5z6 & Bq5yx6);
assign Aov5z6 = (~(Whhov6 | Oaadt6));
assign Whhov6 = (!Tlmov6);
assign Mbhiw6 = (W5q7z6[1] ? Qov5z6 : Iov5z6);
assign Qov5z6 = (W5q7z6[0] ? U9p7z6[28] : U9p7z6[26]);
assign Iov5z6 = (W5q7z6[0] & U9p7z6[24]);
assign F9i7v6 = (Yov5z6 | Op5ov6);
assign Yov5z6 = (B63yx6 ? F2f7v6 : Gpv5z6);
assign Gpv5z6 = (~(Opv5z6 & Wpv5z6));
assign Wpv5z6 = (~(Eqv5z6 & Mqv5z6));
assign Mqv5z6 = (Dxiyx6 | D53yx6);
assign Opv5z6 = (~(Dxiyx6 & Fo5ov6));
assign Y8i7v6 = (~(Uqv5z6 & Crv5z6));
assign Crv5z6 = (Zyiyx6 & Krv5z6);
assign Uqv5z6 = (Srv5z6 & Asv5z6);
assign Asv5z6 = (~(J7f7v6 & Isv5z6));
assign Isv5z6 = (~(Qsv5z6 & Ysv5z6));
assign Ysv5z6 = (Gtv5z6 | Otv5z6);
assign Gtv5z6 = (~(M8e7v6 | I6e7v6));
assign Srv5z6 = (~(Wtv5z6 & Mo5ov6));
assign Wtv5z6 = (~(Euv5z6 & Muv5z6));
assign Muv5z6 = (Uuv5z6 & Cvv5z6);
assign Cvv5z6 = (~(Kvv5z6 & L9e7v6));
assign Kvv5z6 = (I6e7v6 & Svv5z6);
assign Uuv5z6 = (Ju2yx6 & Awv5z6);
assign Awv5z6 = (!F2f7v6);
assign Euv5z6 = (~(D53yx6 | Fo5ov6));
assign R8i7v6 = (!Iwv5z6);
assign Iwv5z6 = (B63yx6 ? F8iyx6 : T5iyx6);
assign K8i7v6 = (Mo5ov6 ? Eqv5z6 : Qa2nz6[1]);
assign Eqv5z6 = (!Hp5ov6);
assign D8i7v6 = (!Qwv5z6);
assign Qwv5z6 = (Kf2nz6[0] ? Gxv5z6 : Ywv5z6);
assign Gxv5z6 = (Oxv5z6 & Wxv5z6);
assign Oxv5z6 = (Xjjyx6 & P7jyx6);
assign P7jyx6 = (!P3jyx6);
assign Xjjyx6 = (!Z6jyx6);
assign Z6jyx6 = (Iy1nz6[1] & M81nv6);
assign W7i7v6 = (~(Eyv5z6 & Myv5z6));
assign Myv5z6 = (~(P3jyx6 & Wxv5z6));
assign P3jyx6 = (Gie7v6 & M81nv6);
assign Eyv5z6 = (~(Uyv5z6 ^ Pfjyx6));
assign P7i7v6 = (~(Czv5z6 & Kzv5z6));
assign Kzv5z6 = (~(Kf2nz6[2] & Szv5z6));
assign Szv5z6 = (Uyv5z6 | Pfjyx6);
assign Pfjyx6 = (!Kf2nz6[1]);
assign Uyv5z6 = (~(Wxv5z6 & Kf2nz6[0]));
assign Czv5z6 = (~(T5jyx6 & Wxv5z6));
assign T5jyx6 = (A0w5z6 & Kf2nz6[1]);
assign A0w5z6 = (~(Dp2yx6 | Kf2nz6[2]));
assign Dp2yx6 = (!Kf2nz6[0]);
assign I7i7v6 = (D92nz6[0] ^ I0w5z6);
assign B7i7v6 = (~(Q0w5z6 & Y0w5z6));
assign Y0w5z6 = (~(I0w5z6 & Svv5z6));
assign Svv5z6 = (!Lb1nv6);
assign Lb1nv6 = (Ec2nz6[1] ? O1w5z6 : G1w5z6);
assign O1w5z6 = (Ec2nz6[0] & Otv5z6);
assign G1w5z6 = (W1w5z6 & Ns2yx6);
assign W1w5z6 = (~(Ec2nz6[2] | Ec2nz6[3]));
assign Q0w5z6 = (E2w5z6 ^ D92nz6[1]);
assign E2w5z6 = (~(I0w5z6 & D92nz6[0]));
assign I0w5z6 = (V91nv6 & Xrjyx6);
assign U6i7v6 = (Mo5ov6 ? Dxiyx6 : Qa2nz6[0]);
assign N6i7v6 = (Mo5ov6 ? M2w5z6 : A4f7v6);
assign Mo5ov6 = (!B63yx6);
assign M2w5z6 = (Vwiyx6 ? C3w5z6 : U2w5z6);
assign Vwiyx6 = (K3w5z6 & T5f7v6);
assign K3w5z6 = (Ec2nz6[0] & X7iyx6);
assign C3w5z6 = (S3w5z6 & Nwiyx6);
assign U2w5z6 = (Vp5ov6 & Hp5ov6);
assign G6i7v6 = (~(A4w5z6 & I4w5z6));
assign I4w5z6 = (Q4w5z6 | Ik77z6);
assign Q4w5z6 = (~(Vs2yx6 | Od77z6));
assign A4w5z6 = (~(Y4w5z6 & G5w5z6));
assign G5w5z6 = (O5w5z6 & W5w5z6);
assign W5w5z6 = (~(E6w5z6 & J23yx6));
assign E6w5z6 = (~(M6w5z6 & Ec2nz6[0]));
assign M6w5z6 = (R0f7v6 ? Op5ov6 : F8iyx6);
assign O5w5z6 = (U6w5z6 & X7iyx6);
assign U6w5z6 = (~(Qa2nz6[0] & Ns2yx6));
assign Y4w5z6 = (Qsv5z6 & H7iyx6);
assign Qsv5z6 = (~(B63yx6 | L5iyx6));
assign Z5i7v6 = (Lhliw6 ? Tjr7z6[4] : ETMINTNUM[2]);
assign Lhliw6 = (~(C7w5z6 & Xkq7z6[16]));
assign C7w5z6 = (HTMDHBURST[0] & Yohiy6);
assign Yohiy6 = (Ehliw6 | W3wnv6);
assign W3wnv6 = (!Skh7v6);
assign Ehliw6 = (!Zkh7v6);
assign S5i7v6 = (Kjv5z6 ? Hcymz6[4] : K7w5z6);
assign Kjv5z6 = (~(Xid8x6 & Hjpyx6));
assign Hjpyx6 = (S7w5z6 & A8w5z6);
assign A8w5z6 = (Xfymz6[2] & J6yyx6);
assign J6yyx6 = (!Xfymz6[4]);
assign S7w5z6 = (Kb1jy6 & Xfymz6[3]);
assign Kb1jy6 = (~(Qgv5z6 | R6pyx6));
assign R6pyx6 = (!Xfymz6[5]);
assign Qgv5z6 = (~(I8w5z6 & U6v5z6));
assign U6v5z6 = (Kfv5z6 & Ic2jy6);
assign Ic2jy6 = (!Xfymz6[7]);
assign Kfv5z6 = (Q8w5z6 & Sb2jy6);
assign Sb2jy6 = (!Xfymz6[10]);
assign Q8w5z6 = (~(Xfymz6[11] | Xfymz6[9]));
assign I8w5z6 = (Aslhy6 & I81jy6);
assign I81jy6 = (!Xfymz6[8]);
assign Aslhy6 = (!Xfymz6[6]);
assign Xid8x6 = (~(Yohiw6 | Xu67v6));
assign Yohiw6 = (!L877v6);
assign K7w5z6 = (~(Mmv5z6 & Zaeiw6));
assign Zaeiw6 = (!W52nv6);
assign Mmv5z6 = (Y8w5z6 & G9w5z6);
assign G9w5z6 = (V12nv6 & O9w5z6);
assign O9w5z6 = (W9w5z6 & I42jy6);
assign I42jy6 = (Gp1jy6 & Eaw5z6);
assign Eaw5z6 = (Maw5z6 & Uaw5z6);
assign Uaw5z6 = (M5giw6 & Wagiw6);
assign Wagiw6 = (!Ro3iw6);
assign Ro3iw6 = (~(Cbw5z6 & Kbw5z6));
assign Kbw5z6 = (~(Uiv5z6 & Vxq7x6));
assign Cbw5z6 = (~(Itb7z6[30] & Cjv5z6));
assign M5giw6 = (!E64iw6);
assign E64iw6 = (~(Sbw5z6 & Acw5z6));
assign Acw5z6 = (~(Uiv5z6 & Mbq7x6));
assign Sbw5z6 = (~(Itb7z6[26] & Cjv5z6));
assign Maw5z6 = (L1giw6 & U2giw6);
assign U2giw6 = (!Wf4iw6);
assign Wf4iw6 = (~(Icw5z6 & Qcw5z6));
assign Qcw5z6 = (~(Uiv5z6 & Yqonv6));
assign Icw5z6 = (~(Itb7z6[24] & Cjv5z6));
assign L1giw6 = (!Cx4iw6);
assign Cx4iw6 = (~(Ycw5z6 & Gdw5z6));
assign Gdw5z6 = (~(Uiv5z6 & Xzp7x6));
assign Ycw5z6 = (~(Itb7z6[23] & Cjv5z6));
assign Gp1jy6 = (Odw5z6 & D4giw6);
assign D4giw6 = (!Iklov6);
assign Iklov6 = (~(Wdw5z6 & Eew5z6));
assign Eew5z6 = (~(Uiv5z6 & C6q7x6));
assign Wdw5z6 = (~(Itb7z6[25] & Cjv5z6));
assign Odw5z6 = (V6giw6 & E8giw6);
assign E8giw6 = (!W14iw6);
assign W14iw6 = (~(Mew5z6 & Uew5z6));
assign Uew5z6 = (~(Uiv5z6 & Gmq7x6));
assign Mew5z6 = (~(Itb7z6[28] & Cjv5z6));
assign V6giw6 = (!H44iw6);
assign H44iw6 = (~(Cfw5z6 & Kfw5z6));
assign Kfw5z6 = (~(Uiv5z6 & Wgq7x6));
assign Cfw5z6 = (~(Itb7z6[27] & Cjv5z6));
assign W9w5z6 = (Tyfiw6 & Sfw5z6);
assign Sfw5z6 = (~(W52nv6 & P52nv6));
assign P52nv6 = (~(Agw5z6 & Igw5z6));
assign Igw5z6 = (~(Uiv5z6 & Fiq7x6));
assign Agw5z6 = (~(Itb7z6[3] & Cjv5z6));
assign W52nv6 = (~(Qgw5z6 & Ygw5z6));
assign Ygw5z6 = (~(Uiv5z6 & Pnq7x6));
assign Qgw5z6 = (~(Itb7z6[4] & Cjv5z6));
assign Tyfiw6 = (!Ej5iw6);
assign Ej5iw6 = (~(Ghw5z6 & Ohw5z6));
assign Ohw5z6 = (~(Uiv5z6 & Mpq7x6));
assign Ghw5z6 = (~(Itb7z6[21] & Cjv5z6));
assign V12nv6 = (Umhiw6 & Whw5z6);
assign Whw5z6 = (Eiw5z6 & Miw5z6);
assign Miw5z6 = (Wifiw6 & Nhfiw6);
assign Nhfiw6 = (!U47iw6);
assign U47iw6 = (~(Uiw5z6 & Cjw5z6));
assign Cjw5z6 = (~(Uiv5z6 & Kqonv6));
assign Uiw5z6 = (~(Itb7z6[8] & Cjv5z6));
assign Wifiw6 = (!J27iw6);
assign J27iw6 = (~(Kjw5z6 & Sjw5z6));
assign Sjw5z6 = (~(Uiv5z6 & H5q7x6));
assign Kjw5z6 = (~(Itb7z6[9] & Cjv5z6));
assign Eiw5z6 = (N9giw6 & Fcgiw6);
assign Fcgiw6 = (!X0hov6);
assign X0hov6 = (~(Akw5z6 & Ikw5z6));
assign Ikw5z6 = (~(Uiv5z6 & Ht1ov6));
assign Akw5z6 = (~(Itb7z6[31] & Cjv5z6));
assign N9giw6 = (!Zz3iw6);
assign Zz3iw6 = (~(Qkw5z6 & Ykw5z6));
assign Ykw5z6 = (~(Uiv5z6 & Qrq7x6));
assign Qkw5z6 = (~(Itb7z6[29] & Cjv5z6));
assign Umhiw6 = (Xmfiw6 & C0giw6);
assign C0giw6 = (!D85iw6);
assign D85iw6 = (~(Glw5z6 & Olw5z6));
assign Olw5z6 = (~(Uiv5z6 & Wuq7x6));
assign Glw5z6 = (~(Itb7z6[22] & Cjv5z6));
assign Xmfiw6 = (!Emhov6);
assign Emhov6 = (~(Wlw5z6 & Emw5z6));
assign Emw5z6 = (~(Uiv5z6 & Llq7x6));
assign Wlw5z6 = (~(Itb7z6[12] & Cjv5z6));
assign Y8w5z6 = (Mmw5z6 & Umw5z6);
assign Umw5z6 = (Z32nv6 & Egfiw6);
assign Egfiw6 = (!R62nv6);
assign R62nv6 = (~(Cnw5z6 & Knw5z6));
assign Knw5z6 = (~(Uiv5z6 & Kwp7x6));
assign Cnw5z6 = (~(Itb7z6[7] & Cjv5z6));
assign Z32nv6 = (~(Snw5z6 | Aow5z6));
assign Aow5z6 = (~(Iow5z6 & Qow5z6));
assign Qow5z6 = (Yow5z6 & Oyhov6);
assign Oyhov6 = (!Gr5iw6);
assign Gr5iw6 = (~(Gpw5z6 & Opw5z6));
assign Opw5z6 = (~(Uiv5z6 & Y3q7x6));
assign Gpw5z6 = (~(Itb7z6[17] & Cjv5z6));
assign Yow5z6 = (Kxfiw6 & Bwfiw6);
assign Bwfiw6 = (!Mn5iw6);
assign Mn5iw6 = (~(Wpw5z6 & Eqw5z6));
assign Eqw5z6 = (~(Uiv5z6 & Seq7x6));
assign Wpw5z6 = (~(Itb7z6[19] & Cjv5z6));
assign Kxfiw6 = (!Bl5iw6);
assign Bl5iw6 = (~(Mqw5z6 & Uqw5z6));
assign Uqw5z6 = (~(Uiv5z6 & Ckq7x6));
assign Mqw5z6 = (~(Itb7z6[20] & Cjv5z6));
assign Iow5z6 = (Hsfiw6 & Sufiw6);
assign Sufiw6 = (!Jp5iw6);
assign Jp5iw6 = (~(Crw5z6 & Krw5z6));
assign Krw5z6 = (~(Uiv5z6 & I9q7x6));
assign Crw5z6 = (~(Itb7z6[18] & Cjv5z6));
assign Hsfiw6 = (!Is5iw6);
assign Is5iw6 = (~(Srw5z6 & Asw5z6));
assign Asw5z6 = (~(Uiv5z6 & V4r7x6));
assign Srw5z6 = (~(Itb7z6[16] & Cjv5z6));
assign Snw5z6 = (~(Isw5z6 & Qsw5z6));
assign Qsw5z6 = (Ysw5z6 & Gofiw6);
assign Gofiw6 = (!Guhov6);
assign Guhov6 = (~(Gtw5z6 & Otw5z6));
assign Otw5z6 = (~(Uiv5z6 & Vqq7x6));
assign Gtw5z6 = (~(Itb7z6[13] & Cjv5z6));
assign Ysw5z6 = (Yqfiw6 & Ppfiw6);
assign Ppfiw6 = (!Bk6iw6);
assign Bk6iw6 = (~(Wtw5z6 & Euw5z6));
assign Euw5z6 = (~(Uiv5z6 & Twq7x6));
assign Wtw5z6 = (~(Itb7z6[14] & Cjv5z6));
assign Yqfiw6 = (!Z0iov6);
assign Z0iov6 = (~(Muw5z6 & Uuw5z6));
assign Uuw5z6 = (~(Uiv5z6 & Oyp7x6));
assign Muw5z6 = (~(Itb7z6[15] & Cjv5z6));
assign Isw5z6 = (Olfiw6 & Fkfiw6);
assign Fkfiw6 = (!H17iw6);
assign H17iw6 = (~(Cvw5z6 & Kvw5z6));
assign Kvw5z6 = (~(Uiv5z6 & Raq7x6));
assign Cvw5z6 = (~(Itb7z6[10] & Cjv5z6));
assign Olfiw6 = (!Dz6iw6);
assign Dz6iw6 = (~(Svw5z6 & Aww5z6));
assign Aww5z6 = (~(Uiv5z6 & Bgq7x6));
assign Svw5z6 = (~(Itb7z6[11] & Cjv5z6));
assign Mmw5z6 = (Gbeiw6 & Tdfiw6);
assign Tdfiw6 = (!D62nv6);
assign D62nv6 = (~(Iww5z6 & Qww5z6));
assign Qww5z6 = (~(Uiv5z6 & Zsq7x6));
assign Iww5z6 = (~(Itb7z6[5] & Cjv5z6));
assign Gbeiw6 = (!K62nv6);
assign K62nv6 = (~(Yww5z6 & Gxw5z6));
assign Gxw5z6 = (~(Uiv5z6 & Lzq7x6));
assign Uiv5z6 = (C1o7z6[0] & Q497z6);
assign Yww5z6 = (~(Itb7z6[6] & Cjv5z6));
assign Cjv5z6 = (C1o7z6[1] & Q497z6);
assign L5i7v6 = (Zmbyx6 ? Vcxmz6[0] : TSVALUEB[0]);
assign E5i7v6 = (Zmbyx6 ? Vcxmz6[47] : TSVALUEB[47]);
assign X4i7v6 = (Zmbyx6 ? Vcxmz6[46] : TSVALUEB[46]);
assign Q4i7v6 = (Zmbyx6 ? Vcxmz6[45] : TSVALUEB[45]);
assign J4i7v6 = (Zmbyx6 ? Vcxmz6[44] : TSVALUEB[44]);
assign C4i7v6 = (Zmbyx6 ? Vcxmz6[43] : TSVALUEB[43]);
assign V3i7v6 = (Zmbyx6 ? Vcxmz6[42] : TSVALUEB[42]);
assign O3i7v6 = (Zmbyx6 ? Vcxmz6[41] : TSVALUEB[41]);
assign H3i7v6 = (Zmbyx6 ? Vcxmz6[40] : TSVALUEB[40]);
assign A3i7v6 = (Zmbyx6 ? Vcxmz6[39] : TSVALUEB[39]);
assign T2i7v6 = (Zmbyx6 ? Vcxmz6[38] : TSVALUEB[38]);
assign M2i7v6 = (Zmbyx6 ? Vcxmz6[37] : TSVALUEB[37]);
assign F2i7v6 = (Zmbyx6 ? Vcxmz6[36] : TSVALUEB[36]);
assign Y1i7v6 = (Zmbyx6 ? Vcxmz6[35] : TSVALUEB[35]);
assign R1i7v6 = (Zmbyx6 ? Vcxmz6[34] : TSVALUEB[34]);
assign K1i7v6 = (Zmbyx6 ? Vcxmz6[33] : TSVALUEB[33]);
assign D1i7v6 = (Zmbyx6 ? Vcxmz6[32] : TSVALUEB[32]);
assign W0i7v6 = (Zmbyx6 ? Vcxmz6[31] : TSVALUEB[31]);
assign P0i7v6 = (Zmbyx6 ? Vcxmz6[30] : TSVALUEB[30]);
assign I0i7v6 = (Zmbyx6 ? Vcxmz6[29] : TSVALUEB[29]);
assign B0i7v6 = (Zmbyx6 ? Vcxmz6[28] : TSVALUEB[28]);
assign Uzh7v6 = (Zmbyx6 ? Vcxmz6[27] : TSVALUEB[27]);
assign Nzh7v6 = (Zmbyx6 ? Vcxmz6[26] : TSVALUEB[26]);
assign Gzh7v6 = (Zmbyx6 ? Vcxmz6[25] : TSVALUEB[25]);
assign Zyh7v6 = (Zmbyx6 ? Vcxmz6[24] : TSVALUEB[24]);
assign Syh7v6 = (Zmbyx6 ? Vcxmz6[23] : TSVALUEB[23]);
assign Lyh7v6 = (Zmbyx6 ? Vcxmz6[22] : TSVALUEB[22]);
assign Eyh7v6 = (Zmbyx6 ? Vcxmz6[21] : TSVALUEB[21]);
assign Xxh7v6 = (Zmbyx6 ? Vcxmz6[20] : TSVALUEB[20]);
assign Qxh7v6 = (Zmbyx6 ? Vcxmz6[19] : TSVALUEB[19]);
assign Jxh7v6 = (Zmbyx6 ? Vcxmz6[18] : TSVALUEB[18]);
assign Cxh7v6 = (Zmbyx6 ? Vcxmz6[17] : TSVALUEB[17]);
assign Vwh7v6 = (Zmbyx6 ? Vcxmz6[16] : TSVALUEB[16]);
assign Owh7v6 = (Zmbyx6 ? Vcxmz6[15] : TSVALUEB[15]);
assign Hwh7v6 = (Zmbyx6 ? Vcxmz6[14] : TSVALUEB[14]);
assign Awh7v6 = (Zmbyx6 ? Vcxmz6[13] : TSVALUEB[13]);
assign Tvh7v6 = (Zmbyx6 ? Vcxmz6[12] : TSVALUEB[12]);
assign Mvh7v6 = (Zmbyx6 ? Vcxmz6[11] : TSVALUEB[11]);
assign Fvh7v6 = (Zmbyx6 ? Vcxmz6[10] : TSVALUEB[10]);
assign Yuh7v6 = (Zmbyx6 ? Vcxmz6[9] : TSVALUEB[9]);
assign Ruh7v6 = (Zmbyx6 ? Vcxmz6[8] : TSVALUEB[8]);
assign Kuh7v6 = (Zmbyx6 ? Vcxmz6[7] : TSVALUEB[7]);
assign Duh7v6 = (Zmbyx6 ? Vcxmz6[6] : TSVALUEB[6]);
assign Wth7v6 = (Zmbyx6 ? Vcxmz6[5] : TSVALUEB[5]);
assign Pth7v6 = (Zmbyx6 ? Vcxmz6[4] : TSVALUEB[4]);
assign Zmbyx6 = (!Oxw5z6);
assign Ith7v6 = (Oxw5z6 ? TSVALUEB[3] : Vcxmz6[3]);
assign Bth7v6 = (Oxw5z6 ? TSVALUEB[2] : Vcxmz6[2]);
assign Ush7v6 = (Oxw5z6 ? TSVALUEB[1] : Vcxmz6[1]);
assign Oxw5z6 = (Wxw5z6 & Fho7v6);
assign Fho7v6 = (I96ft6 | D5byx6);
assign D5byx6 = (D86ft6 & Eyw5z6);
assign Eyw5z6 = (~(Myw5z6 & Uyw5z6));
assign Uyw5z6 = (~(Uur7z6[1] | Hsr7z6[1]));
assign Myw5z6 = (Eixiy6 & Nc5yx6);
assign Nc5yx6 = (!C4s7z6[1]);
assign Eixiy6 = (~(Ixr7z6[1] | Xwadt6));
assign Wxw5z6 = (~(Ak77z6 | Fbxmz6[3]));
assign Nsh7v6 = (Vjqnv6 ? J0n7z6[0] : Gfqnv6);
assign Gsh7v6 = (~(Czw5z6 & Kzw5z6));
assign Kzw5z6 = (~(J72nz6[7] & Szw5z6));
assign Czw5z6 = (A0x5z6 & I0x5z6);
assign I0x5z6 = (~(Q0x5z6 & Y0x5z6));
assign Q0x5z6 = (G1x5z6 & O1x5z6);
assign O1x5z6 = (W1x5z6 | E2x5z6);
assign G1x5z6 = (W1x5z6 | Au1nz6[7]);
assign W1x5z6 = (~(M2x5z6 & U2x5z6));
assign U2x5z6 = (~(Qq5ov6 & Zs1nz6[7]));
assign M2x5z6 = (C3x5z6 & K3x5z6);
assign K3x5z6 = (~(S3x5z6 & Yr1nz6[7]));
assign C3x5z6 = (~(Jq5ov6 & Xq1nz6[7]));
assign A0x5z6 = (L53yx6 | Zijyx6);
assign Zijyx6 = (A4x5z6 & I4x5z6);
assign I4x5z6 = (Q4x5z6 & Y4x5z6);
assign Y4x5z6 = (~(G5x5z6 & Mm1nz6[7]));
assign Q4x5z6 = (~(O5x5z6 & Oo1nz6[7]));
assign A4x5z6 = (W5x5z6 & E6x5z6);
assign E6x5z6 = (~(Z63yx6 & Kh1nz6[7]));
assign W5x5z6 = (~(H73yx6 & Nn1nz6[7]));
assign Zrh7v6 = (~(M6x5z6 & U6x5z6));
assign U6x5z6 = (~(J72nz6[2] & Szw5z6));
assign M6x5z6 = (C7x5z6 & K7x5z6);
assign K7x5z6 = (~(Y0x5z6 & S7x5z6));
assign S7x5z6 = (~(A8x5z6 & I8x5z6));
assign I8x5z6 = (Q8x5z6 & Y8x5z6);
assign Y8x5z6 = (~(S3x5z6 & Yr1nz6[2]));
assign Q8x5z6 = (~(E2x5z6 & Au1nz6[2]));
assign A8x5z6 = (G9x5z6 & O9x5z6);
assign O9x5z6 = (~(Jq5ov6 & Xq1nz6[2]));
assign G9x5z6 = (~(Qq5ov6 & Zs1nz6[2]));
assign C7x5z6 = (L53yx6 | Fojyx6);
assign Fojyx6 = (W9x5z6 & Eax5z6);
assign Eax5z6 = (Max5z6 & Uax5z6);
assign Uax5z6 = (~(G5x5z6 & Mm1nz6[2]));
assign Max5z6 = (~(O5x5z6 & Oo1nz6[2]));
assign W9x5z6 = (Cbx5z6 & Kbx5z6);
assign Kbx5z6 = (~(Z63yx6 & Kh1nz6[2]));
assign Cbx5z6 = (~(H73yx6 & Nn1nz6[2]));
assign Srh7v6 = (~(Sbx5z6 & Acx5z6));
assign Acx5z6 = (~(J72nz6[3] & Szw5z6));
assign Sbx5z6 = (Icx5z6 & Qcx5z6);
assign Qcx5z6 = (~(Y0x5z6 & Ycx5z6));
assign Ycx5z6 = (~(Gdx5z6 & Odx5z6));
assign Odx5z6 = (Wdx5z6 & Eex5z6);
assign Eex5z6 = (~(S3x5z6 & Yr1nz6[3]));
assign Wdx5z6 = (~(E2x5z6 & Au1nz6[3]));
assign Gdx5z6 = (Mex5z6 & Uex5z6);
assign Uex5z6 = (~(Jq5ov6 & Xq1nz6[3]));
assign Mex5z6 = (~(Qq5ov6 & Zs1nz6[3]));
assign Icx5z6 = (L53yx6 | Lhjyx6);
assign Lhjyx6 = (Cfx5z6 & Kfx5z6);
assign Kfx5z6 = (Sfx5z6 & Agx5z6);
assign Agx5z6 = (~(G5x5z6 & Mm1nz6[3]));
assign Sfx5z6 = (~(O5x5z6 & Oo1nz6[3]));
assign Cfx5z6 = (Igx5z6 & Qgx5z6);
assign Qgx5z6 = (~(Z63yx6 & Kh1nz6[3]));
assign Igx5z6 = (~(H73yx6 & Nn1nz6[3]));
assign Lrh7v6 = (~(Ygx5z6 & Ghx5z6));
assign Ghx5z6 = (~(J72nz6[5] & Szw5z6));
assign Ygx5z6 = (Ohx5z6 & Whx5z6);
assign Whx5z6 = (~(Y0x5z6 & Eix5z6));
assign Eix5z6 = (~(Mix5z6 & Uix5z6));
assign Uix5z6 = (Cjx5z6 & Kjx5z6);
assign Kjx5z6 = (~(S3x5z6 & Yr1nz6[5]));
assign Cjx5z6 = (~(E2x5z6 & Au1nz6[5]));
assign Mix5z6 = (Sjx5z6 & Akx5z6);
assign Akx5z6 = (~(Jq5ov6 & Xq1nz6[5]));
assign Sjx5z6 = (~(Qq5ov6 & Zs1nz6[5]));
assign Ohx5z6 = (L53yx6 | Ddjyx6);
assign Ddjyx6 = (Ikx5z6 & Qkx5z6);
assign Qkx5z6 = (Ykx5z6 & Glx5z6);
assign Glx5z6 = (~(G5x5z6 & Mm1nz6[5]));
assign Ykx5z6 = (~(O5x5z6 & Oo1nz6[5]));
assign Ikx5z6 = (Olx5z6 & Wlx5z6);
assign Wlx5z6 = (~(Z63yx6 & Kh1nz6[5]));
assign Olx5z6 = (~(H73yx6 & Nn1nz6[5]));
assign Erh7v6 = (~(Emx5z6 & Mmx5z6));
assign Mmx5z6 = (~(J72nz6[0] & Szw5z6));
assign Emx5z6 = (Umx5z6 & Cnx5z6);
assign Cnx5z6 = (~(Y0x5z6 & Knx5z6));
assign Knx5z6 = (~(Snx5z6 & Aox5z6));
assign Aox5z6 = (Iox5z6 & Qox5z6);
assign Qox5z6 = (~(S3x5z6 & Yr1nz6[0]));
assign Iox5z6 = (~(E2x5z6 & Au1nz6[0]));
assign Snx5z6 = (Yox5z6 & Gpx5z6);
assign Gpx5z6 = (~(Jq5ov6 & Bv1nz6[0]));
assign Yox5z6 = (~(Qq5ov6 & Zs1nz6[0]));
assign Umx5z6 = (L53yx6 | Hrjyx6);
assign Hrjyx6 = (Opx5z6 & Wpx5z6);
assign Wpx5z6 = (Eqx5z6 & Mqx5z6);
assign Mqx5z6 = (~(G5x5z6 & Mm1nz6[0]));
assign Eqx5z6 = (~(O5x5z6 & Oo1nz6[0]));
assign Opx5z6 = (Uqx5z6 & Crx5z6);
assign Crx5z6 = (~(Z63yx6 & Pp1nz6[0]));
assign Uqx5z6 = (~(H73yx6 & Nn1nz6[0]));
assign Xqh7v6 = (Dt2yx6 ? N52nz6[5] : N52nz6[6]);
assign Qqh7v6 = (Dt2yx6 ? N52nz6[4] : N52nz6[5]);
assign Jqh7v6 = (Dt2yx6 ? N52nz6[3] : N52nz6[4]);
assign Cqh7v6 = (Dt2yx6 ? N52nz6[2] : N52nz6[3]);
assign Vph7v6 = (Dt2yx6 ? N52nz6[1] : N52nz6[2]);
assign Oph7v6 = (Dt2yx6 ? N52nz6[0] : N52nz6[1]);
assign Dt2yx6 = (!Krx5z6);
assign Hph7v6 = (Krx5z6 ? N52nz6[0] : Wye7v6);
assign Krx5z6 = (~(Vs2yx6 | Ns2yx6));
assign Vs2yx6 = (~(Srx5z6 & Bejyx6));
assign Bejyx6 = (~(Xrjyx6 | B63yx6));
assign Srx5z6 = (V91nv6 & J7f7v6);
assign Aph7v6 = (Vjqnv6 ? J0n7z6[1] : Qdqnv6);
assign Vjqnv6 = (!Gmnet6);
assign Toh7v6 = (~(Asx5z6 & Isx5z6));
assign Isx5z6 = (~(J72nz6[4] & Szw5z6));
assign Asx5z6 = (Qsx5z6 & Ysx5z6);
assign Ysx5z6 = (~(Y0x5z6 & Gtx5z6));
assign Gtx5z6 = (~(Otx5z6 & Wtx5z6));
assign Wtx5z6 = (Eux5z6 & Mux5z6);
assign Mux5z6 = (~(S3x5z6 & Yr1nz6[4]));
assign Eux5z6 = (~(E2x5z6 & Au1nz6[4]));
assign Otx5z6 = (Uux5z6 & Cvx5z6);
assign Cvx5z6 = (~(Jq5ov6 & Xq1nz6[4]));
assign Uux5z6 = (~(Qq5ov6 & Zs1nz6[4]));
assign Qsx5z6 = (L53yx6 | Bqjyx6);
assign Bqjyx6 = (Kvx5z6 & Svx5z6);
assign Svx5z6 = (Awx5z6 & Iwx5z6);
assign Iwx5z6 = (~(G5x5z6 & Mm1nz6[4]));
assign Awx5z6 = (~(O5x5z6 & Oo1nz6[4]));
assign Kvx5z6 = (Qwx5z6 & Ywx5z6);
assign Ywx5z6 = (~(Z63yx6 & Kh1nz6[4]));
assign Qwx5z6 = (~(H73yx6 & Nn1nz6[4]));
assign Moh7v6 = (~(Gxx5z6 & Oxx5z6));
assign Oxx5z6 = (~(J72nz6[6] & Szw5z6));
assign Gxx5z6 = (Wxx5z6 & Eyx5z6);
assign Eyx5z6 = (~(Y0x5z6 & Myx5z6));
assign Myx5z6 = (~(Uyx5z6 & Czx5z6));
assign Czx5z6 = (Kzx5z6 & Szx5z6);
assign Szx5z6 = (~(S3x5z6 & Yr1nz6[6]));
assign Kzx5z6 = (~(E2x5z6 & Au1nz6[6]));
assign Uyx5z6 = (A0y5z6 & I0y5z6);
assign I0y5z6 = (~(Jq5ov6 & Xq1nz6[6]));
assign A0y5z6 = (~(Qq5ov6 & Zs1nz6[6]));
assign Wxx5z6 = (~(Q0y5z6 & Zmjyx6));
assign Zmjyx6 = (~(Y0y5z6 & G1y5z6));
assign G1y5z6 = (O1y5z6 & W1y5z6);
assign W1y5z6 = (~(G5x5z6 & Mm1nz6[6]));
assign O1y5z6 = (~(O5x5z6 & Oo1nz6[6]));
assign Y0y5z6 = (E2y5z6 & M2y5z6);
assign M2y5z6 = (~(Z63yx6 & Kh1nz6[6]));
assign E2y5z6 = (~(H73yx6 & Nn1nz6[6]));
assign Foh7v6 = (Cxtet6 & Mr9ov6);
assign Ynh7v6 = (Dztet6 & Mr9ov6);
assign Mr9ov6 = (H2kiw6 | F4xnv6);
assign F4xnv6 = (~(H11ov6 & Kconv6));
assign H11ov6 = (Ccnet6 & Rconv6);
assign Rconv6 = (~(U2y5z6 & C3y5z6));
assign C3y5z6 = (K3y5z6 & S3y5z6);
assign S3y5z6 = (~(G7piw6 & HREADYS));
assign K3y5z6 = (A4y5z6 & Kfliy6);
assign Kfliy6 = (~(Kqm7z6[2] & I4y5z6));
assign A4y5z6 = (~(HREADYI & Q4y5z6));
assign Q4y5z6 = (~(Y4y5z6 & Ealiy6));
assign Ealiy6 = (!R9piw6);
assign R9piw6 = (Kqm7z6[0] & I4y5z6);
assign Y4y5z6 = (~(G5y5z6 & Cfliy6));
assign G5y5z6 = (~(G7piw6 | K9piw6));
assign G7piw6 = (Kqm7z6[1] & I4y5z6);
assign I4y5z6 = (Cfliy6 & O5y5z6);
assign U2y5z6 = (X0oet6 & W5y5z6);
assign W5y5z6 = (~(K9piw6 & Q0ziy6));
assign Q0ziy6 = (!E6y5z6);
assign K9piw6 = (M6y5z6 & Cfliy6);
assign M6y5z6 = (!O5y5z6);
assign O5y5z6 = (Cakiw6 | U6y5z6);
assign H2kiw6 = (~(C7y5z6 & K7y5z6));
assign K7y5z6 = (~(Ogkiw6 & S7y5z6));
assign S7y5z6 = (~(A8y5z6 & Vd1ft6));
assign A8y5z6 = (I8y5z6 & Dm1ft6);
assign Ogkiw6 = (Q8y5z6 & Y8y5z6);
assign Y8y5z6 = (~(D7gxx6 | S4gxx6));
assign S4gxx6 = (!U5gxx6);
assign U5gxx6 = (~(G9y5z6 & Pg1ft6));
assign G9y5z6 = (I8y5z6 & Hq1ft6);
assign D7gxx6 = (O9y5z6 & Te1ft6);
assign O9y5z6 = (I8y5z6 & Nn1ft6);
assign Q8y5z6 = (Z4gxx6 & W6gxx6);
assign W6gxx6 = (~(W9y5z6 & Rf1ft6));
assign W9y5z6 = (I8y5z6 & Xo1ft6);
assign Z4gxx6 = (Eay5z6 & E4gxx6);
assign E4gxx6 = (!Mfkiw6);
assign Mfkiw6 = (May5z6 & Li1ft6);
assign May5z6 = (I8y5z6 & Iv1ft6);
assign Eay5z6 = (~(Uay5z6 & Nh1ft6));
assign Uay5z6 = (I8y5z6 & Rr1ft6);
assign I8y5z6 = (Lbkiw6 & Zy1ft6);
assign C7y5z6 = (Kconv6 & Cby5z6);
assign Cby5z6 = (!Dconv6);
assign Dconv6 = (Ccnet6 & Y3xnv6);
assign Y3xnv6 = (~(Kby5z6 & Sby5z6));
assign Sby5z6 = (~(Acy5z6 & Icy5z6));
assign Acy5z6 = (Am1ov6 & Qcy5z6);
assign Qcy5z6 = (~(Ycy5z6 & Ikyiy6));
assign Ycy5z6 = (Ody5z6 ? Gdy5z6 : N0nyx6);
assign Gdy5z6 = (Wdy5z6 & Eey5z6);
assign Eey5z6 = (Mey5z6 & Uey5z6);
assign Uey5z6 = (Cfy5z6 & Kfy5z6);
assign Kfy5z6 = (~(Ltnyx6 & Zlk7z6[23]));
assign Cfy5z6 = (~(Nsnyx6 & Hwk7z6[23]));
assign Mey5z6 = (Sfy5z6 & Agy5z6);
assign Agy5z6 = (~(Junyx6 & P6l7z6[23]));
assign Sfy5z6 = (~(Runyx6 & Xgl7z6[23]));
assign Wdy5z6 = (Igy5z6 & Qgy5z6);
assign Qgy5z6 = (Ygy5z6 & Ghy5z6);
assign Ghy5z6 = (~(Fwnyx6 & Frl7z6[23]));
assign Ygy5z6 = (~(Nwnyx6 & N1m7z6[23]));
assign Igy5z6 = (Ohy5z6 & Why5z6);
assign Why5z6 = (~(Lxnyx6 & Rbk7z6[23]));
assign Ohy5z6 = (~(Txnyx6 & Vbm7z6[23]));
assign N0nyx6 = (~(Xnmyx6 & Eiy5z6));
assign Eiy5z6 = (~(Bkfnv6 & Eg3nv6));
assign Kby5z6 = (~(Miy5z6 & Am1ov6));
assign Miy5z6 = (Uiy5z6 & X3nyx6);
assign X3nyx6 = (!Hnmyx6);
assign Hnmyx6 = (~(Cjy5z6 | Ltmyx6));
assign Ltmyx6 = (Icy5z6 & Ody5z6);
assign Cjy5z6 = (Kjy5z6 & Sjy5z6);
assign Kjy5z6 = (Icy5z6 & Aky5z6);
assign Aky5z6 = (~(Apget6 & HPROTI[1]));
assign Icy5z6 = (!HPROTI[0]);
assign HPROTI[0] = (Crcdt6 ? Fsc7z6[0] : Emoov6);
assign Uiy5z6 = (~(Iky5z6 & Ody5z6));
assign Ody5z6 = (~(Lxnyx6 & Qky5z6));
assign Qky5z6 = (~(Yky5z6 & Gly5z6));
assign Gly5z6 = (Oly5z6 & Wly5z6);
assign Wly5z6 = (Emy5z6 & Mmy5z6);
assign Mmy5z6 = (Umy5z6 & Cny5z6);
assign Cny5z6 = (~(C4het6 | Kny5z6));
assign Kny5z6 = (Sny5z6 & Jienv6);
assign Sny5z6 = (Az3nv6 ^ Aoy5z6);
assign Umy5z6 = (Ioy5z6 & Qoy5z6);
assign Qoy5z6 = (~(Yoy5z6 & O3env6));
assign Yoy5z6 = (HADDRI[7] ^ Dfk7z6[7]);
assign Ioy5z6 = (~(Gpy5z6 & Cbenv6));
assign Gpy5z6 = (HADDRI[6] ^ Dfk7z6[6]);
assign Emy5z6 = (Opy5z6 & Wpy5z6);
assign Wpy5z6 = (Eqy5z6 & Mqy5z6);
assign Mqy5z6 = (~(Uqy5z6 & Nrenv6));
assign Uqy5z6 = (HADDRI[15] ^ Dfk7z6[15]);
assign Eqy5z6 = (~(Cry5z6 & Qwenv6));
assign Cry5z6 = (HADDRI[14] ^ Dfk7z6[14]);
assign Opy5z6 = (Kry5z6 & Sry5z6);
assign Sry5z6 = (~(Asy5z6 & H3env6));
assign Asy5z6 = (HADDRI[13] ^ Dfk7z6[13]);
assign Kry5z6 = (~(Isy5z6 & Vaenv6));
assign Isy5z6 = (HADDRI[12] ^ Dfk7z6[12]);
assign Oly5z6 = (Qsy5z6 & Ysy5z6);
assign Ysy5z6 = (Gty5z6 & Oty5z6);
assign Oty5z6 = (Wty5z6 & Euy5z6);
assign Euy5z6 = (~(Muy5z6 & Qienv6));
assign Muy5z6 = (HADDRI[11] ^ Dfk7z6[11]);
assign Wty5z6 = (~(Uuy5z6 & Fnenv6));
assign Uuy5z6 = (HADDRI[10] ^ Dfk7z6[10]);
assign Gty5z6 = (Cvy5z6 & Kvy5z6);
assign Kvy5z6 = (~(Svy5z6 & Awy5z6));
assign Svy5z6 = (HADDRI[9] ^ Dfk7z6[9]);
assign Cvy5z6 = (~(Iwy5z6 & Cienv6));
assign Iwy5z6 = (HADDRI[8] ^ Dfk7z6[8]);
assign Qsy5z6 = (Qwy5z6 & Ywy5z6);
assign Ywy5z6 = (~(Gxy5z6 & Peenv6));
assign Gxy5z6 = (Dfk7z6[29] ^ Bkfnv6);
assign Qwy5z6 = (Oxy5z6 & Wxy5z6);
assign Wxy5z6 = (~(Eyy5z6 & Nzdnv6));
assign Eyy5z6 = (Njfnv6 ^ Dfk7z6[31]);
assign Oxy5z6 = (~(Myy5z6 & B7env6));
assign Myy5z6 = (Ujfnv6 ^ Dfk7z6[30]);
assign Yky5z6 = (Uyy5z6 & Czy5z6);
assign Czy5z6 = (Kzy5z6 & Szy5z6);
assign Szy5z6 = (A0z5z6 & I0z5z6);
assign I0z5z6 = (Q0z5z6 & Y0z5z6);
assign Y0z5z6 = (~(G1z5z6 & O1z5z6));
assign G1z5z6 = (HADDRI[28] ^ Dfk7z6[28]);
assign Q0z5z6 = (~(W1z5z6 & Dtenv6));
assign W1z5z6 = (HADDRI[27] ^ Dfk7z6[27]);
assign A0z5z6 = (E2z5z6 & M2z5z6);
assign M2z5z6 = (~(U2z5z6 & K0fnv6));
assign U2z5z6 = (HADDRI[26] ^ Dfk7z6[26]);
assign E2z5z6 = (~(C3z5z6 & K1env6));
assign C3z5z6 = (HADDRI[25] ^ Dfk7z6[25]);
assign Kzy5z6 = (K3z5z6 & S3z5z6);
assign S3z5z6 = (~(A4z5z6 & Wlenv6));
assign A4z5z6 = (HADDRI[22] ^ Dfk7z6[22]);
assign K3z5z6 = (I4z5z6 & Q4z5z6);
assign Q4z5z6 = (~(Y4z5z6 & Y8env6));
assign Y4z5z6 = (HADDRI[24] ^ Dfk7z6[24]);
assign I4z5z6 = (~(G5z5z6 & Mgenv6));
assign G5z5z6 = (HADDRI[23] ^ Dfk7z6[23]);
assign Uyy5z6 = (O5z5z6 & W5z5z6);
assign W5z5z6 = (E6z5z6 & M6z5z6);
assign M6z5z6 = (U6z5z6 & C7z5z6);
assign C7z5z6 = (~(K7z5z6 & Grenv6));
assign K7z5z6 = (HADDRI[21] ^ Dfk7z6[21]);
assign U6z5z6 = (~(S7z5z6 & Gyenv6));
assign S7z5z6 = (HADDRI[20] ^ Dfk7z6[20]);
assign E6z5z6 = (A8z5z6 & I8z5z6);
assign I8z5z6 = (~(Q8z5z6 & Q4env6));
assign Q8z5z6 = (HADDRI[19] ^ Dfk7z6[19]);
assign A8z5z6 = (~(Y8z5z6 & Ecenv6));
assign Y8z5z6 = (HADDRI[18] ^ Dfk7z6[18]);
assign O5z5z6 = (G9z5z6 & O9z5z6);
assign G9z5z6 = (W9z5z6 & Eaz5z6);
assign Eaz5z6 = (~(Maz5z6 & Sjenv6));
assign Maz5z6 = (HADDRI[17] ^ Dfk7z6[17]);
assign W9z5z6 = (~(Uaz5z6 & Dmenv6));
assign Uaz5z6 = (HADDRI[16] ^ Dfk7z6[16]);
assign Iky5z6 = (~(Cbz5z6 & Kbz5z6));
assign Kbz5z6 = (Sbz5z6 & Acz5z6);
assign Acz5z6 = (Icz5z6 & Qcz5z6);
assign Qcz5z6 = (~(Junyx6 & P6l7z6[21]));
assign Icz5z6 = (Ycz5z6 & Gdz5z6);
assign Gdz5z6 = (~(Ltnyx6 & Zlk7z6[21]));
assign Ycz5z6 = (~(Nsnyx6 & Hwk7z6[21]));
assign Sbz5z6 = (Odz5z6 & Wdz5z6);
assign Wdz5z6 = (~(Runyx6 & Xgl7z6[21]));
assign Odz5z6 = (~(Fwnyx6 & Frl7z6[21]));
assign Cbz5z6 = (Eez5z6 & Mez5z6);
assign Mez5z6 = (Uez5z6 & Cfz5z6);
assign Cfz5z6 = (~(Nwnyx6 & N1m7z6[21]));
assign Uez5z6 = (~(Lxnyx6 & Rbk7z6[21]));
assign Eez5z6 = (Kfz5z6 & Sfz5z6);
assign Sfz5z6 = (~(Txnyx6 & Vbm7z6[21]));
assign Kfz5z6 = (Qgz5z6 ? Igz5z6 : Agz5z6);
assign Qgz5z6 = (Ygz5z6 & Ghz5z6);
assign Ghz5z6 = (Ohz5z6 & Whz5z6);
assign Whz5z6 = (Eiz5z6 & Miz5z6);
assign Miz5z6 = (~(Nwnyx6 & N1m7z6[20]));
assign Eiz5z6 = (~(Lxnyx6 & Rbk7z6[20]));
assign Ohz5z6 = (Uiz5z6 & Cjz5z6);
assign Cjz5z6 = (~(Junyx6 & P6l7z6[20]));
assign Uiz5z6 = (~(Nsnyx6 & Hwk7z6[20]));
assign Ygz5z6 = (Kjz5z6 & Sjz5z6);
assign Sjz5z6 = (Akz5z6 & Ikz5z6);
assign Ikz5z6 = (~(Fwnyx6 & Frl7z6[20]));
assign Akz5z6 = (~(Ltnyx6 & Zlk7z6[20]));
assign Kjz5z6 = (Qkz5z6 & Ykz5z6);
assign Ykz5z6 = (~(Txnyx6 & Vbm7z6[20]));
assign Qkz5z6 = (~(Runyx6 & Xgl7z6[20]));
assign Igz5z6 = (Glz5z6 & Olz5z6);
assign Olz5z6 = (Wlz5z6 & Emz5z6);
assign Emz5z6 = (Mmz5z6 & Umz5z6);
assign Umz5z6 = (~(Ltnyx6 & Zlk7z6[22]));
assign Ltnyx6 = (Cnz5z6 & Knz5z6);
assign Cnz5z6 = (Snz5z6 & Aoz5z6);
assign Mmz5z6 = (~(Nsnyx6 & Hwk7z6[22]));
assign Nsnyx6 = (~(Ioz5z6 | Qoz5z6));
assign Wlz5z6 = (Yoz5z6 & Gpz5z6);
assign Gpz5z6 = (~(Junyx6 & P6l7z6[22]));
assign Junyx6 = (~(Opz5z6 | Ioz5z6));
assign Ioz5z6 = (~(Snz5z6 & Wpz5z6));
assign Yoz5z6 = (~(Runyx6 & Xgl7z6[22]));
assign Runyx6 = (Eqz5z6 & Mqz5z6);
assign Eqz5z6 = (~(Uqz5z6 | Crz5z6));
assign Glz5z6 = (Krz5z6 & Srz5z6);
assign Srz5z6 = (Asz5z6 & Isz5z6);
assign Isz5z6 = (~(Fwnyx6 & Frl7z6[22]));
assign Fwnyx6 = (Crz5z6 & Qsz5z6);
assign Asz5z6 = (~(Nwnyx6 & N1m7z6[22]));
assign Nwnyx6 = (~(Txnyx6 | Qsz5z6));
assign Krz5z6 = (Ysz5z6 & Gtz5z6);
assign Gtz5z6 = (~(Lxnyx6 & Rbk7z6[22]));
assign Lxnyx6 = (Otz5z6 & Snz5z6);
assign Snz5z6 = (Wtz5z6 & Qsz5z6);
assign Qsz5z6 = (!Uqz5z6);
assign Uqz5z6 = (~(Euz5z6 & Muz5z6));
assign Muz5z6 = (!Txnyx6);
assign Euz5z6 = (~(Uuz5z6 & Cvz5z6));
assign Cvz5z6 = (Kvz5z6 & Svz5z6);
assign Svz5z6 = (Awz5z6 & Iwz5z6);
assign Iwz5z6 = (Qwz5z6 & Ywz5z6);
assign Ywz5z6 = (~(Cslet6 | Gxz5z6));
assign Gxz5z6 = (Oxz5z6 & Xk5nv6);
assign Oxz5z6 = (Az3nv6 ^ Wxz5z6);
assign Qwz5z6 = (Eyz5z6 & Myz5z6);
assign Myz5z6 = (~(Uyz5z6 & C65nv6));
assign Uyz5z6 = (Usbiw6 ^ HADDRI[7]);
assign Eyz5z6 = (~(Qd5nv6 & Czz5z6));
assign Czz5z6 = (Hpbiw6 ^ HADDRI[6]);
assign Awz5z6 = (Kzz5z6 & Szz5z6);
assign Szz5z6 = (A006z6 & I006z6);
assign I006z6 = (~(Q006z6 & Iu5nv6));
assign Q006z6 = (Ndciw6 ^ HADDRI[15]);
assign A006z6 = (~(Y006z6 & Sz5nv6));
assign Y006z6 = (Cbciw6 ^ HADDRI[14]);
assign Kzz5z6 = (G106z6 & O106z6);
assign O106z6 = (~(W106z6 & V55nv6));
assign W106z6 = (M9ciw6 ^ HADDRI[13]);
assign G106z6 = (~(E206z6 & Jd5nv6));
assign E206z6 = (P7ciw6 ^ HADDRI[12]);
assign Kvz5z6 = (M206z6 & U206z6);
assign U206z6 = (C306z6 & K306z6);
assign K306z6 = (S306z6 & A406z6);
assign A406z6 = (~(I406z6 & El5nv6));
assign I406z6 = (Q4ciw6 ^ HADDRI[11]);
assign S306z6 = (~(Q406z6 & Aq5nv6));
assign Q406z6 = (W0ciw6 ^ HADDRI[10]);
assign C306z6 = (Y406z6 & G506z6);
assign G506z6 = (~(O506z6 & W506z6));
assign O506z6 = (Gzbiw6 ^ HADDRI[9]);
assign Y406z6 = (~(E606z6 & Qk5nv6));
assign E606z6 = (M606z6 ^ U606z6);
assign M206z6 = (C706z6 & K706z6);
assign K706z6 = (~(S706z6 & Dh5nv6));
assign S706z6 = (Bkfnv6 ^ Z4diw6);
assign C706z6 = (A806z6 & I806z6);
assign I806z6 = (~(Q806z6 & B25nv6));
assign Q806z6 = (K787z6 ^ Eg3nv6);
assign A806z6 = (~(Y806z6 & P95nv6));
assign Y806z6 = (P6diw6 ^ Ujfnv6);
assign P6diw6 = (!G987z6);
assign Uuz5z6 = (G906z6 & O906z6);
assign O906z6 = (W906z6 & Ea06z6);
assign Ea06z6 = (Ma06z6 & Ua06z6);
assign Ua06z6 = (Cb06z6 & Kb06z6);
assign Kb06z6 = (~(Sb06z6 & Ac06z6));
assign Sb06z6 = (J3diw6 ^ HADDRI[28]);
assign Cb06z6 = (~(Ic06z6 & Fw5nv6));
assign Ic06z6 = (F1diw6 ^ HADDRI[27]);
assign Ma06z6 = (Qc06z6 & Yc06z6);
assign Yc06z6 = (~(Gd06z6 & M36nv6));
assign Gd06z6 = (Pzciw6 ^ HADDRI[26]);
assign Pzciw6 = (!A887z6);
assign Qc06z6 = (~(Od06z6 & Y35nv6));
assign Od06z6 = (Gyciw6 ^ HADDRI[25]);
assign Gyciw6 = (!S787z6);
assign W906z6 = (Wd06z6 & Ee06z6);
assign Ee06z6 = (~(Me06z6 & Ko5nv6));
assign Me06z6 = (Lqciw6 ^ HADDRI[22]);
assign Wd06z6 = (Ue06z6 & Cf06z6);
assign Cf06z6 = (~(Kf06z6 & Mb5nv6));
assign Kf06z6 = (Rqmyx6 ^ Sf06z6);
assign Ue06z6 = (~(Ag06z6 & Aj5nv6));
assign Ag06z6 = (Isciw6 ^ HADDRI[23]);
assign Isciw6 = (!Gl77z6);
assign G906z6 = (Ig06z6 & Qg06z6);
assign Qg06z6 = (Yg06z6 & Gh06z6);
assign Gh06z6 = (Oh06z6 & Wh06z6);
assign Wh06z6 = (~(Ei06z6 & Bu5nv6));
assign Ei06z6 = (Oociw6 ^ HADDRI[21]);
assign Oociw6 = (!U687z6);
assign Oh06z6 = (~(Mi06z6 & I16nv6));
assign Mi06z6 = (Kmciw6 ^ HADDRI[20]);
assign Kmciw6 = (!O587z6);
assign Yg06z6 = (Ui06z6 & Cj06z6);
assign Cj06z6 = (~(Kj06z6 & E75nv6));
assign Kj06z6 = (Ukciw6 ^ HADDRI[19]);
assign Ui06z6 = (~(Sj06z6 & Se5nv6));
assign Sj06z6 = (Ejciw6 ^ HADDRI[18]);
assign Ig06z6 = (Ak06z6 & Ik06z6);
assign Ak06z6 = (Qk06z6 & Yk06z6);
assign Yk06z6 = (~(Gl06z6 & Gm5nv6));
assign Gl06z6 = (Ohciw6 ^ HADDRI[17]);
assign Ohciw6 = (!M687z6);
assign Qk06z6 = (~(Ol06z6 & Ro5nv6));
assign Ol06z6 = (Wl06z6 ^ Em06z6);
assign Wtz5z6 = (~(Crz5z6 | Mqz5z6));
assign Mqz5z6 = (Mm06z6 & Um06z6);
assign Um06z6 = (Cn06z6 & Kn06z6);
assign Kn06z6 = (Sn06z6 & Ao06z6);
assign Ao06z6 = (Io06z6 & Qo06z6);
assign Qo06z6 = (~(C8ket6 | Yo06z6));
assign Yo06z6 = (Gp06z6 & Pk8nv6);
assign Gp06z6 = (Az3nv6 ^ Op06z6);
assign Io06z6 = (Wp06z6 & Eq06z6);
assign Eq06z6 = (~(Mq06z6 & U58nv6));
assign Mq06z6 = (Kj3nv6 ^ Uq06z6);
assign Kj3nv6 = (!HADDRI[7]);
assign Wp06z6 = (~(Cr06z6 & Id8nv6));
assign Cr06z6 = (Yq3nv6 ^ Kr06z6);
assign Yq3nv6 = (!HADDRI[6]);
assign Sn06z6 = (Sr06z6 & As06z6);
assign As06z6 = (Is06z6 & Qs06z6);
assign Qs06z6 = (~(Ys06z6 & Tt8nv6));
assign Ys06z6 = (Gt06z6 ^ Ot06z6);
assign Gt06z6 = (!HADDRI[15]);
assign Is06z6 = (~(Wt06z6 & Wy8nv6));
assign Wt06z6 = (Eu06z6 ^ Mu06z6);
assign Eu06z6 = (!HADDRI[14]);
assign Sr06z6 = (Uu06z6 & Cv06z6);
assign Cv06z6 = (~(Kv06z6 & N58nv6));
assign Kv06z6 = (Sv06z6 ^ Aw06z6);
assign Sv06z6 = (!HADDRI[13]);
assign Uu06z6 = (~(Iw06z6 & Bd8nv6));
assign Iw06z6 = (Qw06z6 ^ Yw06z6);
assign Qw06z6 = (!HADDRI[12]);
assign Cn06z6 = (Gx06z6 & Ox06z6);
assign Ox06z6 = (Wx06z6 & Ey06z6);
assign Ey06z6 = (My06z6 & Uy06z6);
assign Uy06z6 = (~(Cz06z6 & Wk8nv6));
assign Cz06z6 = (Kz06z6 ^ Sz06z6);
assign Kz06z6 = (!HADDRI[11]);
assign My06z6 = (~(A016z6 & Lp8nv6));
assign A016z6 = (I016z6 ^ Q016z6);
assign I016z6 = (!HADDRI[10]);
assign Wx06z6 = (Y016z6 & G116z6);
assign G116z6 = (~(O116z6 & W116z6));
assign O116z6 = (E216z6 ^ M216z6);
assign E216z6 = (!HADDRI[9]);
assign Y016z6 = (~(U216z6 & Ik8nv6));
assign U216z6 = (M606z6 ^ C316z6);
assign Gx06z6 = (K316z6 & S316z6);
assign S316z6 = (~(A416z6 & Vg8nv6));
assign A416z6 = (I416z6 ^ Bw3nv6);
assign K316z6 = (Q416z6 & Y416z6);
assign Y416z6 = (~(G516z6 & T18nv6));
assign G516z6 = (Eg3nv6 ^ O516z6);
assign Q416z6 = (~(W516z6 & H98nv6));
assign W516z6 = (Zn3nv6 ^ E616z6);
assign Mm06z6 = (M616z6 & U616z6);
assign U616z6 = (C716z6 & K716z6);
assign K716z6 = (S716z6 & A816z6);
assign A816z6 = (I816z6 & Q816z6);
assign Q816z6 = (~(Y816z6 & G916z6));
assign Y816z6 = (Tpmyx6 ^ O916z6);
assign Tpmyx6 = (!HADDRI[28]);
assign I816z6 = (~(W916z6 & Jv8nv6));
assign W916z6 = (Vsmyx6 ^ Ea16z6);
assign Vsmyx6 = (!HADDRI[27]);
assign S716z6 = (Ma16z6 & Ua16z6);
assign Ua16z6 = (~(Cb16z6 & Q29nv6));
assign Cb16z6 = (Dtmyx6 ^ Kb16z6);
assign Dtmyx6 = (!HADDRI[26]);
assign Ma16z6 = (~(Sb16z6 & Q38nv6));
assign Sb16z6 = (Bqmyx6 ^ Ac16z6);
assign C716z6 = (Ic16z6 & Qc16z6);
assign Qc16z6 = (~(Yc16z6 & Co8nv6));
assign Yc16z6 = (Jqmyx6 ^ Gd16z6);
assign Jqmyx6 = (!HADDRI[22]);
assign Ic16z6 = (Od16z6 & Wd16z6);
assign Wd16z6 = (~(Ee16z6 & Eb8nv6));
assign Ee16z6 = (Rqmyx6 ^ Me16z6);
assign Od16z6 = (~(Ue16z6 & Si8nv6));
assign Ue16z6 = (Fsmyx6 ^ Cf16z6);
assign Fsmyx6 = (!HADDRI[23]);
assign M616z6 = (Kf16z6 & Sf16z6);
assign Sf16z6 = (Ag16z6 & Ig16z6);
assign Ig16z6 = (Qg16z6 & Yg16z6);
assign Yg16z6 = (~(Gh16z6 & Mt8nv6));
assign Gh16z6 = (Zqmyx6 ^ Oh16z6);
assign Zqmyx6 = (!HADDRI[21]);
assign Qg16z6 = (~(Wh16z6 & M09nv6));
assign Wh16z6 = (Nsmyx6 ^ Ei16z6);
assign Nsmyx6 = (!HADDRI[20]);
assign Ag16z6 = (Mi16z6 & Ui16z6);
assign Ui16z6 = (~(Cj16z6 & W68nv6));
assign Cj16z6 = (Kj16z6 ^ Sj16z6);
assign Kj16z6 = (!HADDRI[19]);
assign Mi16z6 = (~(Ak16z6 & Ke8nv6));
assign Ak16z6 = (Ik16z6 ^ Qk16z6);
assign Ik16z6 = (!HADDRI[18]);
assign Kf16z6 = (Yk16z6 & Gl16z6);
assign Yk16z6 = (Ol16z6 & Wl16z6);
assign Wl16z6 = (~(Em16z6 & Yl8nv6));
assign Em16z6 = (Mm16z6 ^ Um16z6);
assign Mm16z6 = (!HADDRI[17]);
assign Ol16z6 = (~(Cn16z6 & Jo8nv6));
assign Cn16z6 = (Wl06z6 ^ Kn16z6);
assign Crz5z6 = (Sn16z6 & Ao16z6);
assign Ao16z6 = (Io16z6 & Qo16z6);
assign Qo16z6 = (Yo16z6 & Gp16z6);
assign Gp16z6 = (Op16z6 & Wp16z6);
assign Wp16z6 = (~(C0let6 | Eq16z6));
assign Eq16z6 = (Mq16z6 & T27nv6);
assign Mq16z6 = (Az3nv6 ^ Uq16z6);
assign Op16z6 = (Cr16z6 & Kr16z6);
assign Kr16z6 = (~(Sr16z6 & Yn6nv6));
assign Sr16z6 = (Gsbiw6 ^ HADDRI[7]);
assign Cr16z6 = (~(Mv6nv6 & As16z6));
assign As16z6 = (Apbiw6 ^ HADDRI[6]);
assign Yo16z6 = (Is16z6 & Qs16z6);
assign Qs16z6 = (Ys16z6 & Gt16z6);
assign Gt16z6 = (~(Ot16z6 & Xb7nv6));
assign Ot16z6 = (Zcciw6 ^ HADDRI[15]);
assign Ys16z6 = (~(Wt16z6 & Ah7nv6));
assign Wt16z6 = (Vaciw6 ^ HADDRI[14]);
assign Is16z6 = (Eu16z6 & Mu16z6);
assign Mu16z6 = (~(Uu16z6 & Rn6nv6));
assign Uu16z6 = (F9ciw6 ^ HADDRI[13]);
assign Eu16z6 = (~(Cv16z6 & Fv6nv6));
assign Cv16z6 = (I7ciw6 ^ HADDRI[12]);
assign Io16z6 = (Kv16z6 & Sv16z6);
assign Sv16z6 = (Aw16z6 & Iw16z6);
assign Iw16z6 = (Qw16z6 & Yw16z6);
assign Yw16z6 = (~(Gx16z6 & A37nv6));
assign Gx16z6 = (V3ciw6 ^ HADDRI[11]);
assign Qw16z6 = (~(Ox16z6 & P77nv6));
assign Ox16z6 = (P0ciw6 ^ HADDRI[10]);
assign Aw16z6 = (Wx16z6 & Ey16z6);
assign Ey16z6 = (~(My16z6 & Uy16z6));
assign My16z6 = (Zybiw6 ^ HADDRI[9]);
assign Wx16z6 = (~(Cz16z6 & M27nv6));
assign Cz16z6 = (M606z6 ^ Kz16z6);
assign Kv16z6 = (Sz16z6 & A026z6);
assign A026z6 = (~(I026z6 & Zy6nv6));
assign I026z6 = (Bkfnv6 ^ S4diw6);
assign Sz16z6 = (Q026z6 & Y026z6);
assign Y026z6 = (~(G126z6 & Xj6nv6));
assign G126z6 = (Ee87z6 ^ Eg3nv6);
assign Q026z6 = (~(O126z6 & Lr6nv6));
assign O126z6 = (I6diw6 ^ Ujfnv6);
assign I6diw6 = (!Ag87z6);
assign Sn16z6 = (W126z6 & E226z6);
assign E226z6 = (M226z6 & U226z6);
assign U226z6 = (C326z6 & K326z6);
assign K326z6 = (S326z6 & A426z6);
assign A426z6 = (~(I426z6 & Q426z6));
assign I426z6 = (V2diw6 ^ HADDRI[28]);
assign S326z6 = (~(Y426z6 & Nd7nv6));
assign Y426z6 = (Y0diw6 ^ HADDRI[27]);
assign C326z6 = (G526z6 & O526z6);
assign O526z6 = (~(W526z6 & Bl7nv6));
assign W526z6 = (Izciw6 ^ HADDRI[26]);
assign Izciw6 = (!Ue87z6);
assign G526z6 = (~(E626z6 & Ul6nv6));
assign E626z6 = (Zxciw6 ^ HADDRI[25]);
assign Zxciw6 = (!Me87z6);
assign M226z6 = (M626z6 & U626z6);
assign U626z6 = (~(C726z6 & G67nv6));
assign C726z6 = (Eqciw6 ^ HADDRI[22]);
assign M626z6 = (K726z6 & S726z6);
assign S726z6 = (~(A826z6 & It6nv6));
assign A826z6 = (Rqmyx6 ^ I826z6);
assign K726z6 = (~(Q826z6 & W07nv6));
assign Q826z6 = (Bsciw6 ^ HADDRI[23]);
assign Bsciw6 = (!Ol77z6);
assign W126z6 = (Y826z6 & G926z6);
assign G926z6 = (O926z6 & W926z6);
assign W926z6 = (Ea26z6 & Ma26z6);
assign Ma26z6 = (~(Ua26z6 & Qb7nv6));
assign Ua26z6 = (Aociw6 ^ HADDRI[21]);
assign Aociw6 = (!Od87z6);
assign Ea26z6 = (~(Cb26z6 & Ej7nv6));
assign Cb26z6 = (Dmciw6 ^ HADDRI[20]);
assign Dmciw6 = (!Ic87z6);
assign O926z6 = (Kb26z6 & Sb26z6);
assign Sb26z6 = (~(Ac26z6 & Ap6nv6));
assign Ac26z6 = (Nkciw6 ^ HADDRI[19]);
assign Kb26z6 = (~(Ic26z6 & Ow6nv6));
assign Ic26z6 = (Xiciw6 ^ HADDRI[18]);
assign Y826z6 = (Qc26z6 & Yc26z6);
assign Qc26z6 = (Gd26z6 & Od26z6);
assign Od26z6 = (~(Wd26z6 & C47nv6));
assign Wd26z6 = (Hhciw6 ^ HADDRI[17]);
assign Hhciw6 = (!Gd87z6);
assign Gd26z6 = (~(Ee26z6 & N67nv6));
assign Ee26z6 = (Wl06z6 ^ Me26z6);
assign Otz5z6 = (~(Wpz5z6 | Knz5z6));
assign Knz5z6 = (Ue26z6 & Cf26z6);
assign Cf26z6 = (Kf26z6 & Sf26z6);
assign Sf26z6 = (Ag26z6 & Ig26z6);
assign Ig26z6 = (Qg26z6 & Yg26z6);
assign Yg26z6 = (~(Cwhet6 | Gh26z6));
assign Gh26z6 = (Oh26z6 & U0dnv6);
assign Oh26z6 = (Az3nv6 ^ Wh26z6);
assign Qg26z6 = (Ei26z6 & Mi26z6);
assign Mi26z6 = (~(Ui26z6 & Zlcnv6));
assign Ui26z6 = (Jqbiw6 ^ HADDRI[7]);
assign Ei26z6 = (~(Ntcnv6 & Cj26z6));
assign Cj26z6 = (Fobiw6 ^ HADDRI[6]);
assign Ag26z6 = (Kj26z6 & Sj26z6);
assign Sj26z6 = (Ak26z6 & Ik26z6);
assign Ik26z6 = (~(Qk26z6 & Y9dnv6));
assign Qk26z6 = (Xbciw6 ^ HADDRI[15]);
assign Ak26z6 = (~(Yk26z6 & Bfdnv6));
assign Yk26z6 = (Aaciw6 ^ HADDRI[14]);
assign Kj26z6 = (Gl26z6 & Ol26z6);
assign Ol26z6 = (~(Wl26z6 & Slcnv6));
assign Wl26z6 = (K8ciw6 ^ HADDRI[13]);
assign Gl26z6 = (~(Em26z6 & Gtcnv6));
assign Em26z6 = (L5ciw6 ^ HADDRI[12]);
assign Kf26z6 = (Mm26z6 & Um26z6);
assign Um26z6 = (Cn26z6 & Kn26z6);
assign Kn26z6 = (Sn26z6 & Ao26z6);
assign Ao26z6 = (~(Io26z6 & B1dnv6));
assign Io26z6 = (Y1ciw6 ^ HADDRI[11]);
assign Sn26z6 = (~(Qo26z6 & Q5dnv6));
assign Qo26z6 = (Uzbiw6 ^ HADDRI[10]);
assign Cn26z6 = (Yo26z6 & Gp26z6);
assign Gp26z6 = (~(Op26z6 & Wp26z6));
assign Op26z6 = (Eybiw6 ^ HADDRI[9]);
assign Yo26z6 = (~(Eq26z6 & N0dnv6));
assign Eq26z6 = (M606z6 ^ Mq26z6);
assign Mm26z6 = (Uq26z6 & Cr26z6);
assign Cr26z6 = (~(Kr26z6 & Axcnv6));
assign Kr26z6 = (Bkfnv6 ^ X3diw6);
assign Uq26z6 = (Sr26z6 & As26z6);
assign As26z6 = (~(Is26z6 & Yhcnv6));
assign Is26z6 = (Yk87z6 ^ Eg3nv6);
assign Sr26z6 = (~(Qs26z6 & Mpcnv6));
assign Qs26z6 = (N5diw6 ^ Ujfnv6);
assign N5diw6 = (!Um87z6);
assign Ue26z6 = (Ys26z6 & Gt26z6);
assign Gt26z6 = (Ot26z6 & Wt26z6);
assign Wt26z6 = (Eu26z6 & Mu26z6);
assign Mu26z6 = (Uu26z6 & Cv26z6);
assign Cv26z6 = (~(Kv26z6 & Sv26z6));
assign Kv26z6 = (A2diw6 ^ HADDRI[28]);
assign Uu26z6 = (~(Aw26z6 & Obdnv6));
assign Aw26z6 = (D0diw6 ^ HADDRI[27]);
assign Eu26z6 = (Iw26z6 & Qw26z6);
assign Qw26z6 = (~(Yw26z6 & Vidnv6));
assign Yw26z6 = (Nyciw6 ^ HADDRI[26]);
assign Nyciw6 = (!Ol87z6);
assign Iw26z6 = (~(Gx26z6 & Vjcnv6));
assign Gx26z6 = (Exciw6 ^ HADDRI[25]);
assign Exciw6 = (!Gl87z6);
assign Ot26z6 = (Ox26z6 & Wx26z6);
assign Wx26z6 = (~(Ey26z6 & H4dnv6));
assign Ey26z6 = (Jpciw6 ^ HADDRI[22]);
assign Ox26z6 = (My26z6 & Uy26z6);
assign Uy26z6 = (~(Cz26z6 & Jrcnv6));
assign Cz26z6 = (Rqmyx6 ^ Kz26z6);
assign My26z6 = (~(Sz26z6 & Xycnv6));
assign Sz26z6 = (Grciw6 ^ HADDRI[23]);
assign Grciw6 = (!Mm77z6);
assign Ys26z6 = (A036z6 & I036z6);
assign I036z6 = (Q036z6 & Y036z6);
assign Y036z6 = (G136z6 & O136z6);
assign O136z6 = (~(W136z6 & R9dnv6));
assign W136z6 = (Fnciw6 ^ HADDRI[21]);
assign Fnciw6 = (!Ik87z6);
assign G136z6 = (~(E236z6 & Rgdnv6));
assign E236z6 = (Ilciw6 ^ HADDRI[20]);
assign Ilciw6 = (!Cj87z6);
assign Q036z6 = (M236z6 & U236z6);
assign U236z6 = (~(C336z6 & Bncnv6));
assign C336z6 = (Sjciw6 ^ HADDRI[19]);
assign M236z6 = (~(K336z6 & Pucnv6));
assign K336z6 = (Ciciw6 ^ HADDRI[18]);
assign A036z6 = (S336z6 & A436z6);
assign S336z6 = (I436z6 & Q436z6);
assign Q436z6 = (~(Y436z6 & D2dnv6));
assign Y436z6 = (Mgciw6 ^ HADDRI[17]);
assign Mgciw6 = (!Ak87z6);
assign I436z6 = (~(G536z6 & O4dnv6));
assign G536z6 = (Wl06z6 ^ O536z6);
assign Wpz5z6 = (!Aoz5z6);
assign Aoz5z6 = (~(W536z6 | Qoz5z6));
assign Qoz5z6 = (!Opz5z6);
assign Opz5z6 = (~(E636z6 & M636z6));
assign M636z6 = (U636z6 & C736z6);
assign C736z6 = (K736z6 & S736z6);
assign S736z6 = (A836z6 & I836z6);
assign I836z6 = (~(Cgjet6 | Q836z6));
assign Q836z6 = (Y836z6 & X1anv6);
assign Y836z6 = (Az3nv6 ^ G936z6);
assign A836z6 = (O936z6 & W936z6);
assign W936z6 = (~(Ea36z6 & Cn9nv6));
assign Ea36z6 = (Lrbiw6 ^ HADDRI[7]);
assign O936z6 = (~(Qu9nv6 & Ma36z6));
assign Ma36z6 = (Tobiw6 ^ HADDRI[6]);
assign K736z6 = (Ua36z6 & Cb36z6);
assign Cb36z6 = (Kb36z6 & Sb36z6);
assign Sb36z6 = (~(Ac36z6 & Bbanv6));
assign Ac36z6 = (Lcciw6 ^ HADDRI[15]);
assign Kb36z6 = (~(Ic36z6 & Eganv6));
assign Ic36z6 = (Oaciw6 ^ HADDRI[14]);
assign Ua36z6 = (Qc36z6 & Yc36z6);
assign Yc36z6 = (~(Gd36z6 & Vm9nv6));
assign Gd36z6 = (Y8ciw6 ^ HADDRI[13]);
assign Qc36z6 = (~(Od36z6 & Ju9nv6));
assign Od36z6 = (N6ciw6 ^ HADDRI[12]);
assign U636z6 = (Wd36z6 & Ee36z6);
assign Ee36z6 = (Me36z6 & Ue36z6);
assign Ue36z6 = (Cf36z6 & Kf36z6);
assign Kf36z6 = (~(Sf36z6 & E2anv6));
assign Sf36z6 = (A3ciw6 ^ HADDRI[11]);
assign Cf36z6 = (~(Ag36z6 & T6anv6));
assign Ag36z6 = (I0ciw6 ^ HADDRI[10]);
assign Me36z6 = (Ig36z6 & Qg36z6);
assign Qg36z6 = (~(Yg36z6 & Gh36z6));
assign Yg36z6 = (Sybiw6 ^ HADDRI[9]);
assign Ig36z6 = (~(Oh36z6 & Q1anv6));
assign Oh36z6 = (HADDRI[8] ^ Bal7z6[8]);
assign Wd36z6 = (Wh36z6 & Ei36z6);
assign Ei36z6 = (~(Mi36z6 & Dy9nv6));
assign Mi36z6 = (Bkfnv6 ^ L4diw6);
assign Wh36z6 = (Ui36z6 & Cj36z6);
assign Cj36z6 = (~(Kj36z6 & Bj9nv6));
assign Kj36z6 = (Jadiw6 ^ Njfnv6);
assign Jadiw6 = (!My87z6);
assign Ui36z6 = (~(Sj36z6 & Pq9nv6));
assign Sj36z6 = (B6diw6 ^ Ujfnv6);
assign B6diw6 = (!I097z6);
assign E636z6 = (Ak36z6 & Ik36z6);
assign Ik36z6 = (Qk36z6 & Yk36z6);
assign Yk36z6 = (Gl36z6 & Ol36z6);
assign Ol36z6 = (Wl36z6 & Em36z6);
assign Em36z6 = (~(Mm36z6 & Um36z6));
assign Mm36z6 = (O2diw6 ^ HADDRI[28]);
assign Wl36z6 = (~(Cn36z6 & Rcanv6));
assign Cn36z6 = (R0diw6 ^ HADDRI[27]);
assign Gl36z6 = (Kn36z6 & Sn36z6);
assign Sn36z6 = (~(Ao36z6 & Yjanv6));
assign Ao36z6 = (Bzciw6 ^ HADDRI[26]);
assign Bzciw6 = (!Cz87z6);
assign Kn36z6 = (~(Io36z6 & Yk9nv6));
assign Io36z6 = (Sxciw6 ^ HADDRI[25]);
assign Sxciw6 = (!Uy87z6);
assign Qk36z6 = (Qo36z6 & Yo36z6);
assign Yo36z6 = (~(Gp36z6 & K5anv6));
assign Gp36z6 = (Xpciw6 ^ HADDRI[22]);
assign Qo36z6 = (Op36z6 & Wp36z6);
assign Wp36z6 = (~(Eq36z6 & Ms9nv6));
assign Eq36z6 = (HADDRI[24] ^ Bal7z6[24]);
assign Op36z6 = (~(Mq36z6 & A0anv6));
assign Mq36z6 = (Urciw6 ^ HADDRI[23]);
assign Urciw6 = (!Wl77z6);
assign Ak36z6 = (Uq36z6 & Cr36z6);
assign Cr36z6 = (Kr36z6 & Sr36z6);
assign Sr36z6 = (As36z6 & Is36z6);
assign Is36z6 = (~(Qs36z6 & Uaanv6));
assign Qs36z6 = (Tnciw6 ^ HADDRI[21]);
assign Tnciw6 = (!Wx87z6);
assign As36z6 = (~(Ys36z6 & Uhanv6));
assign Ys36z6 = (Wlciw6 ^ HADDRI[20]);
assign Wlciw6 = (!Qw87z6);
assign Kr36z6 = (Gt36z6 & Ot36z6);
assign Ot36z6 = (~(Wt36z6 & Eo9nv6));
assign Wt36z6 = (Gkciw6 ^ HADDRI[19]);
assign Gt36z6 = (~(Eu36z6 & Sv9nv6));
assign Eu36z6 = (Qiciw6 ^ HADDRI[18]);
assign Uq36z6 = (Mu36z6 & Uu36z6);
assign Mu36z6 = (Cv36z6 & Kv36z6);
assign Kv36z6 = (~(Sv36z6 & G3anv6));
assign Sv36z6 = (Ahciw6 ^ HADDRI[17]);
assign Ahciw6 = (!Ox87z6);
assign Cv36z6 = (~(Aw36z6 & R5anv6));
assign Aw36z6 = (HADDRI[16] ^ Bal7z6[16]);
assign W536z6 = (Iw36z6 & Qw36z6);
assign Qw36z6 = (Yw36z6 & Gx36z6);
assign Gx36z6 = (Ox36z6 & Wx36z6);
assign Wx36z6 = (Ey36z6 & My36z6);
assign My36z6 = (~(Coiet6 | Uy36z6));
assign Uy36z6 = (Cz36z6 & Mjbnv6);
assign Cz36z6 = (Az3nv6 ^ Kz36z6);
assign Ey36z6 = (Sz36z6 & A046z6);
assign A046z6 = (~(I046z6 & R4bnv6));
assign I046z6 = (Xqbiw6 ^ HADDRI[7]);
assign Sz36z6 = (~(Fcbnv6 & Q046z6));
assign Q046z6 = (Mobiw6 ^ HADDRI[6]);
assign Ox36z6 = (Y046z6 & G146z6);
assign G146z6 = (O146z6 & W146z6);
assign W146z6 = (~(E246z6 & Qsbnv6));
assign E246z6 = (Ecciw6 ^ HADDRI[15]);
assign O146z6 = (~(M246z6 & Txbnv6));
assign M246z6 = (Haciw6 ^ HADDRI[14]);
assign Y046z6 = (U246z6 & C346z6);
assign C346z6 = (~(K346z6 & K4bnv6));
assign K346z6 = (R8ciw6 ^ HADDRI[13]);
assign U246z6 = (~(S346z6 & Ybbnv6));
assign S346z6 = (Z5ciw6 ^ HADDRI[12]);
assign Yw36z6 = (A446z6 & I446z6);
assign I446z6 = (Q446z6 & Y446z6);
assign Y446z6 = (G546z6 & O546z6);
assign O546z6 = (~(W546z6 & Tjbnv6));
assign W546z6 = (M2ciw6 ^ HADDRI[11]);
assign G546z6 = (~(E646z6 & Iobnv6));
assign E646z6 = (B0ciw6 ^ HADDRI[10]);
assign Q446z6 = (M646z6 & U646z6);
assign U646z6 = (~(C746z6 & K746z6));
assign C746z6 = (Lybiw6 ^ HADDRI[9]);
assign M646z6 = (~(S746z6 & Fjbnv6));
assign S746z6 = (M606z6 ^ A846z6);
assign A446z6 = (I846z6 & Q846z6);
assign Q846z6 = (~(Y846z6 & Sfbnv6));
assign Y846z6 = (Bkfnv6 ^ E4diw6);
assign I846z6 = (G946z6 & O946z6);
assign O946z6 = (~(W946z6 & Q0bnv6));
assign W946z6 = (Sr87z6 ^ Eg3nv6);
assign G946z6 = (~(Ea46z6 & E8bnv6));
assign Ea46z6 = (U5diw6 ^ Ujfnv6);
assign U5diw6 = (!Ot87z6);
assign Iw36z6 = (Ma46z6 & Ua46z6);
assign Ua46z6 = (Cb46z6 & Kb46z6);
assign Kb46z6 = (Sb46z6 & Ac46z6);
assign Ac46z6 = (Ic46z6 & Qc46z6);
assign Qc46z6 = (~(Yc46z6 & Gd46z6));
assign Yc46z6 = (H2diw6 ^ HADDRI[28]);
assign Ic46z6 = (~(Od46z6 & Gubnv6));
assign Od46z6 = (K0diw6 ^ HADDRI[27]);
assign Sb46z6 = (Wd46z6 & Ee46z6);
assign Ee46z6 = (~(Me46z6 & N1cnv6));
assign Me46z6 = (Uyciw6 ^ HADDRI[26]);
assign Uyciw6 = (!Is87z6);
assign Wd46z6 = (~(Ue46z6 & N2bnv6));
assign Ue46z6 = (Lxciw6 ^ HADDRI[25]);
assign Lxciw6 = (!As87z6);
assign Cb46z6 = (Cf46z6 & Kf46z6);
assign Kf46z6 = (~(Sf46z6 & Zmbnv6));
assign Sf46z6 = (Qpciw6 ^ HADDRI[22]);
assign Cf46z6 = (Ag46z6 & Ig46z6);
assign Ig46z6 = (~(Qg46z6 & Babnv6));
assign Qg46z6 = (Rqmyx6 ^ Yg46z6);
assign Rqmyx6 = (!HADDRI[24]);
assign Ag46z6 = (~(Gh46z6 & Phbnv6));
assign Gh46z6 = (Nrciw6 ^ HADDRI[23]);
assign Nrciw6 = (!Em77z6);
assign Ma46z6 = (Oh46z6 & Wh46z6);
assign Wh46z6 = (Ei46z6 & Mi46z6);
assign Mi46z6 = (Ui46z6 & Cj46z6);
assign Cj46z6 = (~(Kj46z6 & Jsbnv6));
assign Kj46z6 = (Mnciw6 ^ HADDRI[21]);
assign Mnciw6 = (!Cr87z6);
assign Ui46z6 = (~(Sj46z6 & Jzbnv6));
assign Sj46z6 = (Plciw6 ^ HADDRI[20]);
assign Plciw6 = (!Wp87z6);
assign Ei46z6 = (Ak46z6 & Ik46z6);
assign Ik46z6 = (~(Qk46z6 & T5bnv6));
assign Qk46z6 = (Zjciw6 ^ HADDRI[19]);
assign Ak46z6 = (~(Yk46z6 & Hdbnv6));
assign Yk46z6 = (Jiciw6 ^ HADDRI[18]);
assign Oh46z6 = (Gl46z6 & Ol46z6);
assign Gl46z6 = (Wl46z6 & Em46z6);
assign Em46z6 = (~(Mm46z6 & Vkbnv6));
assign Mm46z6 = (Tgciw6 ^ HADDRI[17]);
assign Tgciw6 = (!Uq87z6);
assign Wl46z6 = (~(Um46z6 & Gnbnv6));
assign Um46z6 = (Wl06z6 ^ Cn46z6);
assign Ysz5z6 = (~(Txnyx6 & Vbm7z6[22]));
assign Txnyx6 = (Kn46z6 & Sn46z6);
assign Sn46z6 = (Ao46z6 & Io46z6);
assign Io46z6 = (Qo46z6 & Yo46z6);
assign Yo46z6 = (Gp46z6 & Op46z6);
assign Op46z6 = (~(Ckmet6 | Wp46z6));
assign Wp46z6 = (Eq46z6 & Hz3nv6);
assign Eq46z6 = (Az3nv6 ^ Mq46z6);
assign Az3nv6 = (!HADDRI[5]);
assign HADDRI[5] = (Crcdt6 ? Dvc7z6[5] : X0d7z6[5]);
assign X0d7z6[5] = (~(Uq46z6 & Cr46z6));
assign Cr46z6 = (Kr46z6 & Sr46z6);
assign Sr46z6 = (~(Pic7z6[5] & Ir0ov6));
assign Kr46z6 = (As46z6 & Is46z6);
assign Is46z6 = (Qs46z6 | Ke0ov6);
assign Ke0ov6 = (Ys46z6 & Gt46z6);
assign Gt46z6 = (~(Wkd7z6[5] & Ddmhw6));
assign Ys46z6 = (Ot46z6 & Wt46z6);
assign Wt46z6 = (~(Xhd7z6[5] & Eu46z6));
assign Ot46z6 = (~(Vnd7z6[5] & Jamnv6));
assign As46z6 = (~(Pdc7z6[5] & Mu46z6));
assign Uq46z6 = (Uu46z6 & Cv46z6);
assign Cv46z6 = (~(Znnov6 & P2j7z6[3]));
assign Uu46z6 = (~(Qdcdt6 & Fhc7z6[5]));
assign Gp46z6 = (Kv46z6 & Sv46z6);
assign Sv46z6 = (~(Aw46z6 & Dj3nv6));
assign Aw46z6 = (Btbiw6 ^ HADDRI[7]);
assign HADDRI[7] = (Crcdt6 ? Dvc7z6[7] : X0d7z6[7]);
assign X0d7z6[7] = (~(Iw46z6 & Qw46z6));
assign Qw46z6 = (Yw46z6 & Gx46z6);
assign Gx46z6 = (~(Pdc7z6[7] & Mu46z6));
assign Yw46z6 = (Ox46z6 & Wx46z6);
assign Wx46z6 = (~(Znnov6 & Ey46z6));
assign Ey46z6 = (Qti7z6[7] | P2j7z6[5]);
assign Ox46z6 = (Qs46z6 | I60ov6);
assign I60ov6 = (My46z6 & Uy46z6);
assign Uy46z6 = (~(Wkd7z6[7] & Ddmhw6));
assign My46z6 = (Cz46z6 & Kz46z6);
assign Kz46z6 = (~(Xhd7z6[7] & Eu46z6));
assign Cz46z6 = (~(Vnd7z6[7] & Jamnv6));
assign Iw46z6 = (Sz46z6 & A056z6);
assign A056z6 = (~(Pic7z6[7] & Ir0ov6));
assign Sz46z6 = (~(Qdcdt6 & Fhc7z6[7]));
assign Kv46z6 = (~(Fr3nv6 & I056z6));
assign I056z6 = (Opbiw6 ^ HADDRI[6]);
assign HADDRI[6] = (Crcdt6 ? Dvc7z6[6] : X0d7z6[6]);
assign X0d7z6[6] = (~(Q056z6 & Y056z6));
assign Y056z6 = (G156z6 & O156z6);
assign O156z6 = (~(Pic7z6[6] & Ir0ov6));
assign G156z6 = (W156z6 & E256z6);
assign E256z6 = (Qs46z6 | Ja0ov6);
assign Ja0ov6 = (M256z6 & U256z6);
assign U256z6 = (~(Wkd7z6[6] & Ddmhw6));
assign M256z6 = (C356z6 & K356z6);
assign K356z6 = (~(Xhd7z6[6] & Eu46z6));
assign C356z6 = (~(Vnd7z6[6] & Jamnv6));
assign W156z6 = (~(Pdc7z6[6] & Mu46z6));
assign Q056z6 = (S356z6 & A456z6);
assign A456z6 = (~(Znnov6 & P2j7z6[4]));
assign S356z6 = (~(Qdcdt6 & Fhc7z6[6]));
assign Qo46z6 = (I456z6 & Q456z6);
assign Q456z6 = (Y456z6 & G556z6);
assign G556z6 = (~(O556z6 & Hs3nv6));
assign O556z6 = (Udciw6 ^ HADDRI[15]);
assign HADDRI[15] = (Crcdt6 ? Dvc7z6[15] : X0d7z6[15]);
assign X0d7z6[15] = (~(W556z6 & E656z6));
assign E656z6 = (M656z6 & U656z6);
assign U656z6 = (~(Pic7z6[15] & Ir0ov6));
assign M656z6 = (C756z6 & K756z6);
assign K756z6 = (Qs46z6 | Aaznv6);
assign Aaznv6 = (S756z6 & A856z6);
assign A856z6 = (~(Wkd7z6[15] & Ddmhw6));
assign S756z6 = (I856z6 & Q856z6);
assign Q856z6 = (~(Xhd7z6[15] & Eu46z6));
assign I856z6 = (~(Vnd7z6[15] & Jamnv6));
assign C756z6 = (~(Pdc7z6[15] & Mu46z6));
assign W556z6 = (Y856z6 & G956z6);
assign G956z6 = (~(Pnb7z6[15] & Znnov6));
assign Y856z6 = (~(Qdcdt6 & Fhc7z6[15]));
assign Y456z6 = (~(O956z6 & J04nv6));
assign O956z6 = (Jbciw6 ^ HADDRI[14]);
assign HADDRI[14] = (Crcdt6 ? Dvc7z6[14] : X0d7z6[14]);
assign X0d7z6[14] = (~(W956z6 & Ea56z6));
assign Ea56z6 = (Ma56z6 & Ua56z6);
assign Ua56z6 = (~(Pic7z6[14] & Ir0ov6));
assign Ma56z6 = (Cb56z6 & Kb56z6);
assign Kb56z6 = (Qs46z6 | Beznv6);
assign Beznv6 = (Sb56z6 & Ac56z6);
assign Ac56z6 = (~(Wkd7z6[14] & Ddmhw6));
assign Sb56z6 = (Ic56z6 & Qc56z6);
assign Qc56z6 = (~(Xhd7z6[14] & Eu46z6));
assign Ic56z6 = (~(Vnd7z6[14] & Jamnv6));
assign Cb56z6 = (~(Pdc7z6[14] & Mu46z6));
assign W956z6 = (Yc56z6 & Gd56z6);
assign Gd56z6 = (~(Pnb7z6[14] & Znnov6));
assign Yc56z6 = (~(Qdcdt6 & Fhc7z6[14]));
assign I456z6 = (Od56z6 & Wd56z6);
assign Wd56z6 = (~(Ee56z6 & Wi3nv6));
assign Ee56z6 = (T9ciw6 ^ HADDRI[13]);
assign HADDRI[13] = (Crcdt6 ? Dvc7z6[13] : X0d7z6[13]);
assign X0d7z6[13] = (~(Me56z6 & Ue56z6));
assign Ue56z6 = (Cf56z6 & Kf56z6);
assign Kf56z6 = (~(Pic7z6[13] & Ir0ov6));
assign Cf56z6 = (Sf56z6 & Ag56z6);
assign Ag56z6 = (Qs46z6 | Ciznv6);
assign Ciznv6 = (Ig56z6 & Qg56z6);
assign Qg56z6 = (~(Wkd7z6[13] & Ddmhw6));
assign Ig56z6 = (Yg56z6 & Gh56z6);
assign Gh56z6 = (~(Xhd7z6[13] & Eu46z6));
assign Yg56z6 = (~(Vnd7z6[13] & Jamnv6));
assign Sf56z6 = (~(Pdc7z6[13] & Mu46z6));
assign Me56z6 = (Oh56z6 & Wh56z6);
assign Wh56z6 = (~(Pnb7z6[13] & Znnov6));
assign Oh56z6 = (~(Qdcdt6 & Fhc7z6[13]));
assign Od56z6 = (~(Ei56z6 & Mr3nv6));
assign Ei56z6 = (D8ciw6 ^ HADDRI[12]);
assign HADDRI[12] = (Crcdt6 ? Dvc7z6[12] : X0d7z6[12]);
assign X0d7z6[12] = (~(Mi56z6 & Ui56z6));
assign Ui56z6 = (Cj56z6 & Kj56z6);
assign Kj56z6 = (~(Pic7z6[12] & Ir0ov6));
assign Cj56z6 = (Sj56z6 & Ak56z6);
assign Ak56z6 = (Qs46z6 | Dmznv6);
assign Dmznv6 = (Ik56z6 & Qk56z6);
assign Qk56z6 = (~(Wkd7z6[12] & Ddmhw6));
assign Ik56z6 = (Yk56z6 & Gl56z6);
assign Gl56z6 = (~(Xhd7z6[12] & Eu46z6));
assign Yk56z6 = (~(Vnd7z6[12] & Jamnv6));
assign Sj56z6 = (~(Pdc7z6[12] & Mu46z6));
assign Mi56z6 = (Ol56z6 & Wl56z6);
assign Wl56z6 = (~(Pnb7z6[12] & Znnov6));
assign Ol56z6 = (~(Qdcdt6 & Fhc7z6[12]));
assign Ao46z6 = (Em56z6 & Mm56z6);
assign Mm56z6 = (Um56z6 & Cn56z6);
assign Cn56z6 = (Kn56z6 & Sn56z6);
assign Sn56z6 = (~(Ao56z6 & Oz3nv6));
assign Ao56z6 = (X4ciw6 ^ HADDRI[11]);
assign HADDRI[11] = (Crcdt6 ? Dvc7z6[11] : X0d7z6[11]);
assign X0d7z6[11] = (~(Io56z6 & Qo56z6));
assign Qo56z6 = (Yo56z6 & Gp56z6);
assign Gp56z6 = (~(Pic7z6[11] & Ir0ov6));
assign Yo56z6 = (Op56z6 & Wp56z6);
assign Wp56z6 = (Qs46z6 | Eqznv6);
assign Eqznv6 = (Eq56z6 & Mq56z6);
assign Mq56z6 = (~(Wkd7z6[11] & Ddmhw6));
assign Eq56z6 = (Uq56z6 & Cr56z6);
assign Cr56z6 = (~(Xhd7z6[11] & Eu46z6));
assign Uq56z6 = (~(Vnd7z6[11] & Jamnv6));
assign Op56z6 = (~(Pdc7z6[11] & Mu46z6));
assign Io56z6 = (Kr56z6 & Sr56z6);
assign Sr56z6 = (~(Pnb7z6[11] & Znnov6));
assign Kr56z6 = (~(Qdcdt6 & Fhc7z6[11]));
assign Kn56z6 = (~(As56z6 & Is56z6));
assign As56z6 = (D1ciw6 ^ HADDRI[10]);
assign HADDRI[10] = (Crcdt6 ? Dvc7z6[10] : X0d7z6[10]);
assign X0d7z6[10] = (~(Qs56z6 & Ys56z6));
assign Ys56z6 = (Gt56z6 & Ot56z6);
assign Ot56z6 = (~(Pic7z6[10] & Ir0ov6));
assign Gt56z6 = (Wt56z6 & Eu56z6);
assign Eu56z6 = (Qs46z6 | Fuznv6);
assign Fuznv6 = (Mu56z6 & Uu56z6);
assign Uu56z6 = (~(Wkd7z6[10] & Ddmhw6));
assign Mu56z6 = (Cv56z6 & Kv56z6);
assign Kv56z6 = (~(Xhd7z6[10] & Eu46z6));
assign Cv56z6 = (~(Vnd7z6[10] & Jamnv6));
assign Wt56z6 = (~(Pdc7z6[10] & Mu46z6));
assign Qs56z6 = (Sv56z6 & Aw56z6);
assign Aw56z6 = (~(Pnb7z6[10] & Znnov6));
assign Sv56z6 = (~(Qdcdt6 & Fhc7z6[10]));
assign Um56z6 = (Iw56z6 & Qw56z6);
assign Qw56z6 = (~(Yw56z6 & Rq3nv6));
assign Yw56z6 = (Nzbiw6 ^ HADDRI[9]);
assign HADDRI[9] = (Crcdt6 ? Dvc7z6[9] : X0d7z6[9]);
assign X0d7z6[9] = (~(Gx56z6 & Ox56z6));
assign Ox56z6 = (Wx56z6 & Ey56z6);
assign Ey56z6 = (~(Pic7z6[9] & Ir0ov6));
assign Wx56z6 = (My56z6 & Uy56z6);
assign Uy56z6 = (Qs46z6 | Gyznv6);
assign Gyznv6 = (Cz56z6 & Kz56z6);
assign Kz56z6 = (~(Wkd7z6[9] & Ddmhw6));
assign Cz56z6 = (Sz56z6 & A066z6);
assign A066z6 = (~(Xhd7z6[9] & Eu46z6));
assign Sz56z6 = (~(Vnd7z6[9] & Jamnv6));
assign My56z6 = (~(Pdc7z6[9] & Mu46z6));
assign Gx56z6 = (I066z6 & Q066z6);
assign Q066z6 = (~(Qti7z6[9] & Znnov6));
assign I066z6 = (~(Qdcdt6 & Fhc7z6[9]));
assign Iw56z6 = (~(Y066z6 & Ty3nv6));
assign Y066z6 = (M606z6 ^ G166z6);
assign M606z6 = (!HADDRI[8]);
assign HADDRI[8] = (Crcdt6 ? Dvc7z6[8] : X0d7z6[8]);
assign X0d7z6[8] = (~(O166z6 & W166z6));
assign W166z6 = (E266z6 & M266z6);
assign M266z6 = (~(Pdc7z6[8] & Mu46z6));
assign E266z6 = (U266z6 & C366z6);
assign C366z6 = (~(Znnov6 & K366z6));
assign K366z6 = (Qti7z6[8] | P2j7z6[6]);
assign U266z6 = (Qs46z6 | H20ov6);
assign H20ov6 = (S366z6 & A466z6);
assign A466z6 = (~(Wkd7z6[8] & Ddmhw6));
assign S366z6 = (I466z6 & Q466z6);
assign Q466z6 = (~(Xhd7z6[8] & Eu46z6));
assign I466z6 = (~(Vnd7z6[8] & Jamnv6));
assign O166z6 = (Y466z6 & G566z6);
assign G566z6 = (~(Pic7z6[8] & Ir0ov6));
assign Y466z6 = (~(Qdcdt6 & Fhc7z6[8]));
assign Em56z6 = (O566z6 & W566z6);
assign W566z6 = (~(E666z6 & Gv3nv6));
assign E666z6 = (Bkfnv6 ^ G5diw6);
assign O566z6 = (M666z6 & U666z6);
assign U666z6 = (~(C766z6 & Ve3nv6));
assign C766z6 = (Iw77z6 ^ Eg3nv6);
assign Eg3nv6 = (!Njfnv6);
assign M666z6 = (~(K766z6 & En3nv6));
assign K766z6 = (W6diw6 ^ Ujfnv6);
assign W6diw6 = (!Ey77z6);
assign Kn46z6 = (S766z6 & A866z6);
assign A866z6 = (I866z6 & Q866z6);
assign Q866z6 = (Y866z6 & G966z6);
assign G966z6 = (O966z6 & W966z6);
assign W966z6 = (~(Ea66z6 & Ma66z6));
assign Ea66z6 = (Q3diw6 ^ HADDRI[28]);
assign HADDRI[28] = (Crcdt6 ? Dvc7z6[28] : X0d7z6[28]);
assign X0d7z6[28] = (~(Ua66z6 & Cb66z6));
assign Cb66z6 = (Kb66z6 & Sb66z6);
assign Sb66z6 = (~(Pic7z6[28] & Ir0ov6));
assign Kb66z6 = (Ac66z6 & Ic66z6);
assign Ic66z6 = (Qs46z6 | Bnxnv6);
assign Bnxnv6 = (Qc66z6 & Yc66z6);
assign Yc66z6 = (~(Wkd7z6[28] & Ddmhw6));
assign Qc66z6 = (Gd66z6 & Od66z6);
assign Od66z6 = (~(Xhd7z6[28] & Eu46z6));
assign Gd66z6 = (~(Vnd7z6[28] & Jamnv6));
assign Ac66z6 = (~(Pdc7z6[28] & Mu46z6));
assign Ua66z6 = (Wd66z6 & Ee66z6);
assign Ee66z6 = (~(Pnb7z6[28] & Znnov6));
assign Wd66z6 = (~(Qdcdt6 & Fhc7z6[28]));
assign O966z6 = (~(Me66z6 & Qm3nv6));
assign Me66z6 = (M1diw6 ^ HADDRI[27]);
assign HADDRI[27] = (Crcdt6 ? Dvc7z6[27] : X0d7z6[27]);
assign X0d7z6[27] = (~(Ue66z6 & Cf66z6));
assign Cf66z6 = (Kf66z6 & Sf66z6);
assign Sf66z6 = (~(Pic7z6[27] & Ir0ov6));
assign Kf66z6 = (Ag66z6 & Ig66z6);
assign Ig66z6 = (Qs46z6 | Qrxnv6);
assign Qrxnv6 = (Qg66z6 & Yg66z6);
assign Yg66z6 = (~(Wkd7z6[27] & Ddmhw6));
assign Qg66z6 = (Gh66z6 & Oh66z6);
assign Oh66z6 = (~(Xhd7z6[27] & Eu46z6));
assign Gh66z6 = (~(Vnd7z6[27] & Jamnv6));
assign Ag66z6 = (~(Pdc7z6[27] & Mu46z6));
assign Ue66z6 = (Wh66z6 & Ei66z6);
assign Ei66z6 = (~(Pnb7z6[27] & Znnov6));
assign Wh66z6 = (~(Qdcdt6 & Fhc7z6[27]));
assign Y866z6 = (Mi66z6 & Ui66z6);
assign Ui66z6 = (~(Cj66z6 & Su3nv6));
assign Cj66z6 = (Wzciw6 ^ HADDRI[26]);
assign HADDRI[26] = (Crcdt6 ? Dvc7z6[26] : X0d7z6[26]);
assign X0d7z6[26] = (~(Kj66z6 & Sj66z6));
assign Sj66z6 = (Ak66z6 & Ik66z6);
assign Ik66z6 = (~(Pic7z6[26] & Ir0ov6));
assign Ak66z6 = (Qk66z6 & Yk66z6);
assign Yk66z6 = (Qs46z6 | Fwxnv6);
assign Fwxnv6 = (Gl66z6 & Ol66z6);
assign Ol66z6 = (~(Wkd7z6[26] & Ddmhw6));
assign Gl66z6 = (Wl66z6 & Em66z6);
assign Em66z6 = (~(Xhd7z6[26] & Eu46z6));
assign Wl66z6 = (~(Vnd7z6[26] & Jamnv6));
assign Qk66z6 = (~(Pdc7z6[26] & Mu46z6));
assign Kj66z6 = (Mm66z6 & Um66z6);
assign Um66z6 = (~(Pnb7z6[26] & Znnov6));
assign Mm66z6 = (~(Qdcdt6 & Fhc7z6[26]));
assign Wzciw6 = (!Yw77z6);
assign Mi66z6 = (~(Cn66z6 & Jf3nv6));
assign Cn66z6 = (Bqmyx6 ^ Kn66z6);
assign Bqmyx6 = (!HADDRI[25]);
assign HADDRI[25] = (Crcdt6 ? Dvc7z6[25] : X0d7z6[25]);
assign X0d7z6[25] = (~(Sn66z6 & Ao66z6));
assign Ao66z6 = (Io66z6 & Qo66z6);
assign Qo66z6 = (~(Pic7z6[25] & Ir0ov6));
assign Io66z6 = (Yo66z6 & Gp66z6);
assign Gp66z6 = (Qs46z6 | U0ynv6);
assign U0ynv6 = (Op66z6 & Wp66z6);
assign Wp66z6 = (~(Wkd7z6[25] & Ddmhw6));
assign Op66z6 = (Eq66z6 & Mq66z6);
assign Mq66z6 = (~(Xhd7z6[25] & Eu46z6));
assign Eq66z6 = (~(Vnd7z6[25] & Jamnv6));
assign Yo66z6 = (~(Pdc7z6[25] & Mu46z6));
assign Sn66z6 = (Uq66z6 & Cr66z6);
assign Cr66z6 = (~(Pnb7z6[25] & Znnov6));
assign Uq66z6 = (~(Qdcdt6 & Fhc7z6[25]));
assign I866z6 = (Kr66z6 & Sr66z6);
assign Sr66z6 = (~(As66z6 & Zg3nv6));
assign As66z6 = (Sqciw6 ^ HADDRI[22]);
assign HADDRI[22] = (Crcdt6 ? Dvc7z6[22] : X0d7z6[22]);
assign X0d7z6[22] = (~(Is66z6 & Qs66z6));
assign Qs66z6 = (Ys66z6 & Gt66z6);
assign Gt66z6 = (~(Pic7z6[22] & Ir0ov6));
assign Ys66z6 = (Ot66z6 & Wt66z6);
assign Wt66z6 = (Qs46z6 | Zdynv6);
assign Zdynv6 = (Eu66z6 & Mu66z6);
assign Mu66z6 = (~(Wkd7z6[22] & Ddmhw6));
assign Eu66z6 = (Uu66z6 & Cv66z6);
assign Cv66z6 = (~(Xhd7z6[22] & Eu46z6));
assign Uu66z6 = (~(Vnd7z6[22] & Jamnv6));
assign Ot66z6 = (~(Pdc7z6[22] & Mu46z6));
assign Is66z6 = (Kv66z6 & Sv66z6);
assign Sv66z6 = (~(Pnb7z6[22] & Znnov6));
assign Kv66z6 = (~(Qdcdt6 & Fhc7z6[22]));
assign Kr66z6 = (Aw66z6 & Iw66z6);
assign Iw66z6 = (~(Qw66z6 & Bp3nv6));
assign Qw66z6 = (Xwciw6 ^ HADDRI[24]);
assign HADDRI[24] = (Crcdt6 ? Dvc7z6[24] : X0d7z6[24]);
assign X0d7z6[24] = (~(Yw66z6 & Gx66z6));
assign Gx66z6 = (Ox66z6 & Wx66z6);
assign Wx66z6 = (~(Pic7z6[24] & Ir0ov6));
assign Ox66z6 = (Ey66z6 & My66z6);
assign My66z6 = (Qs46z6 | J5ynv6);
assign J5ynv6 = (Uy66z6 & Cz66z6);
assign Cz66z6 = (~(Wkd7z6[24] & Ddmhw6));
assign Uy66z6 = (Kz66z6 & Sz66z6);
assign Sz66z6 = (~(Xhd7z6[24] & Eu46z6));
assign Kz66z6 = (~(Vnd7z6[24] & Jamnv6));
assign Ey66z6 = (~(Pdc7z6[24] & Mu46z6));
assign Yw66z6 = (A076z6 & I076z6);
assign I076z6 = (~(Pnb7z6[24] & Znnov6));
assign A076z6 = (~(Qdcdt6 & Fhc7z6[24]));
assign Xwciw6 = (!Qw77z6);
assign Aw66z6 = (~(Q076z6 & Kx3nv6));
assign Q076z6 = (Psciw6 ^ HADDRI[23]);
assign HADDRI[23] = (Crcdt6 ? Dvc7z6[23] : X0d7z6[23]);
assign X0d7z6[23] = (~(Y076z6 & G176z6));
assign G176z6 = (O176z6 & W176z6);
assign W176z6 = (~(Pic7z6[23] & Ir0ov6));
assign O176z6 = (E276z6 & M276z6);
assign M276z6 = (Qs46z6 | K9ynv6);
assign K9ynv6 = (U276z6 & C376z6);
assign C376z6 = (~(Wkd7z6[23] & Ddmhw6));
assign U276z6 = (K376z6 & S376z6);
assign S376z6 = (~(Xhd7z6[23] & Eu46z6));
assign K376z6 = (~(Vnd7z6[23] & Jamnv6));
assign E276z6 = (~(Pdc7z6[23] & Mu46z6));
assign Y076z6 = (A476z6 & I476z6);
assign I476z6 = (~(Pnb7z6[23] & Znnov6));
assign A476z6 = (~(Qdcdt6 & Fhc7z6[23]));
assign Psciw6 = (!Yk77z6);
assign S766z6 = (Q476z6 & Y476z6);
assign Y476z6 = (G576z6 & O576z6);
assign O576z6 = (W576z6 & E676z6);
assign E676z6 = (~(M676z6 & U676z6));
assign M676z6 = (Cpciw6 ^ HADDRI[21]);
assign HADDRI[21] = (Crcdt6 ? Dvc7z6[21] : X0d7z6[21]);
assign X0d7z6[21] = (~(C776z6 & K776z6));
assign K776z6 = (S776z6 & A876z6);
assign A876z6 = (~(Pic7z6[21] & Ir0ov6));
assign S776z6 = (I876z6 & Q876z6);
assign Q876z6 = (Qs46z6 | Oiynv6);
assign Oiynv6 = (Y876z6 & G976z6);
assign G976z6 = (~(Wkd7z6[21] & Ddmhw6));
assign Y876z6 = (O976z6 & W976z6);
assign W976z6 = (~(Xhd7z6[21] & Eu46z6));
assign O976z6 = (~(Vnd7z6[21] & Jamnv6));
assign I876z6 = (~(Pdc7z6[21] & Mu46z6));
assign C776z6 = (Ea76z6 & Ma76z6);
assign Ma76z6 = (~(Pnb7z6[21] & Znnov6));
assign Ea76z6 = (~(Qdcdt6 & Fhc7z6[21]));
assign Cpciw6 = (!E287z6);
assign W576z6 = (~(Ua76z6 & Ww3nv6));
assign Ua76z6 = (Rmciw6 ^ HADDRI[20]);
assign HADDRI[20] = (Crcdt6 ? Dvc7z6[20] : X0d7z6[20]);
assign X0d7z6[20] = (~(Cb76z6 & Kb76z6));
assign Kb76z6 = (Sb76z6 & Ac76z6);
assign Ac76z6 = (~(Pic7z6[20] & Ir0ov6));
assign Sb76z6 = (Ic76z6 & Qc76z6);
assign Qc76z6 = (Qs46z6 | Dnynv6);
assign Dnynv6 = (Yc76z6 & Gd76z6);
assign Gd76z6 = (~(Wkd7z6[20] & Ddmhw6));
assign Yc76z6 = (Od76z6 & Wd76z6);
assign Wd76z6 = (~(Xhd7z6[20] & Eu46z6));
assign Od76z6 = (~(Vnd7z6[20] & Jamnv6));
assign Ic76z6 = (~(Pdc7z6[20] & Mu46z6));
assign Cb76z6 = (Ee76z6 & Me76z6);
assign Me76z6 = (~(Pnb7z6[20] & Znnov6));
assign Ee76z6 = (~(Qdcdt6 & Fhc7z6[20]));
assign Rmciw6 = (!G187z6);
assign G576z6 = (Ue76z6 & Cf76z6);
assign Cf76z6 = (~(Kf76z6 & Mk3nv6));
assign Kf76z6 = (Blciw6 ^ HADDRI[19]);
assign HADDRI[19] = (Crcdt6 ? Dvc7z6[19] : X0d7z6[19]);
assign X0d7z6[19] = (~(Sf76z6 & Ag76z6));
assign Ag76z6 = (Ig76z6 & Qg76z6);
assign Qg76z6 = (~(Pic7z6[19] & Ir0ov6));
assign Ig76z6 = (Yg76z6 & Gh76z6);
assign Gh76z6 = (Qs46z6 | Srynv6);
assign Srynv6 = (Oh76z6 & Wh76z6);
assign Wh76z6 = (~(Wkd7z6[19] & Ddmhw6));
assign Oh76z6 = (Ei76z6 & Mi76z6);
assign Mi76z6 = (~(Xhd7z6[19] & Eu46z6));
assign Ei76z6 = (~(Vnd7z6[19] & Jamnv6));
assign Yg76z6 = (~(Pdc7z6[19] & Mu46z6));
assign Sf76z6 = (Ui76z6 & Cj76z6);
assign Cj76z6 = (~(Pnb7z6[19] & Znnov6));
assign Ui76z6 = (~(Qdcdt6 & Fhc7z6[19]));
assign Ue76z6 = (~(Kj76z6 & Vs3nv6));
assign Kj76z6 = (Ljciw6 ^ HADDRI[18]);
assign HADDRI[18] = (Crcdt6 ? Dvc7z6[18] : X0d7z6[18]);
assign X0d7z6[18] = (~(Sj76z6 & Ak76z6));
assign Ak76z6 = (Ik76z6 & Qk76z6);
assign Qk76z6 = (~(Pic7z6[18] & Ir0ov6));
assign Ik76z6 = (Yk76z6 & Gl76z6);
assign Gl76z6 = (Qs46z6 | Hwynv6);
assign Hwynv6 = (Ol76z6 & Wl76z6);
assign Wl76z6 = (~(Wkd7z6[18] & Ddmhw6));
assign Ol76z6 = (Em76z6 & Mm76z6);
assign Mm76z6 = (~(Xhd7z6[18] & Eu46z6));
assign Em76z6 = (~(Vnd7z6[18] & Jamnv6));
assign Yk76z6 = (~(Pdc7z6[18] & Mu46z6));
assign Sj76z6 = (Um76z6 & Cn76z6);
assign Cn76z6 = (~(Pnb7z6[18] & Znnov6));
assign Um76z6 = (~(Qdcdt6 & Fhc7z6[18]));
assign Q476z6 = (Kn76z6 & Sn76z6);
assign Kn76z6 = (Ao76z6 & Io76z6);
assign Io76z6 = (~(Qo76z6 & X04nv6));
assign Qo76z6 = (Vhciw6 ^ HADDRI[17]);
assign HADDRI[17] = (Crcdt6 ? Dvc7z6[17] : X0d7z6[17]);
assign X0d7z6[17] = (~(Yo76z6 & Gp76z6));
assign Gp76z6 = (Op76z6 & Wp76z6);
assign Wp76z6 = (~(Pic7z6[17] & Ir0ov6));
assign Op76z6 = (Eq76z6 & Mq76z6);
assign Mq76z6 = (Qs46z6 | W0znv6);
assign W0znv6 = (Uq76z6 & Cr76z6);
assign Cr76z6 = (~(Wkd7z6[17] & Ddmhw6));
assign Uq76z6 = (Kr76z6 & Sr76z6);
assign Sr76z6 = (~(Xhd7z6[17] & Eu46z6));
assign Kr76z6 = (~(Vnd7z6[17] & Jamnv6));
assign Eq76z6 = (~(Pdc7z6[17] & Mu46z6));
assign Yo76z6 = (As76z6 & Is76z6);
assign Is76z6 = (~(Pnb7z6[17] & Znnov6));
assign As76z6 = (~(Qdcdt6 & Fhc7z6[17]));
assign Vhciw6 = (!W187z6);
assign Ao76z6 = (~(Qs76z6 & Ys76z6));
assign Qs76z6 = (Wl06z6 ^ Gt76z6);
assign Wl06z6 = (!HADDRI[16]);
assign HADDRI[16] = (Crcdt6 ? Dvc7z6[16] : X0d7z6[16]);
assign X0d7z6[16] = (~(Ot76z6 & Wt76z6));
assign Wt76z6 = (Eu76z6 & Mu76z6);
assign Mu76z6 = (~(Pic7z6[16] & Ir0ov6));
assign Eu76z6 = (Uu76z6 & Cv76z6);
assign Cv76z6 = (Qs46z6 | L5znv6);
assign L5znv6 = (Kv76z6 & Sv76z6);
assign Sv76z6 = (~(Wkd7z6[16] & Ddmhw6));
assign Kv76z6 = (Aw76z6 & Iw76z6);
assign Iw76z6 = (~(Xhd7z6[16] & Eu46z6));
assign Aw76z6 = (~(Vnd7z6[16] & Jamnv6));
assign Uu76z6 = (~(Pdc7z6[16] & Mu46z6));
assign Ot76z6 = (Qw76z6 & Yw76z6);
assign Yw76z6 = (~(Pnb7z6[16] & Znnov6));
assign Qw76z6 = (~(Qdcdt6 & Fhc7z6[16]));
assign Agz5z6 = (!HPROTI[1]);
assign Kconv6 = (~(Gx76z6 & Ox76z6));
assign Ox76z6 = (Njkiw6 ? Ey76z6 : Wx76z6);
assign Ey76z6 = (~(My76z6 & Uy76z6));
assign My76z6 = (HREADYI & Cfliy6);
assign Wx76z6 = (~(Cz76z6 & Ykyiy6));
assign Ykyiy6 = (Kz76z6 & Sz76z6);
assign Sz76z6 = (Pbonv6 & Ag0jy6);
assign Pbonv6 = (~(Ewyet6 | Styet6));
assign Kz76z6 = (A086z6 & I086z6);
assign A086z6 = (~(K4bdt6 & Q086z6));
assign Cz76z6 = (~(E6y5z6 | Meoet6));
assign E6y5z6 = (~(D6eiw6 & Y086z6));
assign Y086z6 = (~(Yk0jy6 & G186z6));
assign G186z6 = (Gl0jy6 | Zuixx6);
assign Zuixx6 = (!HREADYS);
assign Gl0jy6 = (~(Qk0jy6 & O186z6));
assign O186z6 = (S3v5z6 | Qln7z6[1]);
assign S3v5z6 = (W186z6 & Bwixx6);
assign Yk0jy6 = (E286z6 & M286z6);
assign M286z6 = (~(U286z6 & HREADYD));
assign U286z6 = (!Qk0jy6);
assign Qk0jy6 = (~(C386z6 & Hm1ov6));
assign C386z6 = (~(Zblov6 | Qln7z6[1]));
assign E286z6 = (A4v5z6 & Ag0jy6);
assign A4v5z6 = (Goonv6 | Ik0jy6);
assign Ik0jy6 = (W186z6 & K386z6);
assign K386z6 = (Bwixx6 | Qln7z6[1]);
assign Bwixx6 = (V4myx6 | Go9ov6);
assign Goonv6 = (!HREADYD);
assign D6eiw6 = (~(Djonv6 | S386z6));
assign S386z6 = (Kb0jy6 & Rxixx6);
assign Gx76z6 = (Lbkiw6 & Ikyiy6);
assign Ikyiy6 = (!Bkkiw6);
assign Bkkiw6 = (A486z6 & Ujfnv6);
assign A486z6 = (Njfnv6 & Bkfnv6);
assign Rnh7v6 = (~(I486z6 & Q486z6));
assign Q486z6 = (~(J72nz6[1] & Szw5z6));
assign I486z6 = (Y486z6 & G586z6);
assign G586z6 = (~(Y0x5z6 & O586z6));
assign O586z6 = (~(W586z6 & E686z6));
assign E686z6 = (M686z6 & U686z6);
assign U686z6 = (~(S3x5z6 & Yr1nz6[1]));
assign S3x5z6 = (Md1nz6[0] & Rn5ov6);
assign M686z6 = (~(E2x5z6 & Au1nz6[1]));
assign E2x5z6 = (~(Rn5ov6 | Md1nz6[0]));
assign W586z6 = (C786z6 & K786z6);
assign K786z6 = (~(Jq5ov6 & Bv1nz6[1]));
assign Jq5ov6 = (Rn5ov6 & S786z6);
assign C786z6 = (~(Qq5ov6 & Zs1nz6[1]));
assign Qq5ov6 = (~(Rn5ov6 | S786z6));
assign S786z6 = (!Md1nz6[0]);
assign Rn5ov6 = (Md1nz6[1] ^ Md1nz6[2]);
assign Y0x5z6 = (~(A886z6 | Szw5z6));
assign A886z6 = (~(Hp5ov6 & Dxiyx6));
assign Dxiyx6 = (!Vp5ov6);
assign Y486z6 = (~(Q0y5z6 & Zejyx6));
assign Zejyx6 = (~(I886z6 & Q886z6));
assign Q886z6 = (Y886z6 & G986z6);
assign G986z6 = (~(G5x5z6 & Mm1nz6[1]));
assign G5x5z6 = (~(O986z6 | N43yx6));
assign Y886z6 = (~(O5x5z6 & Oo1nz6[1]));
assign O5x5z6 = (~(R63yx6 | Yb1nz6[0]));
assign I886z6 = (W986z6 & Ea86z6);
assign Ea86z6 = (~(Z63yx6 & Pp1nz6[1]));
assign Z63yx6 = (R63yx6 & O986z6);
assign O986z6 = (!Yb1nz6[0]);
assign W986z6 = (~(H73yx6 & Nn1nz6[1]));
assign H73yx6 = (N43yx6 & Yb1nz6[0]);
assign N43yx6 = (!R63yx6);
assign R63yx6 = (Yb1nz6[1] ^ Yb1nz6[2]);
assign Q0y5z6 = (!L53yx6);
assign L53yx6 = (~(Ma86z6 & Vp5ov6));
assign Vp5ov6 = (Ua86z6 & Cb86z6);
assign Cb86z6 = (~(Kb86z6 & Qa2nz6[0]));
assign Kb86z6 = (Sb86z6 & Ac86z6);
assign Sb86z6 = (~(Qa2nz6[1] & Ic86z6));
assign Ua86z6 = (Qa2nz6[1] ? Yc86z6 : Qc86z6);
assign Yc86z6 = (Gd86z6 & Od86z6);
assign Gd86z6 = (Wd86z6 | Qc86z6);
assign Wd86z6 = (Qa2nz6[0] ? Me86z6 : Ee86z6);
assign Ee86z6 = (~(X7iyx6 & Ue86z6));
assign Ue86z6 = (~(Ju2yx6 & D53yx6));
assign Qc86z6 = (~(Ic86z6 & Cf86z6));
assign Cf86z6 = (~(Me86z6 & Ju2yx6));
assign Ma86z6 = (~(Szw5z6 | Hp5ov6));
assign Hp5ov6 = (Qa2nz6[1] ? Sf86z6 : Kf86z6);
assign Sf86z6 = (Ag86z6 & Od86z6);
assign Od86z6 = (~(Qa2nz6[0] & Ig86z6));
assign Ig86z6 = (~(X7iyx6 & Ns2yx6));
assign Ag86z6 = (~(Qg86z6 & Yg86z6));
assign Yg86z6 = (~(Gh86z6 & Qa2nz6[0]));
assign Gh86z6 = (Oh86z6 & Ic86z6);
assign Qg86z6 = (D53yx6 | Ac86z6);
assign Ac86z6 = (~(Wh86z6 & Ju2yx6));
assign Wh86z6 = (Ic86z6 & X7iyx6);
assign Kf86z6 = (~(Ei86z6 & Mi86z6));
assign Mi86z6 = (~(Ui86z6 & Qa2nz6[0]));
assign Ei86z6 = (Cj86z6 & Ic86z6);
assign Cj86z6 = (~(Oh86z6 & Ju2yx6));
assign Oh86z6 = (~(Me86z6 & D53yx6));
assign Szw5z6 = (Op5ov6 | B63yx6);
assign B63yx6 = (~(M81nv6 | Lge7v6));
assign M81nv6 = (!Twhiw6);
assign Op5ov6 = (F2f7v6 & Kj86z6);
assign Kj86z6 = (~(Sj86z6 & Ryiyx6));
assign Ryiyx6 = (Lx2yx6 & J23yx6);
assign Lx2yx6 = (~(Ak86z6 & Ik86z6));
assign Ik86z6 = (~(Qk86z6 & L5iyx6));
assign L5iyx6 = (Otv5z6 & Eb1nv6);
assign Eb1nv6 = (!Ec2nz6[1]);
assign Qk86z6 = (J7f7v6 & F8iyx6);
assign F8iyx6 = (!T5f7v6);
assign Ak86z6 = (Yk86z6 & Krv5z6);
assign Yk86z6 = (~(T5iyx6 & J7f7v6));
assign T5iyx6 = (Gl86z6 & Ol86z6);
assign Ol86z6 = (~(Wl86z6 & Em86z6));
assign Em86z6 = (Mm86z6 & Um86z6);
assign Um86z6 = (Otv5z6 & Ec2nz6[1]);
assign Mm86z6 = (T32nz6[0] & Ec2nz6[0]);
assign Wl86z6 = (T13yx6 & T32nz6[3]);
assign T13yx6 = (T32nz6[2] & T32nz6[1]);
assign Gl86z6 = (~(Ui86z6 | H7iyx6));
assign H7iyx6 = (Cn86z6 & Ic86z6);
assign Ic86z6 = (~(Kn86z6 & J7f7v6));
assign Kn86z6 = (Sn86z6 & X7iyx6);
assign X7iyx6 = (!Ui86z6);
assign Sn86z6 = (~(Ao86z6 & Io86z6));
assign Ao86z6 = (V91nv6 & J23yx6);
assign J23yx6 = (~(Qo86z6 & Otv5z6));
assign Qo86z6 = (Ec2nz6[1] & Ns2yx6);
assign Cn86z6 = (~(Yo86z6 & Gp86z6));
assign Gp86z6 = (Me86z6 ? Wp86z6 : Op86z6);
assign Me86z6 = (!Fo5ov6);
assign Fo5ov6 = (~(Eq86z6 & Mq86z6));
assign Mq86z6 = (~(Md1nz6[2] ^ Fg1nz6[2]));
assign Eq86z6 = (Uq86z6 & Cr86z6);
assign Cr86z6 = (~(Md1nz6[1] ^ Fg1nz6[1]));
assign Uq86z6 = (~(Md1nz6[0] ^ Fg1nz6[0]));
assign Wp86z6 = (S3w5z6 & Kr86z6);
assign Kr86z6 = (~(D53yx6 & Nwiyx6));
assign Op86z6 = (~(S3w5z6 & Nwiyx6));
assign Nwiyx6 = (!Qa2nz6[1]);
assign Yo86z6 = (Sr86z6 & Ju2yx6);
assign Ju2yx6 = (~(As86z6 & Is86z6));
assign Is86z6 = (Qs86z6 & Ys86z6);
assign Ys86z6 = (~(Gt86z6 & Ot86z6));
assign Ot86z6 = (~(Ca1nv6 & T81nv6));
assign T81nv6 = (!J7f7v6);
assign Ca1nv6 = (D92nz6[1] & D92nz6[0]);
assign Gt86z6 = (Krv5z6 | Xrjyx6);
assign Xrjyx6 = (!Io86z6);
assign Krv5z6 = (~(J7f7v6 & Ns2yx6));
assign Ns2yx6 = (!Ec2nz6[0]);
assign Qs86z6 = (~(Otv5z6 | B5e7v6));
assign Otv5z6 = (Ec2nz6[3] & Ec2nz6[2]);
assign As86z6 = (M8e7v6 & V91nv6);
assign Sr86z6 = (~(Qa2nz6[1] & Wt86z6));
assign Wt86z6 = (~(S3w5z6 & D53yx6));
assign D53yx6 = (~(Eu86z6 & Mu86z6));
assign Mu86z6 = (~(Yb1nz6[2] ^ Af1nz6[2]));
assign Eu86z6 = (Uu86z6 & Cv86z6);
assign Cv86z6 = (~(Yb1nz6[1] ^ Af1nz6[1]));
assign Uu86z6 = (~(Yb1nz6[0] ^ Af1nz6[0]));
assign S3w5z6 = (!Qa2nz6[0]);
assign Ui86z6 = (T5f7v6 & Od77z6);
assign Sj86z6 = (Kv86z6 & Zyiyx6);
assign Zyiyx6 = (~(J7f7v6 & Sv86z6));
assign Sv86z6 = (~(Io86z6 & V91nv6));
assign V91nv6 = (~(Rm2yx6 | Ywv5z6));
assign Ywv5z6 = (!Wxv5z6);
assign Wxv5z6 = (B2jyx6 & Xf2yx6);
assign Xf2yx6 = (Vuf7v6 & V0jyx6);
assign V0jyx6 = (!Ctf7v6);
assign B2jyx6 = (Pb2yx6 & Tl2yx6);
assign Tl2yx6 = (!Mwf7v6);
assign Pb2yx6 = (!Qk77z6);
assign Rm2yx6 = (!J6jyx6);
assign J6jyx6 = (Aw86z6 & Kf2nz6[2]);
assign Aw86z6 = (Kf2nz6[1] & Kf2nz6[0]);
assign Io86z6 = (~(Xre7v6 | Iw86z6));
assign Iw86z6 = (~(Twhiw6 | J7f7v6));
assign Twhiw6 = (Nl1nz6[0] | Nl1nz6[1]);
assign Kv86z6 = (~(A4f7v6 & Ik77z6));
assign Py9dt6 = (~(Olvnv6 & Qw86z6));
assign Qw86z6 = (~(Ez9dt6 & Xkqnv6));
assign Ox9dt6 = (~(Olvnv6 & Yw86z6));
assign Yw86z6 = (~(Cy9dt6 & Xkqnv6));
assign Sz9dt6 = (~(Olvnv6 & Gx86z6));
assign Gx86z6 = (~(G0adt6 & Xkqnv6));
assign Xkqnv6 = (!RSTBYPASS);
assign Olvnv6 = (~(RSTBYPASS & PORESETn));
assign Tib7z6[9] = (Kn97z6 | INTISR[9]);
assign Tib7z6[8] = (Sn97z6 | INTISR[8]);
assign Tib7z6[7] = (Ao97z6 | INTISR[7]);
assign Tib7z6[6] = (Io97z6 | INTISR[6]);
assign Tib7z6[63] = (U697z6 | INTISR[63]);
assign Tib7z6[62] = (C797z6 | INTISR[62]);
assign Tib7z6[61] = (K797z6 | INTISR[61]);
assign Tib7z6[60] = (S797z6 | INTISR[60]);
assign Tib7z6[5] = (Qo97z6 | INTISR[5]);
assign Tib7z6[59] = (A897z6 | INTISR[59]);
assign Tib7z6[58] = (I897z6 | INTISR[58]);
assign Tib7z6[57] = (Q897z6 | INTISR[57]);
assign Tib7z6[56] = (Y897z6 | INTISR[56]);
assign Tib7z6[55] = (G997z6 | INTISR[55]);
assign Tib7z6[54] = (O997z6 | INTISR[54]);
assign Tib7z6[53] = (W997z6 | INTISR[53]);
assign Tib7z6[52] = (Ea97z6 | INTISR[52]);
assign Tib7z6[51] = (Ma97z6 | INTISR[51]);
assign Tib7z6[50] = (Ua97z6 | INTISR[50]);
assign Tib7z6[4] = (Yo97z6 | INTISR[4]);
assign Tib7z6[49] = (Cb97z6 | INTISR[49]);
assign Tib7z6[48] = (Kb97z6 | INTISR[48]);
assign Tib7z6[47] = (Sb97z6 | INTISR[47]);
assign Tib7z6[46] = (Ac97z6 | INTISR[46]);
assign Tib7z6[45] = (Ic97z6 | INTISR[45]);
assign Tib7z6[44] = (Qc97z6 | INTISR[44]);
assign Tib7z6[43] = (Yc97z6 | INTISR[43]);
assign Tib7z6[42] = (Gd97z6 | INTISR[42]);
assign Tib7z6[41] = (Od97z6 | INTISR[41]);
assign Tib7z6[40] = (Wd97z6 | INTISR[40]);
assign Tib7z6[3] = (Gp97z6 | INTISR[3]);
assign Tib7z6[39] = (Ee97z6 | INTISR[39]);
assign Tib7z6[38] = (Me97z6 | INTISR[38]);
assign Tib7z6[37] = (Ue97z6 | INTISR[37]);
assign Tib7z6[36] = (Cf97z6 | INTISR[36]);
assign Tib7z6[35] = (Kf97z6 | INTISR[35]);
assign Tib7z6[34] = (Sf97z6 | INTISR[34]);
assign Tib7z6[33] = (Ag97z6 | INTISR[33]);
assign Tib7z6[32] = (Ig97z6 | INTISR[32]);
assign Tib7z6[31] = (Qg97z6 | INTISR[31]);
assign Tib7z6[30] = (Yg97z6 | INTISR[30]);
assign Tib7z6[2] = (Op97z6 | INTISR[2]);
assign Tib7z6[29] = (Gh97z6 | INTISR[29]);
assign Tib7z6[28] = (Oh97z6 | INTISR[28]);
assign Tib7z6[27] = (Wh97z6 | INTISR[27]);
assign Tib7z6[26] = (Ei97z6 | INTISR[26]);
assign Tib7z6[25] = (Mi97z6 | INTISR[25]);
assign Tib7z6[24] = (Ui97z6 | INTISR[24]);
assign Tib7z6[23] = (Cj97z6 | INTISR[23]);
assign Tib7z6[22] = (Kj97z6 | INTISR[22]);
assign Tib7z6[21] = (Sj97z6 | INTISR[21]);
assign Tib7z6[20] = (Ak97z6 | INTISR[20]);
assign Tib7z6[1] = (Wp97z6 | INTISR[1]);
assign Tib7z6[19] = (Ik97z6 | INTISR[19]);
assign Tib7z6[18] = (Qk97z6 | INTISR[18]);
assign Tib7z6[17] = (Yk97z6 | INTISR[17]);
assign Tib7z6[16] = (Gl97z6 | INTISR[16]);
assign Tib7z6[15] = (Ol97z6 | INTISR[15]);
assign Tib7z6[14] = (Wl97z6 | INTISR[14]);
assign Tib7z6[13] = (Em97z6 | INTISR[13]);
assign Tib7z6[12] = (Mm97z6 | INTISR[12]);
assign Tib7z6[11] = (Um97z6 | INTISR[11]);
assign Tib7z6[10] = (Cn97z6 | INTISR[10]);
assign Tib7z6[0] = (Eq97z6 | INTISR[0]);
assign D4adt6 = (Knbdt6 & Wdtnv6);
assign Wdtnv6 = (!Wfo7v6);
assign S3adt6 = (Jgliw6 & Vb4iw6);
assign Jgliw6 = (~(Wy67v6 & Kygnv6));
assign Kygnv6 = (!HTMDHBURST[0]);
assign WAKEUP = (~(Ox86z6 & Wx86z6));
assign Wx86z6 = (Ey86z6 & My86z6);
assign My86z6 = (Uy86z6 & Cz86z6);
assign Cz86z6 = (Kz86z6 & Sz86z6);
assign Sz86z6 = (A096z6 & I096z6);
assign I096z6 = (Q096z6 & Y096z6);
assign Y096z6 = (~(Fjb7z6[3] & Eq97z6));
assign Q096z6 = (G196z6 & O196z6);
assign O196z6 = (~(Fjb7z6[1] & Uq97z6));
assign G196z6 = (~(Fjb7z6[2] & Mq97z6));
assign A096z6 = (W196z6 & E296z6);
assign E296z6 = (~(Fjb7z6[4] & Wp97z6));
assign W196z6 = (~(Fjb7z6[5] & Op97z6));
assign Kz86z6 = (M296z6 & U296z6);
assign U296z6 = (C396z6 & K396z6);
assign K396z6 = (~(Fjb7z6[6] & Gp97z6));
assign C396z6 = (~(Fjb7z6[7] & Yo97z6));
assign M296z6 = (S396z6 & A496z6);
assign A496z6 = (~(Fjb7z6[8] & Qo97z6));
assign S396z6 = (~(Fjb7z6[9] & Io97z6));
assign Uy86z6 = (I496z6 & Q496z6);
assign Q496z6 = (Y496z6 & G596z6);
assign G596z6 = (O596z6 & W596z6);
assign W596z6 = (~(Fjb7z6[10] & Ao97z6));
assign O596z6 = (~(Fjb7z6[11] & Sn97z6));
assign Y496z6 = (E696z6 & M696z6);
assign M696z6 = (~(Fjb7z6[12] & Kn97z6));
assign E696z6 = (~(Fjb7z6[13] & Cn97z6));
assign I496z6 = (U696z6 & C796z6);
assign C796z6 = (K796z6 & S796z6);
assign S796z6 = (~(Fjb7z6[14] & Um97z6));
assign K796z6 = (~(Fjb7z6[15] & Mm97z6));
assign U696z6 = (A896z6 & I896z6);
assign I896z6 = (~(Fjb7z6[16] & Em97z6));
assign A896z6 = (~(Fjb7z6[17] & Wl97z6));
assign Ey86z6 = (Q896z6 & Y896z6);
assign Y896z6 = (G996z6 & O996z6);
assign O996z6 = (W996z6 & Ea96z6);
assign Ea96z6 = (Ma96z6 & Ua96z6);
assign Ua96z6 = (~(Fjb7z6[20] & Yk97z6));
assign Ma96z6 = (Cb96z6 & Kb96z6);
assign Kb96z6 = (~(Fjb7z6[18] & Ol97z6));
assign Cb96z6 = (~(Fjb7z6[19] & Gl97z6));
assign W996z6 = (Sb96z6 & Ac96z6);
assign Ac96z6 = (~(Fjb7z6[21] & Qk97z6));
assign Sb96z6 = (~(Fjb7z6[22] & Ik97z6));
assign G996z6 = (Ic96z6 & Qc96z6);
assign Qc96z6 = (Yc96z6 & Gd96z6);
assign Gd96z6 = (~(Fjb7z6[23] & Ak97z6));
assign Yc96z6 = (~(Fjb7z6[24] & Sj97z6));
assign Ic96z6 = (Od96z6 & Wd96z6);
assign Wd96z6 = (~(Fjb7z6[25] & Kj97z6));
assign Od96z6 = (~(Fjb7z6[26] & Cj97z6));
assign Q896z6 = (Ee96z6 & Me96z6);
assign Me96z6 = (Ue96z6 & Cf96z6);
assign Cf96z6 = (Kf96z6 & Sf96z6);
assign Sf96z6 = (~(Fjb7z6[27] & Ui97z6));
assign Kf96z6 = (~(Fjb7z6[28] & Mi97z6));
assign Ue96z6 = (Ag96z6 & Ig96z6);
assign Ig96z6 = (~(Fjb7z6[29] & Ei97z6));
assign Ag96z6 = (~(Fjb7z6[30] & Wh97z6));
assign Ee96z6 = (Qg96z6 & Yg96z6);
assign Yg96z6 = (Gh96z6 & Oh96z6);
assign Oh96z6 = (~(Fjb7z6[31] & Oh97z6));
assign Gh96z6 = (~(Fjb7z6[32] & Gh97z6));
assign Qg96z6 = (Wh96z6 & Ei96z6);
assign Ei96z6 = (~(Fjb7z6[33] & Yg97z6));
assign Wh96z6 = (~(Fjb7z6[34] & Qg97z6));
assign Ox86z6 = (Mi96z6 & Ui96z6);
assign Ui96z6 = (Cj96z6 & Kj96z6);
assign Kj96z6 = (Sj96z6 & Ak96z6);
assign Ak96z6 = (Ik96z6 & Qk96z6);
assign Qk96z6 = (Yk96z6 & Gl96z6);
assign Gl96z6 = (~(Fjb7z6[37] & Sf97z6));
assign Yk96z6 = (Ol96z6 & Wl96z6);
assign Wl96z6 = (~(Fjb7z6[35] & Ig97z6));
assign Ol96z6 = (~(Fjb7z6[36] & Ag97z6));
assign Ik96z6 = (Em96z6 & Mm96z6);
assign Mm96z6 = (~(Fjb7z6[38] & Kf97z6));
assign Em96z6 = (~(Fjb7z6[39] & Cf97z6));
assign Sj96z6 = (Um96z6 & Cn96z6);
assign Cn96z6 = (Kn96z6 & Sn96z6);
assign Sn96z6 = (~(Fjb7z6[40] & Ue97z6));
assign Kn96z6 = (~(Fjb7z6[41] & Me97z6));
assign Um96z6 = (Ao96z6 & Io96z6);
assign Io96z6 = (~(Fjb7z6[42] & Ee97z6));
assign Ao96z6 = (~(Fjb7z6[43] & Wd97z6));
assign Cj96z6 = (Qo96z6 & Yo96z6);
assign Yo96z6 = (Gp96z6 & Op96z6);
assign Op96z6 = (Wp96z6 & Eq96z6);
assign Eq96z6 = (~(Fjb7z6[44] & Od97z6));
assign Wp96z6 = (~(Fjb7z6[45] & Gd97z6));
assign Gp96z6 = (Mq96z6 & Uq96z6);
assign Uq96z6 = (~(Fjb7z6[46] & Yc97z6));
assign Mq96z6 = (~(Fjb7z6[47] & Qc97z6));
assign Qo96z6 = (Cr96z6 & Kr96z6);
assign Kr96z6 = (Sr96z6 & As96z6);
assign As96z6 = (~(Fjb7z6[48] & Ic97z6));
assign Sr96z6 = (~(Fjb7z6[49] & Ac97z6));
assign Cr96z6 = (Is96z6 & Qs96z6);
assign Qs96z6 = (~(Fjb7z6[50] & Sb97z6));
assign Is96z6 = (~(Fjb7z6[51] & Kb97z6));
assign Mi96z6 = (Ys96z6 & Gt96z6);
assign Gt96z6 = (Ot96z6 & Wt96z6);
assign Wt96z6 = (Eu96z6 & Mu96z6);
assign Mu96z6 = (Uu96z6 & Cv96z6);
assign Cv96z6 = (~(Fjb7z6[52] & Cb97z6));
assign Uu96z6 = (~(Fjb7z6[53] & Ua97z6));
assign Eu96z6 = (Kv96z6 & Sv96z6);
assign Sv96z6 = (~(Fjb7z6[54] & Ma97z6));
assign Kv96z6 = (~(Fjb7z6[55] & Ea97z6));
assign Ot96z6 = (Aw96z6 & Iw96z6);
assign Iw96z6 = (Qw96z6 & Yw96z6);
assign Yw96z6 = (~(Fjb7z6[56] & W997z6));
assign Qw96z6 = (~(Fjb7z6[57] & O997z6));
assign Aw96z6 = (Gx96z6 & Ox96z6);
assign Ox96z6 = (~(Fjb7z6[58] & G997z6));
assign Gx96z6 = (~(Fjb7z6[59] & Y897z6));
assign Ys96z6 = (Wx96z6 & Ey96z6);
assign Ey96z6 = (My96z6 & Uy96z6);
assign Uy96z6 = (Cz96z6 & Kz96z6);
assign Kz96z6 = (~(Fjb7z6[60] & Q897z6));
assign Cz96z6 = (~(Fjb7z6[61] & I897z6));
assign My96z6 = (Sz96z6 & A0a6z6);
assign A0a6z6 = (~(Fjb7z6[62] & A897z6));
assign Sz96z6 = (~(Fjb7z6[63] & S797z6));
assign Wx96z6 = (I0a6z6 & Q0a6z6);
assign Q0a6z6 = (Y0a6z6 & G1a6z6);
assign G1a6z6 = (~(Fjb7z6[64] & K797z6));
assign Y0a6z6 = (~(Fjb7z6[65] & C797z6));
assign I0a6z6 = (O1a6z6 & W1a6z6);
assign W1a6z6 = (~(Fjb7z6[66] & U697z6));
assign O1a6z6 = (~(Ei77z6 & Fjb7z6[0]));
assign TXEV = (I2edt6 & Pxfov6);
assign SLEEPDEEP = (SLEEPING & U3cet6);
assign MEMATTRS[1] = (~(E2a6z6 & M2a6z6));
assign M2a6z6 = (~(Rj9ov6 & Qdqnv6));
assign Qdqnv6 = (~(U2a6z6 & C3a6z6));
assign C3a6z6 = (~(K3a6z6 & S3a6z6));
assign S3a6z6 = (A4a6z6 & Cmm7z6[29]);
assign A4a6z6 = (Yygnv6 & I4a6z6);
assign K3a6z6 = (Q4a6z6 & Cmm7z6[31]);
assign U2a6z6 = (Y4a6z6 & G5a6z6);
assign G5a6z6 = (~(O5a6z6 & W5a6z6));
assign W5a6z6 = (V5k7z6[31] & E6a6z6);
assign O5a6z6 = (~(M6a6z6 | U6a6z6));
assign Y4a6z6 = (~(C7a6z6 & K7a6z6));
assign C7a6z6 = (S7a6z6 & A8a6z6);
assign A8a6z6 = (~(I8a6z6 & Q8a6z6));
assign Q8a6z6 = (Y8a6z6 & G9a6z6);
assign G9a6z6 = (O9a6z6 & W9a6z6);
assign W9a6z6 = (~(P6l7z6[16] & Eaa6z6));
assign O9a6z6 = (Maa6z6 & Uaa6z6);
assign Uaa6z6 = (~(Cba6z6 & Kba6z6));
assign Maa6z6 = (~(Hwk7z6[16] & Sba6z6));
assign Y8a6z6 = (Aca6z6 & Ica6z6);
assign Ica6z6 = (~(Xgl7z6[16] & Qca6z6));
assign Aca6z6 = (~(Frl7z6[16] & Yca6z6));
assign I8a6z6 = (Gda6z6 & Oda6z6);
assign Oda6z6 = (Wda6z6 & Eea6z6);
assign Eea6z6 = (~(N1m7z6[16] & Mea6z6));
assign Wda6z6 = (~(Zlk7z6[16] & Uea6z6));
assign Gda6z6 = (Cfa6z6 & Kfa6z6);
assign Kfa6z6 = (~(Rbk7z6[16] & Sfa6z6));
assign Cfa6z6 = (~(Vbm7z6[16] & Aga6z6));
assign S7a6z6 = (~(Iga6z6 & Qga6z6));
assign Iga6z6 = (Kba6z6 & Yga6z6);
assign E2a6z6 = (~(Opoet6 & J0jxx6));
assign MEMATTRS[0] = (~(Gha6z6 & Oha6z6));
assign Oha6z6 = (~(Rj9ov6 & Gfqnv6));
assign Gfqnv6 = (~(Wha6z6 & Eia6z6));
assign Wha6z6 = (Mia6z6 | Uia6z6);
assign Mia6z6 = (Kja6z6 ? Cja6z6 : Cba6z6);
assign Cja6z6 = (~(Sja6z6 & Cba6z6));
assign Sja6z6 = (Aka6z6 & Ika6z6);
assign Gha6z6 = (~(Proet6 & J0jxx6));
assign JTAGNSW = (!Dz1nv6);
assign Dz1nv6 = (Qka6z6 | Fqxmz6[5]);
assign Qka6z6 = (Fqxmz6[4] & Yka6z6);
assign Yka6z6 = (~(Gla6z6 & Ola6z6));
assign Ola6z6 = (~(Fqxmz6[2] | Fqxmz6[3]));
assign Gla6z6 = (~(Fqxmz6[0] | Fqxmz6[1]));
assign HWRITES = (~(Wla6z6 & Ema6z6));
assign Ema6z6 = (~(Mma6z6 & L3bdt6));
assign Wla6z6 = (Uma6z6 & Cna6z6);
assign Cna6z6 = (~(J0jxx6 & Kna6z6));
assign Kna6z6 = (Qo8iy6 | Sna6z6);
assign Sna6z6 = (~(Kxixx6 | Xvgxx6));
assign Kxixx6 = (!I2yet6);
assign Uma6z6 = (~(Aoa6z6 & Lhmov6));
assign HWDATAS[9] = (~(Ioa6z6 & Qoa6z6));
assign Qoa6z6 = (~(Yoa6z6 & H5q7x6));
assign Ioa6z6 = (Gpa6z6 & Opa6z6);
assign Opa6z6 = (~(Wpa6z6 & Itb7z6[9]));
assign Gpa6z6 = (~(Tim7z6[9] & Eqa6z6));
assign HWDATAS[8] = (~(Mqa6z6 & Uqa6z6));
assign Uqa6z6 = (~(Yoa6z6 & Kqonv6));
assign Mqa6z6 = (Cra6z6 & Kra6z6);
assign Kra6z6 = (~(Wpa6z6 & Itb7z6[8]));
assign Cra6z6 = (~(Tim7z6[8] & Eqa6z6));
assign HWDATAS[7] = (~(Sra6z6 & Asa6z6));
assign Asa6z6 = (~(Yoa6z6 & Kwp7x6));
assign Sra6z6 = (Isa6z6 & Qsa6z6);
assign Qsa6z6 = (~(Wpa6z6 & Itb7z6[7]));
assign Isa6z6 = (~(Tim7z6[7] & Eqa6z6));
assign HWDATAS[6] = (~(Ysa6z6 & Gta6z6));
assign Gta6z6 = (~(Yoa6z6 & Lzq7x6));
assign Ysa6z6 = (Ota6z6 & Wta6z6);
assign Wta6z6 = (~(Wpa6z6 & Itb7z6[6]));
assign Ota6z6 = (~(Tim7z6[6] & Eqa6z6));
assign HWDATAS[5] = (~(Eua6z6 & Mua6z6));
assign Mua6z6 = (~(Yoa6z6 & Zsq7x6));
assign Eua6z6 = (Uua6z6 & Cva6z6);
assign Cva6z6 = (~(Wpa6z6 & Itb7z6[5]));
assign Uua6z6 = (~(Tim7z6[5] & Eqa6z6));
assign HWDATAS[4] = (~(Kva6z6 & Sva6z6));
assign Sva6z6 = (~(Yoa6z6 & Pnq7x6));
assign Kva6z6 = (Awa6z6 & Iwa6z6);
assign Iwa6z6 = (~(Wpa6z6 & Itb7z6[4]));
assign Awa6z6 = (~(Tim7z6[4] & Eqa6z6));
assign HWDATAS[3] = (~(Qwa6z6 & Ywa6z6));
assign Ywa6z6 = (~(Yoa6z6 & Fiq7x6));
assign Qwa6z6 = (Gxa6z6 & Oxa6z6);
assign Oxa6z6 = (~(Wpa6z6 & Itb7z6[3]));
assign Gxa6z6 = (~(Tim7z6[3] & Eqa6z6));
assign HWDATAS[31] = (~(Wxa6z6 & Eya6z6));
assign Eya6z6 = (~(Yoa6z6 & Ht1ov6));
assign Wxa6z6 = (Mya6z6 & Uya6z6);
assign Uya6z6 = (~(Wpa6z6 & Itb7z6[31]));
assign Mya6z6 = (~(Tim7z6[31] & Eqa6z6));
assign HWDATAS[30] = (~(Cza6z6 & Kza6z6));
assign Kza6z6 = (~(Yoa6z6 & Vxq7x6));
assign Cza6z6 = (Sza6z6 & A0b6z6);
assign A0b6z6 = (~(Wpa6z6 & Itb7z6[30]));
assign Sza6z6 = (~(Tim7z6[30] & Eqa6z6));
assign HWDATAS[2] = (~(I0b6z6 & Q0b6z6));
assign Q0b6z6 = (~(Yoa6z6 & Vcq7x6));
assign I0b6z6 = (Y0b6z6 & G1b6z6);
assign G1b6z6 = (~(Wpa6z6 & Itb7z6[2]));
assign Y0b6z6 = (~(Tim7z6[2] & Eqa6z6));
assign HWDATAS[29] = (~(O1b6z6 & W1b6z6));
assign W1b6z6 = (~(Yoa6z6 & Qrq7x6));
assign O1b6z6 = (E2b6z6 & M2b6z6);
assign M2b6z6 = (~(Wpa6z6 & Itb7z6[29]));
assign E2b6z6 = (~(Tim7z6[29] & Eqa6z6));
assign HWDATAS[28] = (~(U2b6z6 & C3b6z6));
assign C3b6z6 = (~(Yoa6z6 & Gmq7x6));
assign U2b6z6 = (K3b6z6 & S3b6z6);
assign S3b6z6 = (~(Wpa6z6 & Itb7z6[28]));
assign K3b6z6 = (~(Tim7z6[28] & Eqa6z6));
assign HWDATAS[27] = (~(A4b6z6 & I4b6z6));
assign I4b6z6 = (~(Yoa6z6 & Wgq7x6));
assign A4b6z6 = (Q4b6z6 & Y4b6z6);
assign Y4b6z6 = (~(Wpa6z6 & Itb7z6[27]));
assign Q4b6z6 = (~(Tim7z6[27] & Eqa6z6));
assign HWDATAS[26] = (~(G5b6z6 & O5b6z6));
assign O5b6z6 = (~(Yoa6z6 & Mbq7x6));
assign G5b6z6 = (W5b6z6 & E6b6z6);
assign E6b6z6 = (~(Wpa6z6 & Itb7z6[26]));
assign W5b6z6 = (~(Tim7z6[26] & Eqa6z6));
assign HWDATAS[25] = (~(M6b6z6 & U6b6z6));
assign U6b6z6 = (~(Yoa6z6 & C6q7x6));
assign M6b6z6 = (C7b6z6 & K7b6z6);
assign K7b6z6 = (~(Wpa6z6 & Itb7z6[25]));
assign C7b6z6 = (~(Tim7z6[25] & Eqa6z6));
assign HWDATAS[24] = (~(S7b6z6 & A8b6z6));
assign A8b6z6 = (~(Yoa6z6 & Yqonv6));
assign S7b6z6 = (I8b6z6 & Q8b6z6);
assign Q8b6z6 = (~(Wpa6z6 & Itb7z6[24]));
assign I8b6z6 = (~(Tim7z6[24] & Eqa6z6));
assign HWDATAS[23] = (~(Y8b6z6 & G9b6z6));
assign G9b6z6 = (~(Yoa6z6 & Xzp7x6));
assign Y8b6z6 = (O9b6z6 & W9b6z6);
assign W9b6z6 = (~(Wpa6z6 & Itb7z6[23]));
assign O9b6z6 = (~(Tim7z6[23] & Eqa6z6));
assign HWDATAS[22] = (~(Eab6z6 & Mab6z6));
assign Mab6z6 = (~(Yoa6z6 & Wuq7x6));
assign Eab6z6 = (Uab6z6 & Cbb6z6);
assign Cbb6z6 = (~(Wpa6z6 & Itb7z6[22]));
assign Uab6z6 = (~(Tim7z6[22] & Eqa6z6));
assign HWDATAS[21] = (~(Kbb6z6 & Sbb6z6));
assign Sbb6z6 = (~(Yoa6z6 & Mpq7x6));
assign Kbb6z6 = (Acb6z6 & Icb6z6);
assign Icb6z6 = (~(Wpa6z6 & Itb7z6[21]));
assign Acb6z6 = (~(Tim7z6[21] & Eqa6z6));
assign HWDATAS[20] = (~(Qcb6z6 & Ycb6z6));
assign Ycb6z6 = (~(Yoa6z6 & Ckq7x6));
assign Qcb6z6 = (Gdb6z6 & Odb6z6);
assign Odb6z6 = (~(Wpa6z6 & Itb7z6[20]));
assign Gdb6z6 = (~(Tim7z6[20] & Eqa6z6));
assign HWDATAS[1] = (~(Wdb6z6 & Eeb6z6));
assign Eeb6z6 = (~(Yoa6z6 & L7q7x6));
assign Wdb6z6 = (Meb6z6 & Ueb6z6);
assign Ueb6z6 = (~(Wpa6z6 & Itb7z6[1]));
assign Meb6z6 = (~(Tim7z6[1] & Eqa6z6));
assign HWDATAS[19] = (~(Cfb6z6 & Kfb6z6));
assign Kfb6z6 = (~(Yoa6z6 & Seq7x6));
assign Cfb6z6 = (Sfb6z6 & Agb6z6);
assign Agb6z6 = (~(Wpa6z6 & Itb7z6[19]));
assign Sfb6z6 = (~(Tim7z6[19] & Eqa6z6));
assign HWDATAS[18] = (~(Igb6z6 & Qgb6z6));
assign Qgb6z6 = (~(Yoa6z6 & I9q7x6));
assign Igb6z6 = (Ygb6z6 & Ghb6z6);
assign Ghb6z6 = (~(Wpa6z6 & Itb7z6[18]));
assign Ygb6z6 = (~(Tim7z6[18] & Eqa6z6));
assign HWDATAS[17] = (~(Ohb6z6 & Whb6z6));
assign Whb6z6 = (~(Yoa6z6 & Y3q7x6));
assign Ohb6z6 = (Eib6z6 & Mib6z6);
assign Mib6z6 = (~(Wpa6z6 & Itb7z6[17]));
assign Eib6z6 = (~(Tim7z6[17] & Eqa6z6));
assign HWDATAS[16] = (~(Uib6z6 & Cjb6z6));
assign Cjb6z6 = (~(Yoa6z6 & V4r7x6));
assign Uib6z6 = (Kjb6z6 & Sjb6z6);
assign Sjb6z6 = (~(Wpa6z6 & Itb7z6[16]));
assign Kjb6z6 = (~(Tim7z6[16] & Eqa6z6));
assign HWDATAS[15] = (~(Akb6z6 & Ikb6z6));
assign Ikb6z6 = (~(Yoa6z6 & Oyp7x6));
assign Akb6z6 = (Qkb6z6 & Ykb6z6);
assign Ykb6z6 = (~(Wpa6z6 & Itb7z6[15]));
assign Qkb6z6 = (~(Tim7z6[15] & Eqa6z6));
assign HWDATAS[14] = (~(Glb6z6 & Olb6z6));
assign Olb6z6 = (~(Yoa6z6 & Twq7x6));
assign Glb6z6 = (Wlb6z6 & Emb6z6);
assign Emb6z6 = (~(Wpa6z6 & Itb7z6[14]));
assign Wlb6z6 = (~(Tim7z6[14] & Eqa6z6));
assign HWDATAS[13] = (~(Mmb6z6 & Umb6z6));
assign Umb6z6 = (~(Yoa6z6 & Vqq7x6));
assign Mmb6z6 = (Cnb6z6 & Knb6z6);
assign Knb6z6 = (~(Wpa6z6 & Itb7z6[13]));
assign Cnb6z6 = (~(Tim7z6[13] & Eqa6z6));
assign HWDATAS[12] = (~(Snb6z6 & Aob6z6));
assign Aob6z6 = (~(Yoa6z6 & Llq7x6));
assign Snb6z6 = (Iob6z6 & Qob6z6);
assign Qob6z6 = (~(Wpa6z6 & Itb7z6[12]));
assign Iob6z6 = (~(Tim7z6[12] & Eqa6z6));
assign HWDATAS[11] = (~(Yob6z6 & Gpb6z6));
assign Gpb6z6 = (~(Yoa6z6 & Bgq7x6));
assign Yob6z6 = (Opb6z6 & Wpb6z6);
assign Wpb6z6 = (~(Wpa6z6 & Itb7z6[11]));
assign Opb6z6 = (~(Tim7z6[11] & Eqa6z6));
assign HWDATAS[10] = (~(Eqb6z6 & Mqb6z6));
assign Mqb6z6 = (~(Yoa6z6 & Raq7x6));
assign Eqb6z6 = (Uqb6z6 & Crb6z6);
assign Crb6z6 = (~(Wpa6z6 & Itb7z6[10]));
assign Uqb6z6 = (~(Tim7z6[10] & Eqa6z6));
assign HWDATAS[0] = (~(Krb6z6 & Srb6z6));
assign Srb6z6 = (~(Yoa6z6 & I8r7x6));
assign Yoa6z6 = (Svn7z6[0] & Asb6z6);
assign Krb6z6 = (Isb6z6 & Qsb6z6);
assign Qsb6z6 = (~(Wpa6z6 & Itb7z6[0]));
assign Wpa6z6 = (Svn7z6[1] & Asb6z6);
assign Isb6z6 = (~(Tim7z6[0] & Eqa6z6));
assign Eqa6z6 = (~(P3jxx6 & Asb6z6));
assign Asb6z6 = (~(Sb0jy6 & Qln7z6[1]));
assign P3jxx6 = (!Svn7z6[2]);
assign HWDATAD[9] = (~(Ysb6z6 & Gtb6z6));
assign Gtb6z6 = (~(Tim7z6[9] & Otb6z6));
assign Ysb6z6 = (Wtb6z6 & Eub6z6);
assign Eub6z6 = (~(Mub6z6 & H5q7x6));
assign H5q7x6 = (!Uub6z6);
assign Uub6z6 = (No7et6 ? Kvb6z6 : Cvb6z6);
assign Wtb6z6 = (~(Svb6z6 & Itb7z6[9]));
assign HWDATAD[8] = (~(Awb6z6 & Iwb6z6));
assign Iwb6z6 = (~(Tim7z6[8] & Otb6z6));
assign Awb6z6 = (Qwb6z6 & Ywb6z6);
assign Ywb6z6 = (~(Mub6z6 & Kqonv6));
assign Kqonv6 = (!Gxb6z6);
assign Gxb6z6 = (No7et6 ? Wxb6z6 : Oxb6z6);
assign Qwb6z6 = (~(Svb6z6 & Itb7z6[8]));
assign HWDATAD[7] = (~(Eyb6z6 & Myb6z6));
assign Myb6z6 = (~(Tim7z6[7] & Otb6z6));
assign Eyb6z6 = (Uyb6z6 & Czb6z6);
assign Czb6z6 = (~(Mub6z6 & Kwp7x6));
assign Kwp7x6 = (!Kzb6z6);
assign Kzb6z6 = (No7et6 ? A0c6z6 : Szb6z6);
assign Uyb6z6 = (~(Svb6z6 & Itb7z6[7]));
assign HWDATAD[6] = (~(I0c6z6 & Q0c6z6));
assign Q0c6z6 = (~(Tim7z6[6] & Otb6z6));
assign I0c6z6 = (Y0c6z6 & G1c6z6);
assign G1c6z6 = (~(Mub6z6 & Lzq7x6));
assign Lzq7x6 = (!O1c6z6);
assign O1c6z6 = (No7et6 ? E2c6z6 : W1c6z6);
assign Y0c6z6 = (~(Svb6z6 & Itb7z6[6]));
assign HWDATAD[5] = (~(M2c6z6 & U2c6z6));
assign U2c6z6 = (~(Tim7z6[5] & Otb6z6));
assign M2c6z6 = (C3c6z6 & K3c6z6);
assign K3c6z6 = (~(Mub6z6 & Zsq7x6));
assign Zsq7x6 = (!S3c6z6);
assign S3c6z6 = (No7et6 ? I4c6z6 : A4c6z6);
assign C3c6z6 = (~(Svb6z6 & Itb7z6[5]));
assign HWDATAD[4] = (~(Q4c6z6 & Y4c6z6));
assign Y4c6z6 = (~(Tim7z6[4] & Otb6z6));
assign Q4c6z6 = (G5c6z6 & O5c6z6);
assign O5c6z6 = (~(Mub6z6 & Pnq7x6));
assign Pnq7x6 = (!W5c6z6);
assign W5c6z6 = (No7et6 ? M6c6z6 : E6c6z6);
assign G5c6z6 = (~(Svb6z6 & Itb7z6[4]));
assign HWDATAD[3] = (~(U6c6z6 & C7c6z6));
assign C7c6z6 = (~(Tim7z6[3] & Otb6z6));
assign U6c6z6 = (K7c6z6 & S7c6z6);
assign S7c6z6 = (~(Mub6z6 & Fiq7x6));
assign Fiq7x6 = (!A8c6z6);
assign A8c6z6 = (No7et6 ? Q8c6z6 : I8c6z6);
assign K7c6z6 = (~(Svb6z6 & Itb7z6[3]));
assign HWDATAD[31] = (~(Y8c6z6 & G9c6z6));
assign G9c6z6 = (~(Tim7z6[31] & Otb6z6));
assign Y8c6z6 = (O9c6z6 & W9c6z6);
assign W9c6z6 = (~(Mub6z6 & Ht1ov6));
assign Ht1ov6 = (!Eac6z6);
assign Eac6z6 = (No7et6 ? Szb6z6 : A0c6z6);
assign Szb6z6 = (Mac6z6 & Uac6z6);
assign Uac6z6 = (Cbc6z6 & Kbc6z6);
assign Kbc6z6 = (~(Sbc6z6 & Acc6z6));
assign Cbc6z6 = (Icc6z6 & Qcc6z6);
assign Qcc6z6 = (~(Ddo6x6 & Ycc6z6));
assign Ddo6x6 = (Nob7z6[7] & Rslov6);
assign Icc6z6 = (~(Gdc6z6 & Odc6z6));
assign Mac6z6 = (Wdc6z6 & Eec6z6);
assign Eec6z6 = (~(Kxb7z6[7] & Mec6z6));
assign Wdc6z6 = (Uec6z6 & Cfc6z6);
assign Cfc6z6 = (~(Kfc6z6 & Sfc6z6));
assign Uec6z6 = (~(Agc6z6 & Igc6z6));
assign A0c6z6 = (Qgc6z6 & Ygc6z6);
assign Ygc6z6 = (Ghc6z6 & Ohc6z6);
assign Ohc6z6 = (~(Whc6z6 & Sfc6z6));
assign Ghc6z6 = (Eic6z6 & Mic6z6);
assign Mic6z6 = (~(Uic6z6 & Odc6z6));
assign Eic6z6 = (~(Cjc6z6 & Acc6z6));
assign Qgc6z6 = (Kjc6z6 & Sjc6z6);
assign Sjc6z6 = (~(O4gdt6 & Ycc6z6));
assign Kjc6z6 = (Akc6z6 & Ikc6z6);
assign Ikc6z6 = (~(Gdc6z6 & Igc6z6));
assign Akc6z6 = (~(Kxb7z6[31] & Mec6z6));
assign O9c6z6 = (~(Svb6z6 & Itb7z6[31]));
assign HWDATAD[30] = (~(Qkc6z6 & Ykc6z6));
assign Ykc6z6 = (~(Tim7z6[30] & Otb6z6));
assign Qkc6z6 = (Glc6z6 & Olc6z6);
assign Olc6z6 = (~(Mub6z6 & Vxq7x6));
assign Vxq7x6 = (!Wlc6z6);
assign Wlc6z6 = (No7et6 ? W1c6z6 : E2c6z6);
assign W1c6z6 = (Emc6z6 & Mmc6z6);
assign Mmc6z6 = (Umc6z6 & Cnc6z6);
assign Cnc6z6 = (~(Sbc6z6 & Knc6z6));
assign Umc6z6 = (Snc6z6 & Aoc6z6);
assign Aoc6z6 = (~(Nob7z6[6] & Ioc6z6));
assign Snc6z6 = (~(Gdc6z6 & Qoc6z6));
assign Emc6z6 = (Yoc6z6 & Gpc6z6);
assign Gpc6z6 = (~(Kxb7z6[6] & Mec6z6));
assign Yoc6z6 = (Opc6z6 & Wpc6z6);
assign Wpc6z6 = (~(Kfc6z6 & Eqc6z6));
assign Opc6z6 = (~(Agc6z6 & Mqc6z6));
assign E2c6z6 = (Uqc6z6 & Crc6z6);
assign Crc6z6 = (Krc6z6 & Src6z6);
assign Src6z6 = (~(Whc6z6 & Eqc6z6));
assign Krc6z6 = (Asc6z6 & Isc6z6);
assign Isc6z6 = (~(Uic6z6 & Qoc6z6));
assign Asc6z6 = (~(Cjc6z6 & Knc6z6));
assign Uqc6z6 = (Qsc6z6 & Ysc6z6);
assign Ysc6z6 = (~(D6gdt6 & Ycc6z6));
assign Qsc6z6 = (Gtc6z6 & Otc6z6);
assign Otc6z6 = (~(Gdc6z6 & Mqc6z6));
assign Gtc6z6 = (~(Kxb7z6[30] & Mec6z6));
assign Glc6z6 = (~(Svb6z6 & Itb7z6[30]));
assign HWDATAD[2] = (~(Wtc6z6 & Euc6z6));
assign Euc6z6 = (~(Tim7z6[2] & Otb6z6));
assign Wtc6z6 = (Muc6z6 & Uuc6z6);
assign Uuc6z6 = (~(Mub6z6 & Vcq7x6));
assign Vcq7x6 = (!Cvc6z6);
assign Cvc6z6 = (No7et6 ? Svc6z6 : Kvc6z6);
assign Muc6z6 = (~(Svb6z6 & Itb7z6[2]));
assign HWDATAD[29] = (~(Awc6z6 & Iwc6z6));
assign Iwc6z6 = (~(Tim7z6[29] & Otb6z6));
assign Awc6z6 = (Qwc6z6 & Ywc6z6);
assign Ywc6z6 = (~(Mub6z6 & Qrq7x6));
assign Qrq7x6 = (!Gxc6z6);
assign Gxc6z6 = (No7et6 ? A4c6z6 : I4c6z6);
assign A4c6z6 = (Oxc6z6 & Wxc6z6);
assign Wxc6z6 = (Eyc6z6 & Myc6z6);
assign Myc6z6 = (~(Sbc6z6 & Uyc6z6));
assign Eyc6z6 = (Czc6z6 & Kzc6z6);
assign Kzc6z6 = (~(Jti6x6 & Ycc6z6));
assign Jti6x6 = (Nob7z6[5] & Rslov6);
assign Czc6z6 = (~(Gdc6z6 & Szc6z6));
assign Oxc6z6 = (A0d6z6 & I0d6z6);
assign I0d6z6 = (~(Kxb7z6[5] & Mec6z6));
assign A0d6z6 = (Q0d6z6 & Y0d6z6);
assign Y0d6z6 = (~(Kfc6z6 & G1d6z6));
assign Q0d6z6 = (~(Agc6z6 & O1d6z6));
assign I4c6z6 = (W1d6z6 & E2d6z6);
assign E2d6z6 = (M2d6z6 & U2d6z6);
assign U2d6z6 = (~(Whc6z6 & G1d6z6));
assign M2d6z6 = (C3d6z6 & K3d6z6);
assign K3d6z6 = (~(Uic6z6 & Szc6z6));
assign C3d6z6 = (~(Cjc6z6 & Uyc6z6));
assign W1d6z6 = (S3d6z6 & A4d6z6);
assign A4d6z6 = (~(S7gdt6 & Ycc6z6));
assign S3d6z6 = (I4d6z6 & Q4d6z6);
assign Q4d6z6 = (~(Gdc6z6 & O1d6z6));
assign I4d6z6 = (~(Kxb7z6[29] & Mec6z6));
assign Qwc6z6 = (~(Svb6z6 & Itb7z6[29]));
assign HWDATAD[28] = (~(Y4d6z6 & G5d6z6));
assign G5d6z6 = (~(Tim7z6[28] & Otb6z6));
assign Y4d6z6 = (O5d6z6 & W5d6z6);
assign W5d6z6 = (~(Mub6z6 & Gmq7x6));
assign Gmq7x6 = (!E6d6z6);
assign E6d6z6 = (No7et6 ? E6c6z6 : M6c6z6);
assign E6c6z6 = (M6d6z6 & U6d6z6);
assign U6d6z6 = (C7d6z6 & K7d6z6);
assign K7d6z6 = (~(Sbc6z6 & S7d6z6));
assign C7d6z6 = (A8d6z6 & I8d6z6);
assign I8d6z6 = (~(Nob7z6[4] & Ioc6z6));
assign A8d6z6 = (~(Gdc6z6 & Q8d6z6));
assign M6d6z6 = (Y8d6z6 & G9d6z6);
assign G9d6z6 = (~(Kxb7z6[4] & Mec6z6));
assign Y8d6z6 = (O9d6z6 & W9d6z6);
assign W9d6z6 = (~(Kfc6z6 & Ead6z6));
assign O9d6z6 = (~(Agc6z6 & Mad6z6));
assign M6c6z6 = (Uad6z6 & Cbd6z6);
assign Cbd6z6 = (Kbd6z6 & Sbd6z6);
assign Sbd6z6 = (~(Whc6z6 & Ead6z6));
assign Kbd6z6 = (Acd6z6 & Icd6z6);
assign Icd6z6 = (~(Uic6z6 & Q8d6z6));
assign Acd6z6 = (~(Cjc6z6 & S7d6z6));
assign Uad6z6 = (Qcd6z6 & Ycd6z6);
assign Ycd6z6 = (~(H9gdt6 & Ycc6z6));
assign Qcd6z6 = (Gdd6z6 & Odd6z6);
assign Odd6z6 = (~(Gdc6z6 & Mad6z6));
assign Gdd6z6 = (~(Kxb7z6[28] & Mec6z6));
assign O5d6z6 = (~(Svb6z6 & Itb7z6[28]));
assign HWDATAD[27] = (~(Wdd6z6 & Eed6z6));
assign Eed6z6 = (~(Tim7z6[27] & Otb6z6));
assign Wdd6z6 = (Med6z6 & Ued6z6);
assign Ued6z6 = (~(Mub6z6 & Wgq7x6));
assign Wgq7x6 = (!Cfd6z6);
assign Cfd6z6 = (No7et6 ? I8c6z6 : Q8c6z6);
assign I8c6z6 = (Kfd6z6 & Sfd6z6);
assign Sfd6z6 = (Agd6z6 & Igd6z6);
assign Igd6z6 = (~(Sbc6z6 & Qgd6z6));
assign Agd6z6 = (Ygd6z6 & Ghd6z6);
assign Ghd6z6 = (~(Nob7z6[3] & Ioc6z6));
assign Ygd6z6 = (~(Gdc6z6 & Ohd6z6));
assign Kfd6z6 = (Whd6z6 & Eid6z6);
assign Eid6z6 = (~(Kxb7z6[3] & Mec6z6));
assign Whd6z6 = (Mid6z6 & Uid6z6);
assign Uid6z6 = (~(Kfc6z6 & Cjd6z6));
assign Mid6z6 = (~(Agc6z6 & Kjd6z6));
assign Q8c6z6 = (Sjd6z6 & Akd6z6);
assign Akd6z6 = (Ikd6z6 & Qkd6z6);
assign Qkd6z6 = (~(Whc6z6 & Cjd6z6));
assign Ikd6z6 = (Ykd6z6 & Gld6z6);
assign Gld6z6 = (~(Uic6z6 & Ohd6z6));
assign Ykd6z6 = (~(Cjc6z6 & Qgd6z6));
assign Sjd6z6 = (Old6z6 & Wld6z6);
assign Wld6z6 = (~(Lsfdt6 & Ycc6z6));
assign Old6z6 = (Emd6z6 & Mmd6z6);
assign Mmd6z6 = (~(Gdc6z6 & Kjd6z6));
assign Emd6z6 = (~(Kxb7z6[27] & Mec6z6));
assign Med6z6 = (~(Svb6z6 & Itb7z6[27]));
assign HWDATAD[26] = (~(Umd6z6 & Cnd6z6));
assign Cnd6z6 = (~(Tim7z6[26] & Otb6z6));
assign Umd6z6 = (Knd6z6 & Snd6z6);
assign Snd6z6 = (~(Mub6z6 & Mbq7x6));
assign Mbq7x6 = (!Aod6z6);
assign Aod6z6 = (No7et6 ? Kvc6z6 : Svc6z6);
assign Kvc6z6 = (Iod6z6 & Qod6z6);
assign Qod6z6 = (Yod6z6 & Gpd6z6);
assign Gpd6z6 = (~(Sbc6z6 & Opd6z6));
assign Yod6z6 = (Wpd6z6 & Eqd6z6);
assign Eqd6z6 = (~(Tx1jw6 & Ycc6z6));
assign Tx1jw6 = (Nob7z6[2] & Rslov6);
assign Wpd6z6 = (~(Gdc6z6 & Mqd6z6));
assign Iod6z6 = (Uqd6z6 & Crd6z6);
assign Crd6z6 = (~(Kxb7z6[2] & Mec6z6));
assign Uqd6z6 = (Krd6z6 & Srd6z6);
assign Srd6z6 = (~(Kfc6z6 & Asd6z6));
assign Krd6z6 = (~(Agc6z6 & Isd6z6));
assign Svc6z6 = (Qsd6z6 & Ysd6z6);
assign Ysd6z6 = (Gtd6z6 & Otd6z6);
assign Otd6z6 = (~(Cjc6z6 & Opd6z6));
assign Gtd6z6 = (Wtd6z6 & Eud6z6);
assign Eud6z6 = (Mud6z6 | Uud6z6);
assign Wtd6z6 = (~(Uic6z6 & Mqd6z6));
assign Qsd6z6 = (Cvd6z6 & Kvd6z6);
assign Kvd6z6 = (~(Kxb7z6[26] & Mec6z6));
assign Cvd6z6 = (Svd6z6 & Awd6z6);
assign Awd6z6 = (~(Whc6z6 & Asd6z6));
assign Svd6z6 = (~(Gdc6z6 & Isd6z6));
assign Knd6z6 = (~(Svb6z6 & Itb7z6[26]));
assign HWDATAD[25] = (~(Iwd6z6 & Qwd6z6));
assign Qwd6z6 = (~(Tim7z6[25] & Otb6z6));
assign Iwd6z6 = (Ywd6z6 & Gxd6z6);
assign Gxd6z6 = (~(Mub6z6 & C6q7x6));
assign C6q7x6 = (!Oxd6z6);
assign Oxd6z6 = (No7et6 ? Eyd6z6 : Wxd6z6);
assign Ywd6z6 = (~(Svb6z6 & Itb7z6[25]));
assign HWDATAD[24] = (~(Myd6z6 & Uyd6z6));
assign Uyd6z6 = (~(Tim7z6[24] & Otb6z6));
assign Myd6z6 = (Czd6z6 & Kzd6z6);
assign Kzd6z6 = (~(Mub6z6 & Yqonv6));
assign Yqonv6 = (!Szd6z6);
assign Szd6z6 = (No7et6 ? I0e6z6 : A0e6z6);
assign Czd6z6 = (~(Svb6z6 & Itb7z6[24]));
assign HWDATAD[23] = (~(Q0e6z6 & Y0e6z6));
assign Y0e6z6 = (~(Tim7z6[23] & Otb6z6));
assign Q0e6z6 = (G1e6z6 & O1e6z6);
assign O1e6z6 = (~(Mub6z6 & Xzp7x6));
assign Xzp7x6 = (!W1e6z6);
assign W1e6z6 = (No7et6 ? M2e6z6 : E2e6z6);
assign G1e6z6 = (~(Svb6z6 & Itb7z6[23]));
assign HWDATAD[22] = (~(U2e6z6 & C3e6z6));
assign C3e6z6 = (~(Tim7z6[22] & Otb6z6));
assign U2e6z6 = (K3e6z6 & S3e6z6);
assign S3e6z6 = (~(Mub6z6 & Wuq7x6));
assign Wuq7x6 = (!A4e6z6);
assign A4e6z6 = (No7et6 ? Q4e6z6 : I4e6z6);
assign K3e6z6 = (~(Svb6z6 & Itb7z6[22]));
assign HWDATAD[21] = (~(Y4e6z6 & G5e6z6));
assign G5e6z6 = (~(Tim7z6[21] & Otb6z6));
assign Y4e6z6 = (O5e6z6 & W5e6z6);
assign W5e6z6 = (~(Mub6z6 & Mpq7x6));
assign Mpq7x6 = (!E6e6z6);
assign E6e6z6 = (No7et6 ? U6e6z6 : M6e6z6);
assign O5e6z6 = (~(Svb6z6 & Itb7z6[21]));
assign HWDATAD[20] = (~(C7e6z6 & K7e6z6));
assign K7e6z6 = (~(Tim7z6[20] & Otb6z6));
assign C7e6z6 = (S7e6z6 & A8e6z6);
assign A8e6z6 = (~(Mub6z6 & Ckq7x6));
assign Ckq7x6 = (!I8e6z6);
assign I8e6z6 = (No7et6 ? Y8e6z6 : Q8e6z6);
assign S7e6z6 = (~(Svb6z6 & Itb7z6[20]));
assign HWDATAD[1] = (~(G9e6z6 & O9e6z6));
assign O9e6z6 = (~(Tim7z6[1] & Otb6z6));
assign G9e6z6 = (W9e6z6 & Eae6z6);
assign Eae6z6 = (~(Mub6z6 & L7q7x6));
assign L7q7x6 = (!Mae6z6);
assign Mae6z6 = (No7et6 ? Wxd6z6 : Eyd6z6);
assign Wxd6z6 = (Uae6z6 & Cbe6z6);
assign Cbe6z6 = (Kbe6z6 & Sbe6z6);
assign Sbe6z6 = (Ace6z6 & Ice6z6);
assign Ice6z6 = (~(Qce6z6 & Ycc6z6));
assign Qce6z6 = (~(Yce6z6 & Gde6z6));
assign Gde6z6 = (~(Ohe7z6[2] & Ode6z6));
assign Ace6z6 = (~(Uic6z6 & Wde6z6));
assign Kbe6z6 = (Eee6z6 & Mee6z6);
assign Mee6z6 = (~(Cjc6z6 & Uee6z6));
assign Eee6z6 = (~(Whc6z6 & Cfe6z6));
assign Uae6z6 = (Kfe6z6 & Sfe6z6);
assign Sfe6z6 = (~(Jjbdt6 & Age6z6));
assign Kfe6z6 = (Ige6z6 & Qge6z6);
assign Qge6z6 = (~(Gdc6z6 & Yge6z6));
assign Ige6z6 = (~(Kxb7z6[25] & Mec6z6));
assign Eyd6z6 = (Ghe6z6 & Ohe6z6);
assign Ohe6z6 = (Whe6z6 & Eie6z6);
assign Eie6z6 = (~(Sbc6z6 & Uee6z6));
assign Whe6z6 = (Mie6z6 & Uie6z6);
assign Uie6z6 = (~(Nob7z6[1] & Ioc6z6));
assign Mie6z6 = (~(Gdc6z6 & Wde6z6));
assign Ghe6z6 = (Cje6z6 & Kje6z6);
assign Kje6z6 = (~(Kxb7z6[1] & Mec6z6));
assign Cje6z6 = (Sje6z6 & Ake6z6);
assign Ake6z6 = (~(Kfc6z6 & Cfe6z6));
assign Sje6z6 = (~(Agc6z6 & Yge6z6));
assign W9e6z6 = (~(Svb6z6 & Itb7z6[1]));
assign HWDATAD[19] = (~(Ike6z6 & Qke6z6));
assign Qke6z6 = (~(Tim7z6[19] & Otb6z6));
assign Ike6z6 = (Yke6z6 & Gle6z6);
assign Gle6z6 = (~(Mub6z6 & Seq7x6));
assign Seq7x6 = (!Ole6z6);
assign Ole6z6 = (No7et6 ? Eme6z6 : Wle6z6);
assign Yke6z6 = (~(Svb6z6 & Itb7z6[19]));
assign HWDATAD[18] = (~(Mme6z6 & Ume6z6));
assign Ume6z6 = (~(Tim7z6[18] & Otb6z6));
assign Mme6z6 = (Cne6z6 & Kne6z6);
assign Kne6z6 = (~(Mub6z6 & I9q7x6));
assign I9q7x6 = (!Sne6z6);
assign Sne6z6 = (No7et6 ? Ioe6z6 : Aoe6z6);
assign Cne6z6 = (~(Svb6z6 & Itb7z6[18]));
assign HWDATAD[17] = (~(Qoe6z6 & Yoe6z6));
assign Yoe6z6 = (~(Tim7z6[17] & Otb6z6));
assign Qoe6z6 = (Gpe6z6 & Ope6z6);
assign Ope6z6 = (~(Mub6z6 & Y3q7x6));
assign Y3q7x6 = (!Wpe6z6);
assign Wpe6z6 = (No7et6 ? Cvb6z6 : Kvb6z6);
assign Cvb6z6 = (Eqe6z6 & Mqe6z6);
assign Mqe6z6 = (Uqe6z6 & Cre6z6);
assign Cre6z6 = (~(Kre6z6 & Uee6z6));
assign Uqe6z6 = (Sre6z6 & Ase6z6);
assign Ase6z6 = (~(Ise6z6 & Ycc6z6));
assign Ise6z6 = (Hfliw6 | Ir7et6);
assign Hfliw6 = (~(R9h7v6 & Qse6z6));
assign Qse6z6 = (~(Ku7et6 & U28et6));
assign Sre6z6 = (~(Agc6z6 & Wde6z6));
assign Eqe6z6 = (Yse6z6 & Gte6z6);
assign Gte6z6 = (~(Kxb7z6[9] & Mec6z6));
assign Yse6z6 = (Ote6z6 & Wte6z6);
assign Wte6z6 = (~(Eue6z6 & Cfe6z6));
assign Ote6z6 = (~(Mue6z6 & Yge6z6));
assign Kvb6z6 = (Uue6z6 & Cve6z6);
assign Cve6z6 = (Kve6z6 & Sve6z6);
assign Sve6z6 = (~(Awe6z6 & Cfe6z6));
assign Cfe6z6 = (~(Iwe6z6 & Qwe6z6));
assign Qwe6z6 = (~(Fhc7z6[9] & Ywe6z6));
assign Iwe6z6 = (Gxe6z6 & Oxe6z6);
assign Oxe6z6 = (~(Kxb7z6[9] & Wxe6z6));
assign Gxe6z6 = (~(Fth7z6[9] & Eye6z6));
assign Kve6z6 = (Mye6z6 & Uye6z6);
assign Uye6z6 = (~(Mue6z6 & Wde6z6));
assign Wde6z6 = (~(Cze6z6 & Kze6z6));
assign Kze6z6 = (~(Fhc7z6[25] & Ywe6z6));
assign Cze6z6 = (Sze6z6 & A0f6z6);
assign A0f6z6 = (~(Kxb7z6[25] & Wxe6z6));
assign Sze6z6 = (~(Fth7z6[25] & Eye6z6));
assign Mye6z6 = (~(I0f6z6 & Uee6z6));
assign Uee6z6 = (~(Q0f6z6 & Y0f6z6));
assign Y0f6z6 = (~(Kxb7z6[1] & Wxe6z6));
assign Q0f6z6 = (G1f6z6 & O1f6z6);
assign O1f6z6 = (~(E3c7z6[1] & Ywe6z6));
assign G1f6z6 = (~(Fth7z6[1] & Eye6z6));
assign Uue6z6 = (W1f6z6 & E2f6z6);
assign E2f6z6 = (~(Uic6z6 & Yge6z6));
assign Yge6z6 = (~(M2f6z6 & U2f6z6));
assign U2f6z6 = (~(Fhc7z6[17] & Ywe6z6));
assign M2f6z6 = (C3f6z6 & K3f6z6);
assign K3f6z6 = (~(Kxb7z6[17] & Wxe6z6));
assign C3f6z6 = (~(Fth7z6[17] & Eye6z6));
assign W1f6z6 = (~(Kxb7z6[17] & Mec6z6));
assign Gpe6z6 = (~(Svb6z6 & Itb7z6[17]));
assign HWDATAD[16] = (~(S3f6z6 & A4f6z6));
assign A4f6z6 = (~(Tim7z6[16] & Otb6z6));
assign S3f6z6 = (I4f6z6 & Q4f6z6);
assign Q4f6z6 = (~(Mub6z6 & V4r7x6));
assign V4r7x6 = (!Y4f6z6);
assign Y4f6z6 = (No7et6 ? Oxb6z6 : Wxb6z6);
assign Oxb6z6 = (G5f6z6 & O5f6z6);
assign O5f6z6 = (W5f6z6 & E6f6z6);
assign E6f6z6 = (~(Eue6z6 & M6f6z6));
assign W5f6z6 = (U6f6z6 & C7f6z6);
assign C7f6z6 = (~(Nob7z6[8] & Ioc6z6));
assign Ioc6z6 = (~(Uud6z6 | J2cdt6));
assign U6f6z6 = (~(Kre6z6 & K7f6z6));
assign G5f6z6 = (S7f6z6 & A8f6z6);
assign A8f6z6 = (~(Kxb7z6[8] & Mec6z6));
assign S7f6z6 = (I8f6z6 & Q8f6z6);
assign Q8f6z6 = (~(Mue6z6 & Y8f6z6));
assign I8f6z6 = (~(Agc6z6 & G9f6z6));
assign Wxb6z6 = (O9f6z6 & W9f6z6);
assign W9f6z6 = (Eaf6z6 & Maf6z6);
assign Maf6z6 = (~(Awe6z6 & M6f6z6));
assign Eaf6z6 = (Uaf6z6 & Cbf6z6);
assign Cbf6z6 = (~(Mue6z6 & G9f6z6));
assign Uaf6z6 = (~(I0f6z6 & K7f6z6));
assign O9f6z6 = (Kbf6z6 & Sbf6z6);
assign Sbf6z6 = (~(Inadt6 & Age6z6));
assign Kbf6z6 = (Acf6z6 & Icf6z6);
assign Icf6z6 = (~(Uic6z6 & Y8f6z6));
assign Acf6z6 = (~(Kxb7z6[16] & Mec6z6));
assign I4f6z6 = (~(Svb6z6 & Itb7z6[16]));
assign HWDATAD[15] = (~(Qcf6z6 & Ycf6z6));
assign Ycf6z6 = (~(Tim7z6[15] & Otb6z6));
assign Qcf6z6 = (Gdf6z6 & Odf6z6);
assign Odf6z6 = (~(Mub6z6 & Oyp7x6));
assign Oyp7x6 = (!Wdf6z6);
assign Wdf6z6 = (No7et6 ? E2e6z6 : M2e6z6);
assign E2e6z6 = (Eef6z6 & Mef6z6);
assign Mef6z6 = (Uef6z6 & Cff6z6);
assign Cff6z6 = (~(Awe6z6 & Sfc6z6));
assign Uef6z6 = (Kff6z6 & Sff6z6);
assign Sff6z6 = (~(Mue6z6 & Odc6z6));
assign Kff6z6 = (~(I0f6z6 & Acc6z6));
assign Eef6z6 = (Agf6z6 & Igf6z6);
assign Igf6z6 = (~(Uic6z6 & Igc6z6));
assign Agf6z6 = (~(Kxb7z6[23] & Mec6z6));
assign M2e6z6 = (Qgf6z6 & Ygf6z6);
assign Ygf6z6 = (Ghf6z6 & Ohf6z6);
assign Ohf6z6 = (Whf6z6 & Eif6z6);
assign Eif6z6 = (~(Mif6z6 & Mzmov6));
assign Mzmov6 = (~(Uif6z6 & Cjf6z6));
assign Cjf6z6 = (~(Ohe7z6[7] & Kjf6z6));
assign Uif6z6 = (~(Mfe7z6[7] & Ode6z6));
assign Whf6z6 = (~(Agc6z6 & Odc6z6));
assign Odc6z6 = (~(Sjf6z6 & Akf6z6));
assign Akf6z6 = (~(Fhc7z6[31] & Ywe6z6));
assign Sjf6z6 = (Ikf6z6 & Qkf6z6);
assign Qkf6z6 = (~(Kxb7z6[31] & Wxe6z6));
assign Ikf6z6 = (~(Fth7z6[31] & Eye6z6));
assign Ghf6z6 = (Ykf6z6 & Glf6z6);
assign Glf6z6 = (~(Kre6z6 & Acc6z6));
assign Acc6z6 = (~(Olf6z6 & Wlf6z6));
assign Wlf6z6 = (~(Fhc7z6[7] & Ywe6z6));
assign Olf6z6 = (Emf6z6 & Mmf6z6);
assign Mmf6z6 = (~(Kxb7z6[7] & Wxe6z6));
assign Emf6z6 = (~(Fth7z6[7] & Eye6z6));
assign Ykf6z6 = (~(Eue6z6 & Sfc6z6));
assign Sfc6z6 = (~(Umf6z6 & Cnf6z6));
assign Cnf6z6 = (~(Kxb7z6[15] & Wxe6z6));
assign Umf6z6 = (Knf6z6 & Snf6z6);
assign Snf6z6 = (~(Fth7z6[15] & Eye6z6));
assign Knf6z6 = (~(Fhc7z6[15] & Ywe6z6));
assign Qgf6z6 = (Aof6z6 & Iof6z6);
assign Iof6z6 = (Qof6z6 & Yof6z6);
assign Yof6z6 = (~(Mue6z6 & Igc6z6));
assign Igc6z6 = (~(Gpf6z6 & Opf6z6));
assign Opf6z6 = (~(Fhc7z6[23] & Ywe6z6));
assign Gpf6z6 = (Wpf6z6 & Eqf6z6);
assign Eqf6z6 = (~(Kxb7z6[23] & Wxe6z6));
assign Wpf6z6 = (~(Fth7z6[23] & Eye6z6));
assign Qof6z6 = (Mqf6z6 | Dqr8v6);
assign Aof6z6 = (Uqf6z6 & Crf6z6);
assign Crf6z6 = (~(Kxb7z6[15] & Mec6z6));
assign Uqf6z6 = (~(Ppb7z6[7] & Age6z6));
assign Gdf6z6 = (~(Svb6z6 & Itb7z6[15]));
assign HWDATAD[14] = (~(Krf6z6 & Srf6z6));
assign Srf6z6 = (~(Tim7z6[14] & Otb6z6));
assign Krf6z6 = (Asf6z6 & Isf6z6);
assign Isf6z6 = (~(Mub6z6 & Twq7x6));
assign Twq7x6 = (!Qsf6z6);
assign Qsf6z6 = (No7et6 ? I4e6z6 : Q4e6z6);
assign I4e6z6 = (Ysf6z6 & Gtf6z6);
assign Gtf6z6 = (Otf6z6 & Wtf6z6);
assign Wtf6z6 = (~(Awe6z6 & Eqc6z6));
assign Otf6z6 = (Euf6z6 & Muf6z6);
assign Muf6z6 = (~(Mue6z6 & Qoc6z6));
assign Euf6z6 = (~(I0f6z6 & Knc6z6));
assign Ysf6z6 = (Uuf6z6 & Cvf6z6);
assign Cvf6z6 = (~(Uic6z6 & Mqc6z6));
assign Uuf6z6 = (~(Kxb7z6[22] & Mec6z6));
assign Q4e6z6 = (Kvf6z6 & Svf6z6);
assign Svf6z6 = (Awf6z6 & Iwf6z6);
assign Iwf6z6 = (Qwf6z6 & Ywf6z6);
assign Ywf6z6 = (~(Mif6z6 & L2nov6));
assign L2nov6 = (~(Gxf6z6 & Oxf6z6));
assign Oxf6z6 = (~(Ohe7z6[6] & Kjf6z6));
assign Gxf6z6 = (~(Mfe7z6[6] & Ode6z6));
assign Qwf6z6 = (~(Agc6z6 & Qoc6z6));
assign Qoc6z6 = (~(Wxf6z6 & Eyf6z6));
assign Eyf6z6 = (~(Kxb7z6[30] & Wxe6z6));
assign Wxf6z6 = (Myf6z6 & Uyf6z6);
assign Uyf6z6 = (~(Fth7z6[30] & Eye6z6));
assign Myf6z6 = (~(Fhc7z6[30] & Ywe6z6));
assign Awf6z6 = (Czf6z6 & Kzf6z6);
assign Kzf6z6 = (~(Kre6z6 & Knc6z6));
assign Knc6z6 = (~(Szf6z6 & A0g6z6));
assign A0g6z6 = (~(Fhc7z6[6] & Ywe6z6));
assign Szf6z6 = (I0g6z6 & Q0g6z6);
assign Q0g6z6 = (~(Kxb7z6[6] & Wxe6z6));
assign I0g6z6 = (~(Fth7z6[6] & Eye6z6));
assign Czf6z6 = (~(Eue6z6 & Eqc6z6));
assign Eqc6z6 = (~(Y0g6z6 & G1g6z6));
assign G1g6z6 = (~(Kxb7z6[14] & Wxe6z6));
assign Y0g6z6 = (O1g6z6 & W1g6z6);
assign W1g6z6 = (~(Fth7z6[14] & Eye6z6));
assign O1g6z6 = (~(Fhc7z6[14] & Ywe6z6));
assign Kvf6z6 = (E2g6z6 & M2g6z6);
assign M2g6z6 = (U2g6z6 & C3g6z6);
assign C3g6z6 = (~(Mue6z6 & Mqc6z6));
assign Mqc6z6 = (~(K3g6z6 & S3g6z6));
assign S3g6z6 = (~(Fhc7z6[22] & Ywe6z6));
assign K3g6z6 = (A4g6z6 & I4g6z6);
assign I4g6z6 = (~(Kxb7z6[22] & Wxe6z6));
assign A4g6z6 = (~(Fth7z6[22] & Eye6z6));
assign U2g6z6 = (Mqf6z6 | Nnr8v6);
assign E2g6z6 = (Q4g6z6 & Y4g6z6);
assign Y4g6z6 = (~(Kxb7z6[14] & Mec6z6));
assign Q4g6z6 = (~(Ppb7z6[6] & Age6z6));
assign Asf6z6 = (~(Svb6z6 & Itb7z6[14]));
assign HWDATAD[13] = (~(G5g6z6 & O5g6z6));
assign O5g6z6 = (~(Tim7z6[13] & Otb6z6));
assign G5g6z6 = (W5g6z6 & E6g6z6);
assign E6g6z6 = (~(Mub6z6 & Vqq7x6));
assign Vqq7x6 = (!M6g6z6);
assign M6g6z6 = (No7et6 ? M6e6z6 : U6e6z6);
assign M6e6z6 = (U6g6z6 & C7g6z6);
assign C7g6z6 = (K7g6z6 & S7g6z6);
assign S7g6z6 = (~(Awe6z6 & G1d6z6));
assign K7g6z6 = (A8g6z6 & I8g6z6);
assign I8g6z6 = (~(Mue6z6 & Szc6z6));
assign A8g6z6 = (~(I0f6z6 & Uyc6z6));
assign U6g6z6 = (Q8g6z6 & Y8g6z6);
assign Y8g6z6 = (~(Uic6z6 & O1d6z6));
assign Q8g6z6 = (~(Kxb7z6[21] & Mec6z6));
assign U6e6z6 = (G9g6z6 & O9g6z6);
assign O9g6z6 = (W9g6z6 & Eag6z6);
assign Eag6z6 = (Mag6z6 & Uag6z6);
assign Uag6z6 = (~(Mif6z6 & Y5nov6));
assign Y5nov6 = (~(Cbg6z6 & Kbg6z6));
assign Kbg6z6 = (~(Ohe7z6[5] & Kjf6z6));
assign Kjf6z6 = (Sbg6z6 | Acg6z6);
assign Cbg6z6 = (~(Mfe7z6[5] & Ode6z6));
assign Mag6z6 = (~(Agc6z6 & Szc6z6));
assign Szc6z6 = (~(Icg6z6 & Qcg6z6));
assign Qcg6z6 = (~(Fhc7z6[29] & Ywe6z6));
assign Icg6z6 = (Ycg6z6 & Gdg6z6);
assign Gdg6z6 = (~(Kxb7z6[29] & Wxe6z6));
assign Ycg6z6 = (~(Fth7z6[29] & Eye6z6));
assign W9g6z6 = (Odg6z6 & Wdg6z6);
assign Wdg6z6 = (~(Kre6z6 & Uyc6z6));
assign Uyc6z6 = (~(Eeg6z6 & Meg6z6));
assign Meg6z6 = (~(Fhc7z6[5] & Ywe6z6));
assign Eeg6z6 = (Ueg6z6 & Cfg6z6);
assign Cfg6z6 = (~(Kxb7z6[5] & Wxe6z6));
assign Ueg6z6 = (~(Fth7z6[5] & Eye6z6));
assign Odg6z6 = (~(Eue6z6 & G1d6z6));
assign G1d6z6 = (~(Kfg6z6 & Sfg6z6));
assign Sfg6z6 = (~(Fhc7z6[13] & Ywe6z6));
assign Kfg6z6 = (Agg6z6 & Igg6z6);
assign Igg6z6 = (~(Kxb7z6[13] & Wxe6z6));
assign Agg6z6 = (~(Fth7z6[13] & Eye6z6));
assign G9g6z6 = (Qgg6z6 & Ygg6z6);
assign Ygg6z6 = (Ghg6z6 & Ohg6z6);
assign Ohg6z6 = (~(Mue6z6 & O1d6z6));
assign O1d6z6 = (~(Whg6z6 & Eig6z6));
assign Eig6z6 = (~(Fhc7z6[21] & Ywe6z6));
assign Whg6z6 = (Mig6z6 & Uig6z6);
assign Uig6z6 = (~(Kxb7z6[21] & Wxe6z6));
assign Mig6z6 = (~(Fth7z6[21] & Eye6z6));
assign Ghg6z6 = (Mqf6z6 | Xkr8v6);
assign Qgg6z6 = (Cjg6z6 & Kjg6z6);
assign Kjg6z6 = (~(Kxb7z6[13] & Mec6z6));
assign Cjg6z6 = (~(Ppb7z6[5] & Age6z6));
assign W5g6z6 = (~(Svb6z6 & Itb7z6[13]));
assign HWDATAD[12] = (~(Sjg6z6 & Akg6z6));
assign Akg6z6 = (~(Tim7z6[12] & Otb6z6));
assign Sjg6z6 = (Ikg6z6 & Qkg6z6);
assign Qkg6z6 = (~(Mub6z6 & Llq7x6));
assign Llq7x6 = (!Ykg6z6);
assign Ykg6z6 = (No7et6 ? Q8e6z6 : Y8e6z6);
assign Q8e6z6 = (Glg6z6 & Olg6z6);
assign Olg6z6 = (Wlg6z6 & Emg6z6);
assign Emg6z6 = (~(Awe6z6 & Ead6z6));
assign Wlg6z6 = (Mmg6z6 & Umg6z6);
assign Umg6z6 = (~(Mue6z6 & Q8d6z6));
assign Mmg6z6 = (~(I0f6z6 & S7d6z6));
assign Glg6z6 = (Cng6z6 & Kng6z6);
assign Kng6z6 = (~(Uic6z6 & Mad6z6));
assign Cng6z6 = (~(Kxb7z6[20] & Mec6z6));
assign Y8e6z6 = (Sng6z6 & Aog6z6);
assign Aog6z6 = (Iog6z6 & Qog6z6);
assign Qog6z6 = (Yog6z6 & Gpg6z6);
assign Gpg6z6 = (~(Mif6z6 & Gwmov6));
assign Gwmov6 = (~(Opg6z6 & Wpg6z6));
assign Wpg6z6 = (~(Acg6z6 & Ohe7z6[4]));
assign Opg6z6 = (Eqg6z6 & Mqg6z6);
assign Mqg6z6 = (~(Mfe7z6[4] & Ode6z6));
assign Eqg6z6 = (~(N0gdt6 & Sbg6z6));
assign Mif6z6 = (Ycc6z6 & Uqg6z6);
assign Uqg6z6 = (Rysiw6 | Srviy6);
assign Rysiw6 = (!Otsiw6);
assign Yog6z6 = (Mqf6z6 | Hir8v6);
assign Mqf6z6 = (~(Crg6z6 & Otsiw6));
assign Otsiw6 = (Krg6z6 & Srg6z6);
assign Srg6z6 = (~(Asg6z6 | Isg6z6));
assign Asg6z6 = (Qsg6z6 | Ohe7z6[2]);
assign Krg6z6 = (Ysg6z6 & Gtg6z6);
assign Ysg6z6 = (Mud6z6 & Yce6z6);
assign Yce6z6 = (~(Ohe7z6[1] & Sbg6z6));
assign Mud6z6 = (Otg6z6 & Wtg6z6);
assign Wtg6z6 = (~(Acg6z6 & Ohe7z6[1]));
assign Otg6z6 = (Eug6z6 & Mug6z6);
assign Mug6z6 = (~(Ohe7z6[3] & Ode6z6));
assign Eug6z6 = (~(Sbg6z6 & Ohe7z6[2]));
assign Crg6z6 = (~(Srviy6 | Uud6z6));
assign Srviy6 = (Ldo7v6 & Tnzdt6);
assign Iog6z6 = (Uug6z6 & Cvg6z6);
assign Cvg6z6 = (~(Agc6z6 & Q8d6z6));
assign Q8d6z6 = (~(Kvg6z6 & Svg6z6));
assign Svg6z6 = (~(Kxb7z6[28] & Wxe6z6));
assign Kvg6z6 = (Awg6z6 & Iwg6z6);
assign Iwg6z6 = (~(Fth7z6[28] & Eye6z6));
assign Awg6z6 = (~(Fhc7z6[28] & Ywe6z6));
assign Uug6z6 = (~(Kre6z6 & S7d6z6));
assign S7d6z6 = (~(Qwg6z6 & Ywg6z6));
assign Ywg6z6 = (~(Kxb7z6[4] & Wxe6z6));
assign Qwg6z6 = (Gxg6z6 & Oxg6z6);
assign Oxg6z6 = (~(E3c7z6[4] & Ywe6z6));
assign Gxg6z6 = (~(Fth7z6[4] & Eye6z6));
assign Sng6z6 = (Wxg6z6 & Eyg6z6);
assign Eyg6z6 = (~(Kxb7z6[12] & Mec6z6));
assign Wxg6z6 = (Myg6z6 & Uyg6z6);
assign Uyg6z6 = (~(Eue6z6 & Ead6z6));
assign Ead6z6 = (~(Czg6z6 & Kzg6z6));
assign Kzg6z6 = (~(Fhc7z6[12] & Ywe6z6));
assign Czg6z6 = (Szg6z6 & A0h6z6);
assign A0h6z6 = (~(Kxb7z6[12] & Wxe6z6));
assign Szg6z6 = (~(Fth7z6[12] & Eye6z6));
assign Myg6z6 = (~(Mue6z6 & Mad6z6));
assign Mad6z6 = (~(I0h6z6 & Q0h6z6));
assign Q0h6z6 = (~(Fhc7z6[20] & Ywe6z6));
assign I0h6z6 = (Y0h6z6 & G1h6z6);
assign G1h6z6 = (~(Kxb7z6[20] & Wxe6z6));
assign Y0h6z6 = (~(Fth7z6[20] & Eye6z6));
assign Ikg6z6 = (~(Svb6z6 & Itb7z6[12]));
assign HWDATAD[11] = (~(O1h6z6 & W1h6z6));
assign W1h6z6 = (~(Tim7z6[11] & Otb6z6));
assign O1h6z6 = (E2h6z6 & M2h6z6);
assign M2h6z6 = (~(Mub6z6 & Bgq7x6));
assign Bgq7x6 = (!U2h6z6);
assign U2h6z6 = (No7et6 ? Wle6z6 : Eme6z6);
assign Wle6z6 = (C3h6z6 & K3h6z6);
assign K3h6z6 = (S3h6z6 & A4h6z6);
assign A4h6z6 = (~(Awe6z6 & Cjd6z6));
assign S3h6z6 = (I4h6z6 & Q4h6z6);
assign Q4h6z6 = (~(Mue6z6 & Ohd6z6));
assign I4h6z6 = (~(I0f6z6 & Qgd6z6));
assign C3h6z6 = (Y4h6z6 & G5h6z6);
assign G5h6z6 = (~(Uic6z6 & Kjd6z6));
assign Y4h6z6 = (~(Kxb7z6[19] & Mec6z6));
assign Eme6z6 = (O5h6z6 & W5h6z6);
assign W5h6z6 = (E6h6z6 & M6h6z6);
assign M6h6z6 = (~(Kre6z6 & Qgd6z6));
assign Qgd6z6 = (~(U6h6z6 & C7h6z6));
assign C7h6z6 = (~(Kxb7z6[3] & Wxe6z6));
assign U6h6z6 = (K7h6z6 & S7h6z6);
assign S7h6z6 = (~(E3c7z6[3] & Ywe6z6));
assign K7h6z6 = (~(Fth7z6[3] & Eye6z6));
assign E6h6z6 = (A8h6z6 & I8h6z6);
assign I8h6z6 = (Gtg6z6 | Uud6z6);
assign Uud6z6 = (!Ycc6z6);
assign Gtg6z6 = (Q8h6z6 & Y8h6z6);
assign Y8h6z6 = (~(Ohe7z6[3] & Acg6z6));
assign Q8h6z6 = (G9h6z6 & O9h6z6);
assign O9h6z6 = (~(Mfe7z6[3] & Ode6z6));
assign G9h6z6 = (~(Ohe7z6[4] & Sbg6z6));
assign A8h6z6 = (~(Agc6z6 & Ohd6z6));
assign Ohd6z6 = (~(W9h6z6 & Eah6z6));
assign Eah6z6 = (~(Fhc7z6[27] & Ywe6z6));
assign W9h6z6 = (Mah6z6 & Uah6z6);
assign Uah6z6 = (~(Kxb7z6[27] & Wxe6z6));
assign Mah6z6 = (~(Fth7z6[27] & Eye6z6));
assign O5h6z6 = (Cbh6z6 & Kbh6z6);
assign Kbh6z6 = (~(Kxb7z6[11] & Mec6z6));
assign Cbh6z6 = (Sbh6z6 & Ach6z6);
assign Ach6z6 = (~(Eue6z6 & Cjd6z6));
assign Cjd6z6 = (~(Ich6z6 & Qch6z6));
assign Qch6z6 = (~(Fhc7z6[11] & Ywe6z6));
assign Ich6z6 = (Ych6z6 & Gdh6z6);
assign Gdh6z6 = (~(Kxb7z6[11] & Wxe6z6));
assign Ych6z6 = (~(Fth7z6[11] & Eye6z6));
assign Sbh6z6 = (~(Mue6z6 & Kjd6z6));
assign Kjd6z6 = (~(Odh6z6 & Wdh6z6));
assign Wdh6z6 = (~(Fhc7z6[19] & Ywe6z6));
assign Odh6z6 = (Eeh6z6 & Meh6z6);
assign Meh6z6 = (~(Kxb7z6[19] & Wxe6z6));
assign Eeh6z6 = (~(Fth7z6[19] & Eye6z6));
assign E2h6z6 = (~(Svb6z6 & Itb7z6[11]));
assign HWDATAD[10] = (~(Ueh6z6 & Cfh6z6));
assign Cfh6z6 = (~(Tim7z6[10] & Otb6z6));
assign Ueh6z6 = (Kfh6z6 & Sfh6z6);
assign Sfh6z6 = (~(Mub6z6 & Raq7x6));
assign Raq7x6 = (!Agh6z6);
assign Agh6z6 = (No7et6 ? Aoe6z6 : Ioe6z6);
assign Aoe6z6 = (Igh6z6 & Qgh6z6);
assign Qgh6z6 = (Ygh6z6 & Ghh6z6);
assign Ghh6z6 = (~(Awe6z6 & Asd6z6));
assign Awe6z6 = (Ohh6z6 & Whh6z6);
assign Whh6z6 = (~(Eih6z6 & Mih6z6));
assign Ygh6z6 = (Uih6z6 & Cjh6z6);
assign Cjh6z6 = (~(Mue6z6 & Mqd6z6));
assign Uih6z6 = (~(I0f6z6 & Opd6z6));
assign I0f6z6 = (Ohh6z6 & Kjh6z6);
assign Kjh6z6 = (~(Sjh6z6 & Akh6z6));
assign Sjh6z6 = (Ikh6z6 & Qkh6z6);
assign Igh6z6 = (Ykh6z6 & Glh6z6);
assign Glh6z6 = (~(Uic6z6 & Isd6z6));
assign Ykh6z6 = (~(Kxb7z6[18] & Mec6z6));
assign Ioe6z6 = (Olh6z6 & Wlh6z6);
assign Wlh6z6 = (Emh6z6 & Mmh6z6);
assign Mmh6z6 = (~(Eue6z6 & Asd6z6));
assign Asd6z6 = (~(Umh6z6 & Cnh6z6));
assign Cnh6z6 = (~(Fhc7z6[10] & Ywe6z6));
assign Umh6z6 = (Knh6z6 & Snh6z6);
assign Snh6z6 = (~(Kxb7z6[10] & Wxe6z6));
assign Knh6z6 = (~(Fth7z6[10] & Eye6z6));
assign Eue6z6 = (Aoh6z6 & Ioh6z6);
assign Emh6z6 = (Qoh6z6 & Yoh6z6);
assign Yoh6z6 = (~(Gph6z6 & Ycc6z6));
assign Gph6z6 = (~(Oph6z6 & Wph6z6));
assign Wph6z6 = (~(Acg6z6 & Ohe7z6[2]));
assign Oph6z6 = (~(Isg6z6 | Qsg6z6));
assign Qsg6z6 = (Ohe7z6[4] & Ode6z6);
assign Isg6z6 = (Ohe7z6[3] & Sbg6z6);
assign Sbg6z6 = (~(Acg6z6 | Ode6z6));
assign Ode6z6 = (Eqh6z6 & Oyfdt6);
assign Eqh6z6 = (Tnzdt6 & Kgbdt6);
assign Acg6z6 = (~(Gpsiw6 | Ldo7v6));
assign Qoh6z6 = (~(Kre6z6 & Opd6z6));
assign Opd6z6 = (~(Mqh6z6 & Uqh6z6));
assign Uqh6z6 = (~(Kxb7z6[2] & Wxe6z6));
assign Mqh6z6 = (Crh6z6 & Krh6z6);
assign Krh6z6 = (~(E3c7z6[2] & Ywe6z6));
assign Crh6z6 = (~(Fth7z6[2] & Eye6z6));
assign Kre6z6 = (Ohh6z6 & Srh6z6);
assign Srh6z6 = (~(Ash6z6 & Eih6z6));
assign Olh6z6 = (Ish6z6 & Qsh6z6);
assign Qsh6z6 = (~(Kxb7z6[10] & Mec6z6));
assign Ish6z6 = (Ysh6z6 & Gth6z6);
assign Gth6z6 = (~(Agc6z6 & Mqd6z6));
assign Mqd6z6 = (~(Oth6z6 & Wth6z6));
assign Wth6z6 = (~(Fhc7z6[26] & Ywe6z6));
assign Oth6z6 = (Euh6z6 & Muh6z6);
assign Muh6z6 = (~(Kxb7z6[26] & Wxe6z6));
assign Euh6z6 = (~(Fth7z6[26] & Eye6z6));
assign Ysh6z6 = (~(Mue6z6 & Isd6z6));
assign Isd6z6 = (~(Uuh6z6 & Cvh6z6));
assign Cvh6z6 = (~(Fhc7z6[18] & Ywe6z6));
assign Uuh6z6 = (Kvh6z6 & Svh6z6);
assign Svh6z6 = (~(Kxb7z6[18] & Wxe6z6));
assign Kvh6z6 = (~(Fth7z6[18] & Eye6z6));
assign Mue6z6 = (~(Awh6z6 | Iwh6z6));
assign Kfh6z6 = (~(Svb6z6 & Itb7z6[10]));
assign HWDATAD[0] = (~(Qwh6z6 & Ywh6z6));
assign Ywh6z6 = (~(Mub6z6 & I8r7x6));
assign I8r7x6 = (!Gxh6z6);
assign Gxh6z6 = (No7et6 ? A0e6z6 : I0e6z6);
assign A0e6z6 = (Oxh6z6 & Wxh6z6);
assign Wxh6z6 = (Eyh6z6 & Myh6z6);
assign Myh6z6 = (Uyh6z6 & Czh6z6);
assign Czh6z6 = (~(Cjc6z6 & K7f6z6));
assign Cjc6z6 = (Ohh6z6 & Kzh6z6);
assign Kzh6z6 = (~(Ash6z6 & Iwh6z6));
assign Ash6z6 = (Mih6z6 & Qkh6z6);
assign Qkh6z6 = (!Eylxx6);
assign Uyh6z6 = (~(Whc6z6 & M6f6z6));
assign Whc6z6 = (Ohh6z6 & Szh6z6);
assign Szh6z6 = (~(Akh6z6 & Ikh6z6));
assign Eyh6z6 = (A0i6z6 & I0i6z6);
assign I0i6z6 = (~(Gdc6z6 & Y8f6z6));
assign A0i6z6 = (~(Uic6z6 & G9f6z6));
assign Uic6z6 = (Ioh6z6 & Q0i6z6);
assign Q0i6z6 = (~(Y0i6z6 & X7vxx6));
assign Oxh6z6 = (G1i6z6 & O1i6z6);
assign O1i6z6 = (~(Lybdt6 & Ycc6z6));
assign G1i6z6 = (W1i6z6 & E2i6z6);
assign E2i6z6 = (~(Kxb7z6[24] & Mec6z6));
assign W1i6z6 = (~(Tkbdt6 & Age6z6));
assign I0e6z6 = (M2i6z6 & U2i6z6);
assign U2i6z6 = (C3i6z6 & K3i6z6);
assign K3i6z6 = (S3i6z6 & A4i6z6);
assign A4i6z6 = (~(Kfc6z6 & M6f6z6));
assign M6f6z6 = (~(I4i6z6 & Q4i6z6));
assign Q4i6z6 = (~(Fhc7z6[8] & Ywe6z6));
assign I4i6z6 = (Y4i6z6 & G5i6z6);
assign G5i6z6 = (~(Kxb7z6[8] & Wxe6z6));
assign Y4i6z6 = (~(Fth7z6[8] & Eye6z6));
assign Kfc6z6 = (Ohh6z6 & O5i6z6);
assign O5i6z6 = (~(Iwh6z6 & Mih6z6));
assign Mih6z6 = (~(Bqoxx6 & Kih7z6[0]));
assign Iwh6z6 = (Bavxx6 & D9vxx6);
assign D9vxx6 = (~(Dca7x6 & W5i6z6));
assign Bavxx6 = (~(E6i6z6 & Gaa7x6));
assign S3i6z6 = (~(Qm0jw6 & Ycc6z6));
assign Ycc6z6 = (~(M6i6z6 & U6i6z6));
assign U6i6z6 = (~(C7i6z6 & K7i6z6));
assign K7i6z6 = (Fcmyx6 & S7i6z6);
assign Fcmyx6 = (!Qij7z6[2]);
assign C7i6z6 = (Ldmyx6 & Tdmyx6);
assign M6i6z6 = (~(Rioov6 & Gdviy6));
assign Gdviy6 = (!Igniy6);
assign Qm0jw6 = (Nob7z6[0] & Rslov6);
assign Rslov6 = (!J2cdt6);
assign C3i6z6 = (A8i6z6 & I8i6z6);
assign I8i6z6 = (~(Agc6z6 & Y8f6z6));
assign Y8f6z6 = (~(Q8i6z6 & Y8i6z6));
assign Y8i6z6 = (~(Fhc7z6[16] & Ywe6z6));
assign Q8i6z6 = (G9i6z6 & O9i6z6);
assign O9i6z6 = (~(Kxb7z6[16] & Wxe6z6));
assign G9i6z6 = (~(Fth7z6[16] & Eye6z6));
assign Agc6z6 = (~(Akh6z6 | Awh6z6));
assign Akh6z6 = (!L9vxx6);
assign L9vxx6 = (H287x6 & Edh7z6[1]);
assign H287x6 = (~(W9i6z6 | Kih7z6[0]));
assign A8i6z6 = (~(Sbc6z6 & K7f6z6));
assign K7f6z6 = (~(Eai6z6 & Mai6z6));
assign Mai6z6 = (~(Kxb7z6[0] & Wxe6z6));
assign Eai6z6 = (Uai6z6 & Cbi6z6);
assign Cbi6z6 = (~(E3c7z6[0] & Ywe6z6));
assign Uai6z6 = (~(Fth7z6[0] & Eye6z6));
assign Sbc6z6 = (Ioh6z6 & Kbi6z6);
assign Kbi6z6 = (Aoh6z6 | Eylxx6);
assign Eylxx6 = (~(Edh7z6[0] | Edh7z6[1]));
assign Aoh6z6 = (~(Sbi6z6 & Ikh6z6));
assign Ikh6z6 = (~(Bqoxx6 & Aci6z6));
assign Bqoxx6 = (Edh7z6[0] & Ici6z6);
assign Sbi6z6 = (Y0i6z6 & X7vxx6);
assign X7vxx6 = (~(Av77x6 & Edh7z6[1]));
assign Av77x6 = (~(Kih7z6[1] | Kih7z6[0]));
assign Ioh6z6 = (~(Awh6z6 & Y0i6z6));
assign Y0i6z6 = (~(Ow2et6 & X7yxx6));
assign M2i6z6 = (Qci6z6 & Yci6z6);
assign Yci6z6 = (~(Nmadt6 & Age6z6));
assign Age6z6 = (Gdi6z6 & Odi6z6);
assign Odi6z6 = (Tdmyx6 & S7i6z6);
assign Gdi6z6 = (Qij7z6[2] & Ldmyx6);
assign Qci6z6 = (Wdi6z6 & Eei6z6);
assign Eei6z6 = (~(Gdc6z6 & G9f6z6));
assign G9f6z6 = (~(Mei6z6 & Uei6z6));
assign Uei6z6 = (~(Fhc7z6[24] & Ywe6z6));
assign Ywe6z6 = (~(Cfi6z6 | Eye6z6));
assign Cfi6z6 = (!Xnh7z6[0]);
assign Mei6z6 = (Kfi6z6 & Sfi6z6);
assign Sfi6z6 = (~(Kxb7z6[24] & Wxe6z6));
assign Wxe6z6 = (~(Eye6z6 | Xnh7z6[0]));
assign Kfi6z6 = (~(Fth7z6[24] & Eye6z6));
assign Eye6z6 = (~(Agi6z6 & Igi6z6));
assign Igi6z6 = (~(Clhhw6 & Eikiy6));
assign Eikiy6 = (Qgi6z6 & Ygi6z6);
assign Ygi6z6 = (Ghi6z6 & Ohi6z6);
assign Ghi6z6 = (Whi6z6 & Eii6z6);
assign Eii6z6 = (~(P4c7z6[0] & Hir8v6));
assign Qgi6z6 = (Mii6z6 & Glkiy6);
assign Glkiy6 = (~(Mii6z6 & Uii6z6));
assign Uii6z6 = (~(Cji6z6 & Kji6z6));
assign Kji6z6 = (~(Sji6z6 & Aki6z6));
assign Aki6z6 = (~(Iki6z6 & Qki6z6));
assign Qki6z6 = (~(Pxmov6 & C7piy6));
assign C7piy6 = (!P4c7z6[0]);
assign Iki6z6 = (~(Xumov6 & O9kiy6));
assign Sji6z6 = (Ohi6z6 & Whi6z6);
assign Whi6z6 = (Oppiy6 | Kpaov6);
assign Ohi6z6 = (O9kiy6 | Xumov6);
assign Xumov6 = (!Xkr8v6);
assign O9kiy6 = (!P4c7z6[1]);
assign Cji6z6 = (~(Yki6z6 & Gli6z6));
assign Gli6z6 = (~(P4c7z6[3] & Nnr8v6));
assign Yki6z6 = (Oli6z6 & Y8niy6);
assign Y8niy6 = (!Ycniy6);
assign Oli6z6 = (~(P4c7z6[2] & Wli6z6));
assign Wli6z6 = (~(Xlaov6 & Whpiy6));
assign Whpiy6 = (!P4c7z6[3]);
assign Mii6z6 = (~(P4c7z6[3] & Dqr8v6));
assign Agi6z6 = (~(Dzkiw6 | Emi6z6));
assign Emi6z6 = (Mmi6z6 & Ecc7z6[10]);
assign Mmi6z6 = (Vxihw6 & Umi6z6);
assign Umi6z6 = (~(Cni6z6 & Kni6z6));
assign Kni6z6 = (~(Sni6z6 & Aoi6z6));
assign Aoi6z6 = (Ioi6z6 & Qoi6z6);
assign Qoi6z6 = (P4c7z6[0] ^ A8piy6);
assign A8piy6 = (!Pxg7z6[0]);
assign Ioi6z6 = (Yoi6z6 & Ot97x6);
assign Yoi6z6 = (P4c7z6[1] ^ C8a7x6);
assign C8a7x6 = (!Pxg7z6[1]);
assign Sni6z6 = (Gpi6z6 & Opi6z6);
assign Opi6z6 = (~(Oppiy6 ^ Aopiy6));
assign Aopiy6 = (!Pxg7z6[2]);
assign Oppiy6 = (!P4c7z6[2]);
assign Gpi6z6 = (P4c7z6[3] ^ Akpiy6);
assign Akpiy6 = (!Pxg7z6[3]);
assign Cni6z6 = (~(Wpi6z6 & Eqi6z6));
assign Eqi6z6 = (Mqi6z6 & Uqi6z6);
assign Uqi6z6 = (P4c7z6[0] ^ Gclhw6);
assign Gclhw6 = (!Ntg7z6[0]);
assign Mqi6z6 = (Cri6z6 & Yckiy6);
assign Yckiy6 = (Px97x6 & Doihw6);
assign Px97x6 = (~(Zna7x6 | Mpihw6));
assign Cri6z6 = (P4c7z6[1] ^ Pdlhw6);
assign Pdlhw6 = (!Ntg7z6[1]);
assign Wpi6z6 = (Kri6z6 & Sri6z6);
assign Sri6z6 = (P4c7z6[2] ^ Yelhw6);
assign Yelhw6 = (!Ntg7z6[2]);
assign Kri6z6 = (P4c7z6[3] ^ Oglhw6);
assign Oglhw6 = (!Ntg7z6[3]);
assign Vxihw6 = (Ecc7z6[9] & Pbadt6);
assign Dzkiw6 = (Thbet6 & Xnh7z6[1]);
assign Gdc6z6 = (~(Awh6z6 | Eih6z6));
assign Eih6z6 = (P7vxx6 & Zavxx6);
assign Zavxx6 = (~(W5i6z6 & Gaa7x6));
assign Gaa7x6 = (~(W9i6z6 | Aci6z6));
assign W9i6z6 = (!Kih7z6[1]);
assign W5i6z6 = (~(Xgmov6 | Ici6z6));
assign Xgmov6 = (!No7et6);
assign P7vxx6 = (~(E6i6z6 & Dca7x6));
assign Dca7x6 = (~(Aci6z6 | Kih7z6[1]));
assign Aci6z6 = (!Kih7z6[0]);
assign E6i6z6 = (~(Ici6z6 | No7et6));
assign Ici6z6 = (!Edh7z6[1]);
assign Awh6z6 = (!Ohh6z6);
assign Ohh6z6 = (~(Asi6z6 | Spdiw6));
assign Spdiw6 = (!Thbet6);
assign Asi6z6 = (Ztaov6 ? S7i6z6 : Isi6z6);
assign Isi6z6 = (~(Qsi6z6 & Ysi6z6));
assign Ysi6z6 = (Gti6z6 & Oti6z6);
assign Oti6z6 = (X3yxx6 & Qsaov6);
assign Gti6z6 = (T1yxx6 & Ruvxx6);
assign Ruvxx6 = (!Rhihw6);
assign Rhihw6 = (Wti6z6 & Dioov6);
assign Wti6z6 = (Lpwxx6 & Bwvnv6);
assign Qsi6z6 = (Eui6z6 & Mui6z6);
assign Eui6z6 = (~(Uui6z6 | X7yxx6));
assign X7yxx6 = (~(Vkhhw6 & Ajihw6));
assign Ajihw6 = (~(Cvi6z6 & Fulnv6));
assign Cvi6z6 = (Doihw6 & Dwb7z6[3]);
assign Vkhhw6 = (!Ot97x6);
assign Wdi6z6 = (~(Kxb7z6[0] & Mec6z6));
assign Mec6z6 = (~(Kvi6z6 & Svi6z6));
assign Svi6z6 = (Awi6z6 & Iwi6z6);
assign Iwi6z6 = (~(Qwi6z6 & Ldmyx6));
assign Ldmyx6 = (Ywi6z6 & Ztaov6);
assign Ztaov6 = (Kioov6 & G5kiy6);
assign Ywi6z6 = (~(Qij7z6[5] | Qij7z6[6]));
assign Qwi6z6 = (Gxi6z6 & S7i6z6);
assign S7i6z6 = (!X4eet6);
assign Gxi6z6 = (!Tdmyx6);
assign Tdmyx6 = (~(Tdwxx6 | R2vxx6));
assign R2vxx6 = (Qij7z6[1] | Qij7z6[0]);
assign Tdwxx6 = (!Qij7z6[4]);
assign Awi6z6 = (~(Xdphw6 & Oxi6z6));
assign Oxi6z6 = (Uui6z6 | Wxi6z6);
assign Uui6z6 = (~(J1a7x6 & Eyi6z6));
assign Xdphw6 = (!Yioov6);
assign Yioov6 = (Igniy6 | 1'b0);
assign Kvi6z6 = (Mui6z6 & Myi6z6);
assign Myi6z6 = (~(Rioov6 & Igniy6));
assign Mui6z6 = (Uyi6z6 & Czi6z6);
assign Czi6z6 = (~(Ggoov6 & Vqihw6));
assign Uyi6z6 = (Gwsiw6 & Elphw6);
assign Elphw6 = (!Ef47x6);
assign Ef47x6 = (Ggoov6 & Fxaov6);
assign Mub6z6 = (Eqn7z6[0] & Kzi6z6);
assign Qwh6z6 = (Szi6z6 & A0j6z6);
assign A0j6z6 = (~(Svb6z6 & Itb7z6[0]));
assign Svb6z6 = (Eqn7z6[1] & Kzi6z6);
assign Szi6z6 = (~(Tim7z6[0] & Otb6z6));
assign Otb6z6 = (Eqn7z6[2] | I0j6z6);
assign I0j6z6 = (!Kzi6z6);
assign Kzi6z6 = (~(Sb0jy6 & Qln7z6[0]));
assign Sb0jy6 = (Q0j6z6 & Qakiw6);
assign HTRANSS[1] = (Y0j6z6 & G1j6z6);
assign G1j6z6 = (~(O1j6z6 & W1j6z6));
assign W1j6z6 = (Uaonv6 | E2j6z6);
assign HTRANSS[0] = (M2j6z6 & U2j6z6);
assign M2j6z6 = (Aoa6z6 & Y0j6z6);
assign Y0j6z6 = (C3j6z6 & K3j6z6);
assign K3j6z6 = (~(Rj9ov6 & Nhonv6));
assign C3j6z6 = (~(Qmonv6 & J0jxx6));
assign HTRANSI[1] = (Yk1ov6 | S3j6z6);
assign S3j6z6 = (U4zet6 & Am1ov6);
assign Yk1ov6 = (A4j6z6 & I4j6z6);
assign I4j6z6 = (Uy76z6 & Cfliy6);
assign Cfliy6 = (~(Q4j6z6 | Woyet6));
assign Q4j6z6 = (~(Cakiw6 | Benyx6));
assign Uy76z6 = (Y4j6z6 & U6y5z6);
assign Y4j6z6 = (~(DNOTITRANS & HTRANSD[1]));
assign A4j6z6 = (Lbkiw6 & Njkiw6);
assign Njkiw6 = (~(Xnmyx6 | Njfnv6));
assign Njfnv6 = (Crcdt6 ? Dvc7z6[31] : X0d7z6[31]);
assign X0d7z6[31] = (~(G5j6z6 & O5j6z6));
assign O5j6z6 = (W5j6z6 & E6j6z6);
assign E6j6z6 = (~(Pic7z6[31] & Ir0ov6));
assign W5j6z6 = (M6j6z6 & U6j6z6);
assign U6j6z6 = (Qs46z6 | Z0xnv6);
assign Z0xnv6 = (C7j6z6 & K7j6z6);
assign K7j6z6 = (~(Wkd7z6[31] & Ddmhw6));
assign C7j6z6 = (S7j6z6 & A8j6z6);
assign A8j6z6 = (~(Xhd7z6[31] & Eu46z6));
assign S7j6z6 = (~(Vnd7z6[31] & Jamnv6));
assign M6j6z6 = (~(Pdc7z6[31] & Mu46z6));
assign G5j6z6 = (I8j6z6 & Q8j6z6);
assign Q8j6z6 = (~(Pnb7z6[31] & Znnov6));
assign I8j6z6 = (~(Qdcdt6 & Fhc7z6[31]));
assign Xnmyx6 = (~(Bw3nv6 & Zn3nv6));
assign Zn3nv6 = (!Ujfnv6);
assign Ujfnv6 = (Crcdt6 ? Dvc7z6[30] : X0d7z6[30]);
assign X0d7z6[30] = (~(Y8j6z6 & G9j6z6));
assign G9j6z6 = (O9j6z6 & W9j6z6);
assign W9j6z6 = (~(Pic7z6[30] & Ir0ov6));
assign O9j6z6 = (Eaj6z6 & Maj6z6);
assign Maj6z6 = (Qs46z6 | Xdxnv6);
assign Xdxnv6 = (Uaj6z6 & Cbj6z6);
assign Cbj6z6 = (~(Wkd7z6[30] & Ddmhw6));
assign Uaj6z6 = (Kbj6z6 & Sbj6z6);
assign Sbj6z6 = (~(Xhd7z6[30] & Eu46z6));
assign Kbj6z6 = (~(Vnd7z6[30] & Jamnv6));
assign Eaj6z6 = (~(Pdc7z6[30] & Mu46z6));
assign Y8j6z6 = (Acj6z6 & Icj6z6);
assign Icj6z6 = (~(Pnb7z6[30] & Znnov6));
assign Acj6z6 = (~(Qdcdt6 & Fhc7z6[30]));
assign Bw3nv6 = (!Bkfnv6);
assign Bkfnv6 = (Crcdt6 ? Dvc7z6[29] : X0d7z6[29]);
assign X0d7z6[29] = (~(Qcj6z6 & Ycj6z6));
assign Ycj6z6 = (Gdj6z6 & Odj6z6);
assign Odj6z6 = (~(Pic7z6[29] & Ir0ov6));
assign Gdj6z6 = (Wdj6z6 & Eej6z6);
assign Eej6z6 = (Qs46z6 | Mixnv6);
assign Mixnv6 = (Mej6z6 & Uej6z6);
assign Uej6z6 = (~(Wkd7z6[29] & Ddmhw6));
assign Mej6z6 = (Cfj6z6 & Kfj6z6);
assign Kfj6z6 = (~(Xhd7z6[29] & Eu46z6));
assign Cfj6z6 = (~(Vnd7z6[29] & Jamnv6));
assign Wdj6z6 = (~(Pdc7z6[29] & Mu46z6));
assign Qcj6z6 = (Sfj6z6 & Agj6z6);
assign Agj6z6 = (~(Pnb7z6[29] & Znnov6));
assign Sfj6z6 = (~(Qdcdt6 & Fhc7z6[29]));
assign Lbkiw6 = (Am1ov6 & Ygo7v6);
assign Am1ov6 = (Crcdt6 ? Aocdt6 : Lh1ov6);
assign Lh1ov6 = (~(Igj6z6 & Qgj6z6));
assign Qgj6z6 = (Ygj6z6 & Ghj6z6);
assign Ghj6z6 = (~(Ohj6z6 & Cgc7z6[2]));
assign Ohj6z6 = (Whj6z6 & Eij6z6);
assign Eij6z6 = (~(Mij6z6 & P1piw6));
assign Mij6z6 = (~(Uij6z6 & Ckihw6));
assign Ckihw6 = (Q0wnv6 & Qg2nv6);
assign Q0wnv6 = (!K9d7x6);
assign K9d7x6 = (D9d7x6 | Cubdt6);
assign D9d7x6 = (Cjj6z6 & Kjj6z6);
assign Kjj6z6 = (Sjj6z6 & Akj6z6);
assign Akj6z6 = (Ikj6z6 & Qkj6z6);
assign Qkj6z6 = (Ykj6z6 & Glj6z6);
assign Glj6z6 = (Olj6z6 & Fhc7z6[9]);
assign Olj6z6 = (Fhc7z6[25] & Pxfov6);
assign Pxfov6 = (Uobdt6 ? Wlj6z6 : C7riy6);
assign Wlj6z6 = (Tk8iw6 ^ Ide7z6[0]);
assign C7riy6 = (Knbdt6 ? W9edt6 : Acedt6);
assign Ykj6z6 = (Fhc7z6[27] & Fhc7z6[17]);
assign Ikj6z6 = (Emj6z6 & Mmj6z6);
assign Mmj6z6 = (Fhc7z6[19] & Fhc7z6[11]);
assign Emj6z6 = (E3c7z6[4] & Fhc7z6[28]);
assign Sjj6z6 = (Umj6z6 & Cnj6z6);
assign Cnj6z6 = (Knj6z6 & Snj6z6);
assign Snj6z6 = (Aoj6z6 & Fhc7z6[31]);
assign Aoj6z6 = (Fhc7z6[20] & Fhc7z6[12]);
assign Knj6z6 = (Fhc7z6[15] & Fhc7z6[7]);
assign Umj6z6 = (Ioj6z6 & Qoj6z6);
assign Qoj6z6 = (Fhc7z6[8] & Fhc7z6[23]);
assign Ioj6z6 = (Fhc7z6[24] & Fhc7z6[16]);
assign Cjj6z6 = (Yoj6z6 & Gpj6z6);
assign Gpj6z6 = (Opj6z6 & Wpj6z6);
assign Wpj6z6 = (Eqj6z6 & Mqj6z6);
assign Mqj6z6 = (Uqj6z6 & Fhc7z6[18]);
assign Uqj6z6 = (Fhc7z6[10] & Fhc7z6[26]);
assign Eqj6z6 = (Fhc7z6[6] & Fhc7z6[30]);
assign Opj6z6 = (Crj6z6 & Krj6z6);
assign Krj6z6 = (Fhc7z6[22] & Fhc7z6[14]);
assign Crj6z6 = (Fhc7z6[5] & Fhc7z6[29]);
assign Yoj6z6 = (Srj6z6 & Asj6z6);
assign Asj6z6 = (Isj6z6 & Qsj6z6);
assign Qsj6z6 = (Ysj6z6 & J1gov6);
assign J1gov6 = (!Bdu6x6);
assign Bdu6x6 = (Dte7z6[13] | Dte7z6[14]);
assign Ysj6z6 = (Fhc7z6[21] & Fhc7z6[13]);
assign Isj6z6 = (Oac7z6[2] & Oac7z6[3]);
assign Srj6z6 = (Gtj6z6 & Otj6z6);
assign Otj6z6 = (Oac7z6[0] & Oac7z6[1]);
assign Gtj6z6 = (Bqbdt6 & Qp07x6);
assign Qp07x6 = (Wtj6z6 & Dte7z6[15]);
assign Wtj6z6 = (~(Msziw6 | Dte7z6[16]));
assign Msziw6 = (!Dte7z6[17]);
assign Uij6z6 = (T3jhw6 & Ldo7v6);
assign Whj6z6 = (~(Jv0ov6 & Euj6z6));
assign Euj6z6 = (~(Muj6z6 & Uuj6z6));
assign Uuj6z6 = (Cvj6z6 & Kvj6z6);
assign Kvj6z6 = (~(Efcdt6 | A3ddt6));
assign Cvj6z6 = (Svj6z6 & U5u6x6);
assign U5u6x6 = (!X0wnv6);
assign X0wnv6 = (V5ddt6 & K3jnv6);
assign Svj6z6 = (~(Awj6z6 & Wzcdt6));
assign Awj6z6 = (Pacdt6 & Yiaov6);
assign Muj6z6 = (Iwj6z6 & K3jnv6);
assign Iwj6z6 = (Qwj6z6 & Ywj6z6);
assign Ywj6z6 = (~(Fjaov6 & Gxj6z6));
assign Gxj6z6 = (~(Oxj6z6 & Yiaov6));
assign Oxj6z6 = (Wxj6z6 & Fetov6);
assign Wxj6z6 = (~(Wzcdt6 & Eyj6z6));
assign Qwj6z6 = (~(Hofxx6 & Eyj6z6));
assign Eyj6z6 = (~(Myj6z6 & Uyj6z6));
assign Uyj6z6 = (Czj6z6 & Kzj6z6);
assign Kzj6z6 = (~(Szj6z6 & Isfxx6));
assign Isfxx6 = (D6tov6 & T7tov6);
assign T7tov6 = (!Bfd7z6[5]);
assign Szj6z6 = (Kbriy6 & J9tov6);
assign J9tov6 = (!Bfd7z6[1]);
assign Czj6z6 = (~(Mi77z6 | Zgadt6));
assign Myj6z6 = (Fccdt6 & A0k6z6);
assign A0k6z6 = (~(Hofxx6 & I0k6z6));
assign I0k6z6 = (~(Fjaov6 & Kd1ov6));
assign Kd1ov6 = (!Wzcdt6);
assign Hofxx6 = (G597z6 & Q0k6z6);
assign Q0k6z6 = (~(Y0k6z6 & G1k6z6));
assign G1k6z6 = (~(Pmc7z6[1] & O1k6z6));
assign Y0k6z6 = (~(W1k6z6 & Pmc7z6[2]));
assign Jv0ov6 = (!Af1ov6);
assign Af1ov6 = (~(Eu46z6 & E2k6z6));
assign Ygj6z6 = (~(Qmnov6 | Oznov6));
assign Igj6z6 = (M2k6z6 & U2k6z6);
assign U2k6z6 = (~(Znnov6 & Venov6));
assign M2k6z6 = (Sgcdt6 | C3k6z6);
assign C3k6z6 = (~(K3k6z6 | N9oov6));
assign HTRANSD[1] = (S3k6z6 & A4k6z6);
assign A4k6z6 = (~(I4k6z6 & Q4k6z6));
assign Q4k6z6 = (Ibonv6 | E2j6z6);
assign E2j6z6 = (~(Y4k6z6 | G5k6z6));
assign G5k6z6 = (Znn7z6[1] ? O5k6z6 : Xvgxx6);
assign O5k6z6 = (O3uet6 & Znn7z6[2]);
assign Y4k6z6 = (~(W5k6z6 & Eq0jy6));
assign W5k6z6 = (Xvgxx6 | Sjyet6);
assign HTRANSD[0] = (E6k6z6 & U2j6z6);
assign U2j6z6 = (Jc4iw6 & M6k6z6);
assign M6k6z6 = (!Iynet6);
assign Jc4iw6 = (~(U6k6z6 & C7k6z6));
assign C7k6z6 = (~(K7k6z6 & W13et6));
assign K7k6z6 = (~(S7k6z6 | Ex7et6));
assign S7k6z6 = (A8k6z6 & I8k6z6);
assign I8k6z6 = (~(Q8k6z6 & Igniy6));
assign Igniy6 = (~(Y8k6z6 & Xkr8v6));
assign Y8k6z6 = (Hir8v6 & Ycniy6);
assign Ycniy6 = (Dqr8v6 & Nnr8v6);
assign Q8k6z6 = (~(J8nov6 & G9k6z6));
assign J8nov6 = (Ojphw6 | Aga7z6);
assign U6k6z6 = (~(O9k6z6 & W9k6z6));
assign W9k6z6 = (Eak6z6 & Mak6z6);
assign Mak6z6 = (Rihhw6 | Pxmov6);
assign Pxmov6 = (!Hir8v6);
assign Rihhw6 = (Kihhw6 | Xkr8v6);
assign Kihhw6 = (~(Kpaov6 & Xlaov6));
assign Xlaov6 = (!Dqr8v6);
assign Kpaov6 = (!Nnr8v6);
assign Eak6z6 = (~(Aga7z6 | Ex7et6));
assign Aga7z6 = (!Lxydt6);
assign O9k6z6 = (Dihhw6 & W13et6);
assign E6k6z6 = (S3k6z6 & Hm1ov6);
assign S3k6z6 = (Uak6z6 & Cbk6z6);
assign Cbk6z6 = (~(Nhonv6 & Hm1ov6));
assign Uak6z6 = (~(Qmonv6 & Jn1ov6));
assign Qmonv6 = (Gmnet6 & Nhonv6);
assign Nhonv6 = (!B2jnv6);
assign HTMDHWDATA[9] = (~(Kbk6z6 & Sbk6z6));
assign Sbk6z6 = (Ack6z6 & Ick6z6);
assign Ick6z6 = (~(Qck6z6 & Jexmz6[1]));
assign Ack6z6 = (~(Yck6z6 & Jexmz6[25]));
assign Kbk6z6 = (Gdk6z6 & Odk6z6);
assign Odk6z6 = (~(Wdk6z6 & Jexmz6[17]));
assign Gdk6z6 = (~(Eek6z6 & Jexmz6[9]));
assign HTMDHWDATA[8] = (~(Mek6z6 & Uek6z6));
assign Uek6z6 = (Cfk6z6 & Kfk6z6);
assign Kfk6z6 = (~(Qck6z6 & Jexmz6[0]));
assign Cfk6z6 = (~(Yck6z6 & Jexmz6[24]));
assign Mek6z6 = (Sfk6z6 & Agk6z6);
assign Agk6z6 = (~(Wdk6z6 & Jexmz6[16]));
assign Sfk6z6 = (~(Eek6z6 & Jexmz6[8]));
assign HTMDHWDATA[7] = (~(Igk6z6 & Qgk6z6));
assign Qgk6z6 = (Ygk6z6 & Ghk6z6);
assign Ghk6z6 = (~(Qck6z6 & Jexmz6[31]));
assign Ygk6z6 = (~(Yck6z6 & Jexmz6[23]));
assign Igk6z6 = (Ohk6z6 & Whk6z6);
assign Whk6z6 = (~(Wdk6z6 & Jexmz6[15]));
assign Ohk6z6 = (~(Eek6z6 & Jexmz6[7]));
assign HTMDHWDATA[6] = (~(Eik6z6 & Mik6z6));
assign Mik6z6 = (Uik6z6 & Cjk6z6);
assign Cjk6z6 = (~(Qck6z6 & Jexmz6[30]));
assign Uik6z6 = (~(Yck6z6 & Jexmz6[22]));
assign Eik6z6 = (Kjk6z6 & Sjk6z6);
assign Sjk6z6 = (~(Wdk6z6 & Jexmz6[14]));
assign Kjk6z6 = (~(Eek6z6 & Jexmz6[6]));
assign HTMDHWDATA[5] = (~(Akk6z6 & Ikk6z6));
assign Ikk6z6 = (Qkk6z6 & Ykk6z6);
assign Ykk6z6 = (~(Qck6z6 & Jexmz6[29]));
assign Qkk6z6 = (~(Yck6z6 & Jexmz6[21]));
assign Akk6z6 = (Glk6z6 & Olk6z6);
assign Olk6z6 = (~(Wdk6z6 & Jexmz6[13]));
assign Glk6z6 = (~(Eek6z6 & Jexmz6[5]));
assign HTMDHWDATA[4] = (~(Wlk6z6 & Emk6z6));
assign Emk6z6 = (Mmk6z6 & Umk6z6);
assign Umk6z6 = (~(Qck6z6 & Jexmz6[28]));
assign Mmk6z6 = (~(Yck6z6 & Jexmz6[20]));
assign Wlk6z6 = (Cnk6z6 & Knk6z6);
assign Knk6z6 = (~(Wdk6z6 & Jexmz6[12]));
assign Cnk6z6 = (~(Eek6z6 & Jexmz6[4]));
assign HTMDHWDATA[3] = (~(Snk6z6 & Aok6z6));
assign Aok6z6 = (Iok6z6 & Qok6z6);
assign Qok6z6 = (~(Qck6z6 & Jexmz6[27]));
assign Iok6z6 = (~(Yck6z6 & Jexmz6[19]));
assign Snk6z6 = (Yok6z6 & Gpk6z6);
assign Gpk6z6 = (~(Wdk6z6 & Jexmz6[11]));
assign Yok6z6 = (~(Eek6z6 & Jexmz6[3]));
assign HTMDHWDATA[31] = (~(Opk6z6 & Wpk6z6));
assign Wpk6z6 = (Eqk6z6 & Mqk6z6);
assign Mqk6z6 = (~(Qck6z6 & Jexmz6[23]));
assign Eqk6z6 = (~(Yck6z6 & Jexmz6[15]));
assign Opk6z6 = (Uqk6z6 & Crk6z6);
assign Crk6z6 = (~(Wdk6z6 & Jexmz6[7]));
assign Uqk6z6 = (~(Eek6z6 & Jexmz6[31]));
assign HTMDHWDATA[30] = (~(Krk6z6 & Srk6z6));
assign Srk6z6 = (Ask6z6 & Isk6z6);
assign Isk6z6 = (~(Qck6z6 & Jexmz6[22]));
assign Ask6z6 = (~(Yck6z6 & Jexmz6[14]));
assign Krk6z6 = (Qsk6z6 & Ysk6z6);
assign Ysk6z6 = (~(Wdk6z6 & Jexmz6[6]));
assign Qsk6z6 = (~(Eek6z6 & Jexmz6[30]));
assign HTMDHWDATA[2] = (~(Gtk6z6 & Otk6z6));
assign Otk6z6 = (Wtk6z6 & Euk6z6);
assign Euk6z6 = (~(Qck6z6 & Jexmz6[26]));
assign Wtk6z6 = (~(Yck6z6 & Jexmz6[18]));
assign Gtk6z6 = (Muk6z6 & Uuk6z6);
assign Uuk6z6 = (~(Wdk6z6 & Jexmz6[10]));
assign Muk6z6 = (~(Eek6z6 & Jexmz6[2]));
assign HTMDHWDATA[29] = (~(Cvk6z6 & Kvk6z6));
assign Kvk6z6 = (Svk6z6 & Awk6z6);
assign Awk6z6 = (~(Qck6z6 & Jexmz6[21]));
assign Svk6z6 = (~(Yck6z6 & Jexmz6[13]));
assign Cvk6z6 = (Iwk6z6 & Qwk6z6);
assign Qwk6z6 = (~(Wdk6z6 & Jexmz6[5]));
assign Iwk6z6 = (~(Eek6z6 & Jexmz6[29]));
assign HTMDHWDATA[28] = (~(Ywk6z6 & Gxk6z6));
assign Gxk6z6 = (Oxk6z6 & Wxk6z6);
assign Wxk6z6 = (~(Qck6z6 & Jexmz6[20]));
assign Oxk6z6 = (~(Yck6z6 & Jexmz6[12]));
assign Ywk6z6 = (Eyk6z6 & Myk6z6);
assign Myk6z6 = (~(Wdk6z6 & Jexmz6[4]));
assign Eyk6z6 = (~(Eek6z6 & Jexmz6[28]));
assign HTMDHWDATA[27] = (~(Uyk6z6 & Czk6z6));
assign Czk6z6 = (Kzk6z6 & Szk6z6);
assign Szk6z6 = (~(Qck6z6 & Jexmz6[19]));
assign Kzk6z6 = (~(Yck6z6 & Jexmz6[11]));
assign Uyk6z6 = (A0l6z6 & I0l6z6);
assign I0l6z6 = (~(Wdk6z6 & Jexmz6[3]));
assign A0l6z6 = (~(Eek6z6 & Jexmz6[27]));
assign HTMDHWDATA[26] = (~(Q0l6z6 & Y0l6z6));
assign Y0l6z6 = (G1l6z6 & O1l6z6);
assign O1l6z6 = (~(Qck6z6 & Jexmz6[18]));
assign G1l6z6 = (~(Yck6z6 & Jexmz6[10]));
assign Q0l6z6 = (W1l6z6 & E2l6z6);
assign E2l6z6 = (~(Wdk6z6 & Jexmz6[2]));
assign W1l6z6 = (~(Eek6z6 & Jexmz6[26]));
assign HTMDHWDATA[25] = (~(M2l6z6 & U2l6z6));
assign U2l6z6 = (C3l6z6 & K3l6z6);
assign K3l6z6 = (~(Qck6z6 & Jexmz6[17]));
assign C3l6z6 = (~(Yck6z6 & Jexmz6[9]));
assign M2l6z6 = (S3l6z6 & A4l6z6);
assign A4l6z6 = (~(Wdk6z6 & Jexmz6[1]));
assign S3l6z6 = (~(Eek6z6 & Jexmz6[25]));
assign HTMDHWDATA[24] = (~(I4l6z6 & Q4l6z6));
assign Q4l6z6 = (Y4l6z6 & G5l6z6);
assign G5l6z6 = (~(Qck6z6 & Jexmz6[16]));
assign Y4l6z6 = (~(Yck6z6 & Jexmz6[8]));
assign I4l6z6 = (O5l6z6 & W5l6z6);
assign W5l6z6 = (~(Wdk6z6 & Jexmz6[0]));
assign O5l6z6 = (~(Eek6z6 & Jexmz6[24]));
assign HTMDHWDATA[23] = (~(E6l6z6 & M6l6z6));
assign M6l6z6 = (U6l6z6 & C7l6z6);
assign C7l6z6 = (~(Qck6z6 & Jexmz6[15]));
assign U6l6z6 = (~(Yck6z6 & Jexmz6[7]));
assign E6l6z6 = (K7l6z6 & S7l6z6);
assign S7l6z6 = (~(Wdk6z6 & Jexmz6[31]));
assign K7l6z6 = (~(Eek6z6 & Jexmz6[23]));
assign HTMDHWDATA[22] = (~(A8l6z6 & I8l6z6));
assign I8l6z6 = (Q8l6z6 & Y8l6z6);
assign Y8l6z6 = (~(Qck6z6 & Jexmz6[14]));
assign Q8l6z6 = (~(Yck6z6 & Jexmz6[6]));
assign A8l6z6 = (G9l6z6 & O9l6z6);
assign O9l6z6 = (~(Wdk6z6 & Jexmz6[30]));
assign G9l6z6 = (~(Eek6z6 & Jexmz6[22]));
assign HTMDHWDATA[21] = (~(W9l6z6 & Eal6z6));
assign Eal6z6 = (Mal6z6 & Ual6z6);
assign Ual6z6 = (~(Qck6z6 & Jexmz6[13]));
assign Mal6z6 = (~(Yck6z6 & Jexmz6[5]));
assign W9l6z6 = (Cbl6z6 & Kbl6z6);
assign Kbl6z6 = (~(Wdk6z6 & Jexmz6[29]));
assign Cbl6z6 = (~(Eek6z6 & Jexmz6[21]));
assign HTMDHWDATA[20] = (~(Sbl6z6 & Acl6z6));
assign Acl6z6 = (Icl6z6 & Qcl6z6);
assign Qcl6z6 = (~(Qck6z6 & Jexmz6[12]));
assign Icl6z6 = (~(Yck6z6 & Jexmz6[4]));
assign Sbl6z6 = (Ycl6z6 & Gdl6z6);
assign Gdl6z6 = (~(Wdk6z6 & Jexmz6[28]));
assign Ycl6z6 = (~(Eek6z6 & Jexmz6[20]));
assign HTMDHWDATA[1] = (~(Odl6z6 & Wdl6z6));
assign Wdl6z6 = (Eel6z6 & Mel6z6);
assign Mel6z6 = (~(Qck6z6 & Jexmz6[25]));
assign Eel6z6 = (~(Yck6z6 & Jexmz6[17]));
assign Odl6z6 = (Uel6z6 & Cfl6z6);
assign Cfl6z6 = (~(Wdk6z6 & Jexmz6[9]));
assign Uel6z6 = (~(Eek6z6 & Jexmz6[1]));
assign HTMDHWDATA[19] = (~(Kfl6z6 & Sfl6z6));
assign Sfl6z6 = (Agl6z6 & Igl6z6);
assign Igl6z6 = (~(Qck6z6 & Jexmz6[11]));
assign Agl6z6 = (~(Yck6z6 & Jexmz6[3]));
assign Kfl6z6 = (Qgl6z6 & Ygl6z6);
assign Ygl6z6 = (~(Wdk6z6 & Jexmz6[27]));
assign Qgl6z6 = (~(Eek6z6 & Jexmz6[19]));
assign HTMDHWDATA[18] = (~(Ghl6z6 & Ohl6z6));
assign Ohl6z6 = (Whl6z6 & Eil6z6);
assign Eil6z6 = (~(Qck6z6 & Jexmz6[10]));
assign Whl6z6 = (~(Yck6z6 & Jexmz6[2]));
assign Ghl6z6 = (Mil6z6 & Uil6z6);
assign Uil6z6 = (~(Wdk6z6 & Jexmz6[26]));
assign Mil6z6 = (~(Eek6z6 & Jexmz6[18]));
assign HTMDHWDATA[17] = (~(Cjl6z6 & Kjl6z6));
assign Kjl6z6 = (Sjl6z6 & Akl6z6);
assign Akl6z6 = (~(Qck6z6 & Jexmz6[9]));
assign Sjl6z6 = (~(Yck6z6 & Jexmz6[1]));
assign Cjl6z6 = (Ikl6z6 & Qkl6z6);
assign Qkl6z6 = (~(Wdk6z6 & Jexmz6[25]));
assign Ikl6z6 = (~(Eek6z6 & Jexmz6[17]));
assign HTMDHWDATA[16] = (~(Ykl6z6 & Gll6z6));
assign Gll6z6 = (Oll6z6 & Wll6z6);
assign Wll6z6 = (~(Qck6z6 & Jexmz6[8]));
assign Oll6z6 = (~(Yck6z6 & Jexmz6[0]));
assign Ykl6z6 = (Eml6z6 & Mml6z6);
assign Mml6z6 = (~(Wdk6z6 & Jexmz6[24]));
assign Eml6z6 = (~(Eek6z6 & Jexmz6[16]));
assign HTMDHWDATA[15] = (~(Uml6z6 & Cnl6z6));
assign Cnl6z6 = (Knl6z6 & Snl6z6);
assign Snl6z6 = (~(Qck6z6 & Jexmz6[7]));
assign Knl6z6 = (~(Yck6z6 & Jexmz6[31]));
assign Uml6z6 = (Aol6z6 & Iol6z6);
assign Iol6z6 = (~(Wdk6z6 & Jexmz6[23]));
assign Aol6z6 = (~(Eek6z6 & Jexmz6[15]));
assign HTMDHWDATA[14] = (~(Qol6z6 & Yol6z6));
assign Yol6z6 = (Gpl6z6 & Opl6z6);
assign Opl6z6 = (~(Qck6z6 & Jexmz6[6]));
assign Gpl6z6 = (~(Yck6z6 & Jexmz6[30]));
assign Qol6z6 = (Wpl6z6 & Eql6z6);
assign Eql6z6 = (~(Wdk6z6 & Jexmz6[22]));
assign Wpl6z6 = (~(Eek6z6 & Jexmz6[14]));
assign HTMDHWDATA[13] = (~(Mql6z6 & Uql6z6));
assign Uql6z6 = (Crl6z6 & Krl6z6);
assign Krl6z6 = (~(Qck6z6 & Jexmz6[5]));
assign Crl6z6 = (~(Yck6z6 & Jexmz6[29]));
assign Mql6z6 = (Srl6z6 & Asl6z6);
assign Asl6z6 = (~(Wdk6z6 & Jexmz6[21]));
assign Srl6z6 = (~(Eek6z6 & Jexmz6[13]));
assign HTMDHWDATA[12] = (~(Isl6z6 & Qsl6z6));
assign Qsl6z6 = (Ysl6z6 & Gtl6z6);
assign Gtl6z6 = (~(Qck6z6 & Jexmz6[4]));
assign Ysl6z6 = (~(Yck6z6 & Jexmz6[28]));
assign Isl6z6 = (Otl6z6 & Wtl6z6);
assign Wtl6z6 = (~(Wdk6z6 & Jexmz6[20]));
assign Otl6z6 = (~(Eek6z6 & Jexmz6[12]));
assign HTMDHWDATA[11] = (~(Eul6z6 & Mul6z6));
assign Mul6z6 = (Uul6z6 & Cvl6z6);
assign Cvl6z6 = (~(Qck6z6 & Jexmz6[3]));
assign Uul6z6 = (~(Yck6z6 & Jexmz6[27]));
assign Eul6z6 = (Kvl6z6 & Svl6z6);
assign Svl6z6 = (~(Wdk6z6 & Jexmz6[19]));
assign Kvl6z6 = (~(Eek6z6 & Jexmz6[11]));
assign HTMDHWDATA[10] = (~(Awl6z6 & Iwl6z6));
assign Iwl6z6 = (Qwl6z6 & Ywl6z6);
assign Ywl6z6 = (~(Qck6z6 & Jexmz6[2]));
assign Qwl6z6 = (~(Yck6z6 & Jexmz6[26]));
assign Awl6z6 = (Gxl6z6 & Oxl6z6);
assign Oxl6z6 = (~(Wdk6z6 & Jexmz6[18]));
assign Gxl6z6 = (~(Eek6z6 & Jexmz6[10]));
assign HTMDHWDATA[0] = (~(Wxl6z6 & Eyl6z6));
assign Eyl6z6 = (Myl6z6 & Uyl6z6);
assign Uyl6z6 = (~(Qck6z6 & Jexmz6[24]));
assign Qck6z6 = (~(Ue4iw6 | Ld4iw6));
assign Myl6z6 = (~(Yck6z6 & Jexmz6[16]));
assign Yck6z6 = (~(Ue4iw6 | Fb47v6));
assign Ue4iw6 = (!V947v6);
assign Wxl6z6 = (Czl6z6 & Kzl6z6);
assign Kzl6z6 = (~(Wdk6z6 & Jexmz6[8]));
assign Wdk6z6 = (~(Ld4iw6 | V947v6));
assign Ld4iw6 = (!Fb47v6);
assign Czl6z6 = (~(Eek6z6 & Jexmz6[0]));
assign Eek6z6 = (~(V947v6 | Fb47v6));
assign HSIZES[1] = (~(Szl6z6 & A0m6z6));
assign A0m6z6 = (~(J0jxx6 & I0m6z6));
assign I0m6z6 = (~(Q0m6z6 & Y0m6z6));
assign Q0m6z6 = (G1m6z6 & O1m6z6);
assign O1m6z6 = (~(Gsb7z6[1] & Xvgxx6));
assign G1m6z6 = (Jtonv6 | Vugxx6);
assign Jtonv6 = (!S7n7z6[1]);
assign Szl6z6 = (W1m6z6 & E2m6z6);
assign E2m6z6 = (~(M2m6z6 & Anehw6));
assign M2m6z6 = (~(U2m6z6 & C3m6z6));
assign C3m6z6 = (~(Rj9ov6 & Srhiy6));
assign W1m6z6 = (~(Hub7z6[1] & K3m6z6));
assign K3m6z6 = (~(En9ov6 & S3m6z6));
assign S3m6z6 = (~(Fk9ov6 & Jvdiw6));
assign HSIZES[0] = (~(A4m6z6 & I4m6z6));
assign I4m6z6 = (Q4m6z6 & Y4m6z6);
assign Y4m6z6 = (G5m6z6 | O5m6z6);
assign Q4m6z6 = (W5m6z6 & E6m6z6);
assign E6m6z6 = (~(Mma6z6 & M6m6z6));
assign W5m6z6 = (Uaonv6 | U6m6z6);
assign A4m6z6 = (C7m6z6 & K7m6z6);
assign K7m6z6 = (~(Zmnyx6 & Hub7z6[0]));
assign C7m6z6 = (~(S7m6z6 & Wbhnv6));
assign HSIZED[1] = (~(A8m6z6 & I8m6z6));
assign I8m6z6 = (~(Q8m6z6 & Vm1ov6));
assign Q8m6z6 = (Jvdiw6 & Hub7z6[1]);
assign A8m6z6 = (~(Y8m6z6 & Hm1ov6));
assign Y8m6z6 = (Srhiy6 & Anehw6);
assign HSIZED[0] = (~(G9m6z6 & O9m6z6));
assign O9m6z6 = (Jfonv6 | O5m6z6);
assign O5m6z6 = (W9m6z6 & Eam6z6);
assign Eam6z6 = (~(Mam6z6 & D94iw6));
assign W9m6z6 = (~(Wbhnv6 & Nxdiw6));
assign Wbhnv6 = (!Ta4iw6);
assign G9m6z6 = (Uam6z6 & Cbm6z6);
assign Cbm6z6 = (~(Vm1ov6 & M6m6z6));
assign M6m6z6 = (~(Rzdiw6 & Kbm6z6));
assign Kbm6z6 = (~(Sbm6z6 & Hub7z6[0]));
assign Uam6z6 = (Ibonv6 | U6m6z6);
assign U6m6z6 = (Acm6z6 & Icm6z6);
assign Icm6z6 = (~(S7n7z6[0] & Qo8iy6));
assign Acm6z6 = (Qcm6z6 & Ycm6z6);
assign Ycm6z6 = (~(Gdm6z6 & Znn7z6[1]));
assign Gdm6z6 = (~(Xvgxx6 | Eiliy6));
assign Eiliy6 = (Ven7z6[1] & I8liy6);
assign I8liy6 = (!Ven7z6[2]);
assign Qcm6z6 = (~(Gsb7z6[0] & Qakiw6));
assign HPROTS[3] = (~(Odm6z6 & Wdm6z6));
assign Wdm6z6 = (~(Rj9ov6 & Pgqnv6));
assign Pgqnv6 = (~(Eem6z6 & Mem6z6));
assign Mem6z6 = (~(K7a6z6 & Uem6z6));
assign Uem6z6 = (~(Cfm6z6 & Kja6z6));
assign Cfm6z6 = (Kfm6z6 & Sfm6z6);
assign Sfm6z6 = (~(Agm6z6 & Qga6z6));
assign Agm6z6 = (Cba6z6 & Igm6z6);
assign Eem6z6 = (Qgm6z6 & Eia6z6);
assign Eia6z6 = (~(Ygm6z6 & Ghm6z6));
assign Ghm6z6 = (I4a6z6 ? Ohm6z6 : E6a6z6);
assign Ygm6z6 = (Q4a6z6 & M6a6z6);
assign Qgm6z6 = (~(Q4a6z6 & Whm6z6));
assign Whm6z6 = (~(Eim6z6 & Mim6z6));
assign Mim6z6 = (~(Uim6z6 & Cmm7z6[29]));
assign Uim6z6 = (Rygnv6 & I4a6z6);
assign Eim6z6 = (M6a6z6 | V5k7z6[31]);
assign Odm6z6 = (~(Qtoet6 & J0jxx6));
assign HPROTS[2] = (~(Cjm6z6 & Kjm6z6));
assign Kjm6z6 = (~(Rj9ov6 & Yhqnv6));
assign Yhqnv6 = (~(Sjm6z6 & Akm6z6));
assign Akm6z6 = (~(Ikm6z6 & Q4a6z6));
assign Q4a6z6 = (!U6a6z6);
assign U6a6z6 = (~(Qkm6z6 & Uia6z6));
assign Qkm6z6 = (~(Sjy5z6 & Ykm6z6));
assign Ykm6z6 = (~(Apget6 & Glm6z6));
assign Ikm6z6 = (P1het6 ? Wlm6z6 : Olm6z6);
assign Wlm6z6 = (Emm6z6 & Mmm6z6);
assign Mmm6z6 = (~(Umm6z6 & Cnm6z6));
assign Cnm6z6 = (Knm6z6 & Snm6z6);
assign Knm6z6 = (~(V5k7z6[18] | V5k7z6[19]));
assign Umm6z6 = (~(Jhdiw6 | Aom6z6));
assign Jhdiw6 = (!Ui77z6);
assign Emm6z6 = (V5k7z6[29] | V5k7z6[30]);
assign Olm6z6 = (Lgonv6 & Iom6z6);
assign Sjm6z6 = (~(K7a6z6 & Qom6z6));
assign Qom6z6 = (~(Yom6z6 & Gpm6z6));
assign Gpm6z6 = (~(Kba6z6 & Yga6z6));
assign Yga6z6 = (!Cba6z6);
assign Cba6z6 = (Opm6z6 & Wpm6z6);
assign Wpm6z6 = (Eqm6z6 & Mqm6z6);
assign Mqm6z6 = (Uqm6z6 & Crm6z6);
assign Crm6z6 = (~(Zlk7z6[18] & Uea6z6));
assign Uqm6z6 = (~(Hwk7z6[18] & Sba6z6));
assign Eqm6z6 = (Krm6z6 & Srm6z6);
assign Srm6z6 = (~(Frl7z6[18] & Yca6z6));
assign Krm6z6 = (~(Xgl7z6[18] & Qca6z6));
assign Opm6z6 = (Asm6z6 & Ism6z6);
assign Ism6z6 = (Qsm6z6 & Ysm6z6);
assign Ysm6z6 = (~(Vbm7z6[18] & Aga6z6));
assign Qsm6z6 = (~(Rbk7z6[18] & Sfa6z6));
assign Asm6z6 = (Gtm6z6 & Otm6z6);
assign Otm6z6 = (~(N1m7z6[18] & Mea6z6));
assign Gtm6z6 = (~(P6l7z6[18] & Eaa6z6));
assign Kba6z6 = (Wtm6z6 & Kja6z6);
assign Wtm6z6 = (Kfm6z6 & Aka6z6);
assign Kfm6z6 = (!Ika6z6);
assign Ika6z6 = (~(Eum6z6 & Mum6z6));
assign Mum6z6 = (Uum6z6 & Cvm6z6);
assign Cvm6z6 = (Kvm6z6 & Svm6z6);
assign Svm6z6 = (~(Rbk7z6[15] & Sfa6z6));
assign Kvm6z6 = (~(Hwk7z6[15] & Sba6z6));
assign Uum6z6 = (Awm6z6 & Iwm6z6);
assign Iwm6z6 = (~(Frl7z6[15] & Yca6z6));
assign Awm6z6 = (~(Xgl7z6[15] & Qca6z6));
assign Eum6z6 = (Qwm6z6 & Ywm6z6);
assign Ywm6z6 = (Gxm6z6 & Oxm6z6);
assign Oxm6z6 = (~(Vbm7z6[15] & Aga6z6));
assign Gxm6z6 = (~(P6l7z6[15] & Eaa6z6));
assign Qwm6z6 = (Wxm6z6 & Eym6z6);
assign Eym6z6 = (~(Zlk7z6[15] & Uea6z6));
assign Wxm6z6 = (~(N1m7z6[15] & Mea6z6));
assign Yom6z6 = (Kja6z6 ? Qga6z6 : Aka6z6);
assign Kja6z6 = (Mym6z6 & Uym6z6);
assign Uym6z6 = (Czm6z6 & Kzm6z6);
assign Kzm6z6 = (Szm6z6 & A0n6z6);
assign A0n6z6 = (~(Zlk7z6[19] & Uea6z6));
assign Szm6z6 = (~(Hwk7z6[19] & Sba6z6));
assign Czm6z6 = (I0n6z6 & Q0n6z6);
assign Q0n6z6 = (~(Frl7z6[19] & Yca6z6));
assign I0n6z6 = (~(Xgl7z6[19] & Qca6z6));
assign Mym6z6 = (Y0n6z6 & G1n6z6);
assign G1n6z6 = (O1n6z6 & W1n6z6);
assign W1n6z6 = (~(Vbm7z6[19] & Aga6z6));
assign O1n6z6 = (~(Rbk7z6[19] & Sfa6z6));
assign Y0n6z6 = (E2n6z6 & M2n6z6);
assign M2n6z6 = (~(N1m7z6[19] & Mea6z6));
assign E2n6z6 = (~(P6l7z6[19] & Eaa6z6));
assign Qga6z6 = (U2n6z6 & C3n6z6);
assign C3n6z6 = (K3n6z6 & S3n6z6);
assign S3n6z6 = (A4n6z6 & I4n6z6);
assign I4n6z6 = (~(Rbk7z6[14] & Sfa6z6));
assign A4n6z6 = (~(Hwk7z6[14] & Sba6z6));
assign K3n6z6 = (Q4n6z6 & Y4n6z6);
assign Y4n6z6 = (~(Frl7z6[14] & Yca6z6));
assign Q4n6z6 = (~(Xgl7z6[14] & Qca6z6));
assign U2n6z6 = (G5n6z6 & O5n6z6);
assign O5n6z6 = (W5n6z6 & E6n6z6);
assign E6n6z6 = (~(Vbm7z6[14] & Aga6z6));
assign W5n6z6 = (~(P6l7z6[14] & Eaa6z6));
assign G5n6z6 = (M6n6z6 & U6n6z6);
assign U6n6z6 = (~(Zlk7z6[14] & Uea6z6));
assign M6n6z6 = (~(N1m7z6[14] & Mea6z6));
assign Aka6z6 = (!Igm6z6);
assign Igm6z6 = (~(C7n6z6 & K7n6z6));
assign K7n6z6 = (S7n6z6 & A8n6z6);
assign A8n6z6 = (I8n6z6 & Q8n6z6);
assign Q8n6z6 = (~(Hwk7z6[17] & Sba6z6));
assign I8n6z6 = (~(P6l7z6[17] & Eaa6z6));
assign S7n6z6 = (Y8n6z6 & G9n6z6);
assign G9n6z6 = (~(Xgl7z6[17] & Qca6z6));
assign Qca6z6 = (O9n6z6 & W9n6z6);
assign O9n6z6 = (Ean6z6 & Man6z6);
assign Y8n6z6 = (~(Frl7z6[17] & Yca6z6));
assign Yca6z6 = (~(Man6z6 | Uan6z6));
assign Uan6z6 = (!W9n6z6);
assign C7n6z6 = (Cbn6z6 & Kbn6z6);
assign Kbn6z6 = (Sbn6z6 & Acn6z6);
assign Acn6z6 = (~(N1m7z6[17] & Mea6z6));
assign Sbn6z6 = (~(Zlk7z6[17] & Uea6z6));
assign Uea6z6 = (Icn6z6 & Qcn6z6);
assign Icn6z6 = (~(Ean6z6 | Ycn6z6));
assign Cbn6z6 = (Gdn6z6 & Odn6z6);
assign Odn6z6 = (~(Rbk7z6[17] & Sfa6z6));
assign Gdn6z6 = (~(Vbm7z6[17] & Aga6z6));
assign K7a6z6 = (!Uia6z6);
assign Uia6z6 = (~(Wdn6z6 & Een6z6));
assign Wdn6z6 = (I4a6z6 ? Lgonv6 : Aom6z6);
assign Cjm6z6 = (~(Rvoet6 & J0jxx6));
assign HPROTS[1] = (~(Men6z6 & Uen6z6));
assign Uen6z6 = (~(Sxoet6 & J0jxx6));
assign Men6z6 = (Cfn6z6 & Kfn6z6);
assign Kfn6z6 = (~(Rj9ov6 & Hjqnv6));
assign Cfn6z6 = (~(K2bdt6 & Fk9ov6));
assign HPROTS[0] = (~(O1j6z6 & Sfn6z6));
assign Sfn6z6 = (~(Tzoet6 & J0jxx6));
assign O1j6z6 = (Cfonv6 & Zn9ov6);
assign HPROTI[1] = (Crcdt6 ? Fsc7z6[1] : Ghnov6);
assign Ghnov6 = (~(Gbo6x6 & Agn6z6));
assign Agn6z6 = (Xbmyx6 | Bpnov6);
assign Bpnov6 = (!Hkoov6);
assign Hkoov6 = (~(Ign6z6 & T3jhw6));
assign Ign6z6 = (Cgc7z6[2] & P1piw6);
assign Xbmyx6 = (~(Iooov6 & Lqfxx6));
assign Lqfxx6 = (~(Qloov6 & T3jhw6));
assign T3jhw6 = (~(O4jhw6 | Cgc7z6[3]));
assign Qloov6 = (Cgc7z6[2] & Cgc7z6[1]);
assign HPROTD[1] = (~(Qgn6z6 & Ygn6z6));
assign Ygn6z6 = (~(Sxoet6 & Jn1ov6));
assign Qgn6z6 = (Ghn6z6 & Ohn6z6);
assign Ohn6z6 = (~(Hm1ov6 & Hjqnv6));
assign Ghn6z6 = (~(K2bdt6 & Vm1ov6));
assign HPROTD[0] = (~(I4k6z6 & Whn6z6));
assign Whn6z6 = (~(Tzoet6 & Jn1ov6));
assign I4k6z6 = (Jfonv6 & V4myx6);
assign HMASTLOCKS = (~(T9nyx6 & Luixx6));
assign T9nyx6 = (Ein6z6 & Min6z6);
assign Min6z6 = (~(Ngnyx6 & Lhmov6));
assign Ngnyx6 = (S7m6z6 & B2jnv6);
assign B2jnv6 = (~(Uin6z6 & Senet6));
assign Uin6z6 = (Mfdiw6 & K9h7v6);
assign Mfdiw6 = (Tfdiw6 | Bkdiw6);
assign Bkdiw6 = (Cjn6z6 & Kjn6z6);
assign Kjn6z6 = (Sjn6z6 & Lgonv6);
assign Sjn6z6 = (Vb4iw6 & I4a6z6);
assign Cjn6z6 = (Akn6z6 & Ikn6z6);
assign Ikn6z6 = (~(Qkn6z6 & Ikoiy6));
assign Qkn6z6 = (Apget6 & Hjqnv6);
assign Tfdiw6 = (Ykn6z6 & Gln6z6);
assign Gln6z6 = (Oln6z6 & Aom6z6);
assign Aom6z6 = (~(Wln6z6 & Emn6z6));
assign Emn6z6 = (Mmn6z6 & Umn6z6);
assign Umn6z6 = (Cnn6z6 & Knn6z6);
assign Cnn6z6 = (~(V5k7z6[27] | V5k7z6[28]));
assign Mmn6z6 = (Snn6z6 & Aon6z6);
assign Snn6z6 = (~(V5k7z6[22] | V5k7z6[24]));
assign Wln6z6 = (Ion6z6 & Qon6z6);
assign Qon6z6 = (Yon6z6 & V5k7z6[31]);
assign Yon6z6 = (V5k7z6[29] & V5k7z6[30]);
assign Ion6z6 = (Gpn6z6 & Cj77z6);
assign Gpn6z6 = (Kj77z6 & U297z6);
assign Oln6z6 = (~(Opn6z6 & Dzget6));
assign Opn6z6 = (Ikoiy6 & Apget6);
assign Ikoiy6 = (!Een6z6);
assign Ykn6z6 = (Akn6z6 & P1het6);
assign Akn6z6 = (Sjy5z6 & Wpn6z6);
assign Wpn6z6 = (~(Eqn6z6 & Mqn6z6));
assign Mqn6z6 = (Uqn6z6 & Crn6z6);
assign Crn6z6 = (~(Eaa6z6 & Krn6z6));
assign Krn6z6 = (~(Srn6z6 & Asn6z6));
assign Asn6z6 = (P6l7z6[22] ? Qsn6z6 : Isn6z6);
assign Qsn6z6 = (~(Ysn6z6 & Isn6z6));
assign Isn6z6 = (P6l7z6[21] | P6l7z6[20]);
assign Srn6z6 = (P6l7z6[21] ? Otn6z6 : Gtn6z6);
assign Otn6z6 = (Wtn6z6 | P6l7z6[20]);
assign Gtn6z6 = (~(P6l7z6[20] & Eun6z6));
assign Eaa6z6 = (~(Mun6z6 | Uun6z6));
assign Mun6z6 = (!Cvn6z6);
assign Uqn6z6 = (Kvn6z6 & Een6z6);
assign Een6z6 = (~(Sfa6z6 & Svn6z6));
assign Svn6z6 = (~(Awn6z6 & Iwn6z6));
assign Iwn6z6 = (Qwn6z6 & Ywn6z6);
assign Ywn6z6 = (Gxn6z6 & Oxn6z6);
assign Oxn6z6 = (Wxn6z6 & Eyn6z6);
assign Eyn6z6 = (~(Cihet6 | Myn6z6));
assign Myn6z6 = (Uyn6z6 & Jienv6);
assign Jienv6 = (Czn6z6 & Kzn6z6);
assign Czn6z6 = (Szn6z6 & A0o6z6);
assign Uyn6z6 = (Ak4nv6 ^ Aoy5z6);
assign Aoy5z6 = (!Dfk7z6[5]);
assign Wxn6z6 = (I0o6z6 & Q0o6z6);
assign Q0o6z6 = (~(Y0o6z6 & O3env6));
assign O3env6 = (G1o6z6 | Cbenv6);
assign G1o6z6 = (Kzn6z6 & A0o6z6);
assign Y0o6z6 = (Dfk7z6[7] ^ Tp5nv6);
assign I0o6z6 = (~(Cbenv6 & O1o6z6));
assign O1o6z6 = (Dfk7z6[6] ^ Kv5nv6);
assign Cbenv6 = (Cienv6 & Szn6z6);
assign Gxn6z6 = (W1o6z6 & E2o6z6);
assign E2o6z6 = (M2o6z6 & U2o6z6);
assign U2o6z6 = (~(C3o6z6 & Nrenv6));
assign Nrenv6 = (Qwenv6 | Kzn6z6);
assign C3o6z6 = (Dfk7z6[15] ^ Je4nv6);
assign M2o6z6 = (~(K3o6z6 & Qwenv6));
assign Qwenv6 = (~(X4env6 & S3o6z6));
assign S3o6z6 = (~(Szn6z6 & Dmenv6));
assign X4env6 = (!H3env6);
assign K3o6z6 = (Dfk7z6[14] ^ Jl4nv6);
assign W1o6z6 = (A4o6z6 & I4o6z6);
assign I4o6z6 = (~(Q4o6z6 & H3env6));
assign H3env6 = (~(Lcenv6 & Y4o6z6));
assign Y4o6z6 = (~(Kzn6z6 & Szn6z6));
assign Lcenv6 = (!Vaenv6);
assign Q4o6z6 = (Dfk7z6[13] ^ Q74nv6);
assign A4o6z6 = (~(G5o6z6 & Vaenv6));
assign Vaenv6 = (~(Zjenv6 & O5o6z6));
assign O5o6z6 = (~(W5o6z6 & Dmenv6));
assign Zjenv6 = (!Qienv6);
assign G5o6z6 = (Dfk7z6[12] ^ Ce4nv6);
assign Qwn6z6 = (E6o6z6 & M6o6z6);
assign M6o6z6 = (U6o6z6 & C7o6z6);
assign C7o6z6 = (K7o6z6 & S7o6z6);
assign S7o6z6 = (~(A8o6z6 & Qienv6));
assign Qienv6 = (~(A3env6 & I8o6z6));
assign I8o6z6 = (~(Kzn6z6 & W5o6z6));
assign A3env6 = (!Fnenv6);
assign A8o6z6 = (Dfk7z6[11] ^ Cl4nv6);
assign K7o6z6 = (~(Q8o6z6 & Fnenv6));
assign Fnenv6 = (~(Oaenv6 & Y8o6z6));
assign Y8o6z6 = (~(G9o6z6 & Dmenv6));
assign Oaenv6 = (!Awy5z6);
assign Q8o6z6 = (Dfk7z6[10] ^ H64nv6);
assign U6o6z6 = (O9o6z6 & W9o6z6);
assign W9o6z6 = (~(Eao6z6 & Awy5z6));
assign Awy5z6 = (~(Mao6z6 & Pzenv6));
assign Pzenv6 = (!Cienv6);
assign Mao6z6 = (~(G9o6z6 & Kzn6z6));
assign Kzn6z6 = (Uao6z6 & Dmenv6);
assign Eao6z6 = (Dfk7z6[9] ^ Hd4nv6);
assign O9o6z6 = (~(Cienv6 & Cbo6z6));
assign Cbo6z6 = (Dfk7z6[8] ^ Hk4nv6);
assign Cienv6 = (A0o6z6 & Dmenv6);
assign E6o6z6 = (Kbo6z6 & Sbo6z6);
assign Sbo6z6 = (~(Aco6z6 & Peenv6));
assign Aco6z6 = (Ico6z6 ^ Dfk7z6[29]);
assign Kbo6z6 = (Qco6z6 & Yco6z6);
assign Yco6z6 = (~(Gdo6z6 & Nzdnv6));
assign Nzdnv6 = (!Jpenv6);
assign Jpenv6 = (Tuenv6 & Odo6z6);
assign Gdo6z6 = (~(Dfk7z6[31] ^ W34nv6));
assign Qco6z6 = (~(Wdo6z6 & B7env6));
assign B7env6 = (!Tuenv6);
assign Tuenv6 = (D0fnv6 & Eeo6z6);
assign D0fnv6 = (!Peenv6);
assign Peenv6 = (~(Gzdnv6 & Meo6z6));
assign Meo6z6 = (~(Szn6z6 & Uao6z6));
assign Wdo6z6 = (~(Dfk7z6[30] ^ Pa4nv6));
assign Awn6z6 = (Ueo6z6 & Cfo6z6);
assign Cfo6z6 = (Kfo6z6 & Sfo6z6);
assign Sfo6z6 = (Ago6z6 & Igo6z6);
assign Igo6z6 = (Qgo6z6 & Ygo6z6);
assign Ygo6z6 = (~(Gho6z6 & O1z5z6));
assign O1z5z6 = (!Gzdnv6);
assign Gzdnv6 = (Rbk7z6[3] & U6env6);
assign U6env6 = (!Dtenv6);
assign Gho6z6 = (Dfk7z6[28] ^ U24nv6);
assign Qgo6z6 = (~(Oho6z6 & Dtenv6));
assign Dtenv6 = (~(Ieenv6 & Who6z6));
assign Who6z6 = (~(W5o6z6 & Uao6z6));
assign Oho6z6 = (Dfk7z6[27] ^ U94nv6);
assign Ago6z6 = (Eio6z6 & Mio6z6);
assign Mio6z6 = (~(Uio6z6 & K0fnv6));
assign K0fnv6 = (!Ieenv6);
assign Ieenv6 = (Uzdnv6 & Cjo6z6);
assign Cjo6z6 = (!G9o6z6);
assign Uzdnv6 = (!K1env6);
assign Uio6z6 = (~(Dfk7z6[26] ^ Ng4nv6));
assign Eio6z6 = (~(Kjo6z6 & K1env6));
assign K1env6 = (~(I7env6 & Sjo6z6));
assign Sjo6z6 = (~(G9o6z6 & Uao6z6));
assign Kjo6z6 = (~(Dfk7z6[25] ^ B34nv6));
assign Kfo6z6 = (Ako6z6 & Iko6z6);
assign Iko6z6 = (~(Qko6z6 & Wlenv6));
assign Qko6z6 = (Dfk7z6[22] ^ Y44nv6);
assign Ako6z6 = (Yko6z6 & Glo6z6);
assign Glo6z6 = (~(Olo6z6 & Y8env6));
assign Y8env6 = (!I7env6);
assign I7env6 = (Weenv6 & Wlo6z6);
assign Olo6z6 = (Dfk7z6[24] ^ N94nv6);
assign Yko6z6 = (~(Emo6z6 & Mgenv6));
assign Mgenv6 = (!Weenv6);
assign Weenv6 = (~(Wlenv6 | Mmo6z6));
assign Wlenv6 = (~(R8env6 & Umo6z6));
assign Umo6z6 = (~(Szn6z6 & A0o6z6));
assign R8env6 = (!Grenv6);
assign Emo6z6 = (~(Dfk7z6[23] ^ Gg4nv6));
assign Ueo6z6 = (Cno6z6 & Kno6z6);
assign Kno6z6 = (Sno6z6 & Aoo6z6);
assign Aoo6z6 = (Ioo6z6 & Qoo6z6);
assign Qoo6z6 = (~(Yoo6z6 & Grenv6));
assign Grenv6 = (~(Fgenv6 & Gpo6z6));
assign Gpo6z6 = (~(Mmo6z6 & Szn6z6));
assign Fgenv6 = (!Gyenv6);
assign Yoo6z6 = (~(Dfk7z6[21] ^ Kb4nv6));
assign Ioo6z6 = (~(Opo6z6 & Gyenv6));
assign Gyenv6 = (~(R1env6 & Wpo6z6));
assign Wpo6z6 = (~(W5o6z6 & A0o6z6));
assign R1env6 = (!Q4env6);
assign Opo6z6 = (~(Dfk7z6[20] ^ Ri4nv6));
assign Sno6z6 = (Eqo6z6 & Mqo6z6);
assign Mqo6z6 = (~(Uqo6z6 & Q4env6));
assign Q4env6 = (~(F9env6 & Cro6z6));
assign Cro6z6 = (~(Mmo6z6 & W5o6z6));
assign F9env6 = (!Ecenv6);
assign Uqo6z6 = (Dfk7z6[19] ^ R44nv6);
assign Eqo6z6 = (~(Kro6z6 & Ecenv6));
assign Ecenv6 = (~(Tgenv6 & Sro6z6));
assign Sro6z6 = (~(G9o6z6 & A0o6z6));
assign Tgenv6 = (!Sjenv6);
assign Kro6z6 = (Dfk7z6[18] ^ Rb4nv6);
assign Cno6z6 = (Aso6z6 & O9z5z6);
assign Aso6z6 = (Iso6z6 & Qso6z6);
assign Qso6z6 = (~(Yso6z6 & Sjenv6));
assign Sjenv6 = (~(J4env6 & Gto6z6));
assign Gto6z6 = (~(Mmo6z6 & G9o6z6));
assign G9o6z6 = (Szn6z6 & W5o6z6);
assign Szn6z6 = (!Eeo6z6);
assign Eeo6z6 = (Rbk7z6[2] & O9z5z6);
assign Mmo6z6 = (Uao6z6 & A0o6z6);
assign A0o6z6 = (!Wlo6z6);
assign Wlo6z6 = (Rbk7z6[4] & O9z5z6);
assign Uao6z6 = (!Odo6z6);
assign Odo6z6 = (Rbk7z6[1] & O9z5z6);
assign Yso6z6 = (~(Dfk7z6[17] ^ Ki4nv6));
assign Iso6z6 = (~(Oto6z6 & Dmenv6));
assign Dmenv6 = (!J4env6);
assign J4env6 = (Rbk7z6[5] & O9z5z6);
assign O9z5z6 = (Wto6z6 & Rbk7z6[0]);
assign Wto6z6 = (Sjy5z6 & Euo6z6);
assign Euo6z6 = (~(Xafnv6 & W5o6z6));
assign W5o6z6 = (!Rbk7z6[3]);
assign Xafnv6 = (Muo6z6 & Uuo6z6);
assign Uuo6z6 = (!Rbk7z6[5]);
assign Muo6z6 = (!Rbk7z6[4]);
assign Oto6z6 = (~(Dfk7z6[16] ^ J74nv6));
assign Sfa6z6 = (~(Cvo6z6 | Ean6z6));
assign Cvo6z6 = (Ycn6z6 | Qcn6z6);
assign Ycn6z6 = (!Kvo6z6);
assign Kvn6z6 = (~(Sba6z6 & Svo6z6));
assign Svo6z6 = (~(Awo6z6 & Iwo6z6));
assign Iwo6z6 = (Hwk7z6[22] ? Ywo6z6 : Qwo6z6);
assign Ywo6z6 = (~(Ysn6z6 & Qwo6z6));
assign Qwo6z6 = (Hwk7z6[21] | Hwk7z6[20]);
assign Awo6z6 = (Hwk7z6[21] ? Oxo6z6 : Gxo6z6);
assign Oxo6z6 = (Wtn6z6 | Hwk7z6[20]);
assign Gxo6z6 = (~(Hwk7z6[20] & Eun6z6));
assign Sba6z6 = (~(Uun6z6 | Cvn6z6));
assign Uun6z6 = (Ean6z6 | Kvo6z6);
assign Eqn6z6 = (Wxo6z6 & Eyo6z6);
assign Eyo6z6 = (Ean6z6 ? Uyo6z6 : Myo6z6);
assign Ean6z6 = (~(Czo6z6 & W9n6z6));
assign Czo6z6 = (Kzo6z6 & Man6z6);
assign Kzo6z6 = (~(Szo6z6 & A0p6z6));
assign A0p6z6 = (I0p6z6 & Q0p6z6);
assign Q0p6z6 = (Y0p6z6 & G1p6z6);
assign G1p6z6 = (O1p6z6 & W1p6z6);
assign W1p6z6 = (~(Cmket6 | E2p6z6));
assign E2p6z6 = (M2p6z6 & Pk8nv6);
assign Pk8nv6 = (U2p6z6 & C3p6z6);
assign U2p6z6 = (K3p6z6 & S3p6z6);
assign M2p6z6 = (Ak4nv6 ^ Op06z6);
assign Op06z6 = (!Jkl7z6[5]);
assign O1p6z6 = (A4p6z6 & I4p6z6);
assign I4p6z6 = (~(Q4p6z6 & U58nv6));
assign U58nv6 = (Y4p6z6 | Id8nv6);
assign Y4p6z6 = (C3p6z6 & S3p6z6);
assign Q4p6z6 = (Uq06z6 ^ O64nv6);
assign O64nv6 = (!Tp5nv6);
assign Uq06z6 = (!Jkl7z6[7]);
assign A4p6z6 = (~(Id8nv6 & G5p6z6));
assign G5p6z6 = (Kr06z6 ^ Ad4nv6);
assign Ad4nv6 = (!Kv5nv6);
assign Kr06z6 = (!Jkl7z6[6]);
assign Id8nv6 = (Ik8nv6 & K3p6z6);
assign Y0p6z6 = (O5p6z6 & W5p6z6);
assign W5p6z6 = (E6p6z6 & M6p6z6);
assign M6p6z6 = (~(U6p6z6 & Tt8nv6));
assign Tt8nv6 = (Wy8nv6 | C3p6z6);
assign U6p6z6 = (Ot06z6 ^ C7p6z6);
assign C7p6z6 = (!Je4nv6);
assign Ot06z6 = (!Jkl7z6[15]);
assign E6p6z6 = (~(K7p6z6 & Wy8nv6));
assign Wy8nv6 = (~(D78nv6 & S7p6z6));
assign S7p6z6 = (~(K3p6z6 & Jo8nv6));
assign D78nv6 = (!N58nv6);
assign K7p6z6 = (Mu06z6 ^ A8p6z6);
assign A8p6z6 = (!Jl4nv6);
assign Mu06z6 = (!Jkl7z6[14]);
assign O5p6z6 = (I8p6z6 & Q8p6z6);
assign Q8p6z6 = (~(Y8p6z6 & N58nv6));
assign N58nv6 = (~(Re8nv6 & G9p6z6));
assign G9p6z6 = (~(C3p6z6 & K3p6z6));
assign Re8nv6 = (!Bd8nv6);
assign Y8p6z6 = (Aw06z6 ^ O9p6z6);
assign O9p6z6 = (!Q74nv6);
assign Aw06z6 = (!Jkl7z6[13]);
assign I8p6z6 = (~(W9p6z6 & Bd8nv6));
assign Bd8nv6 = (~(Fm8nv6 & Eap6z6));
assign Eap6z6 = (~(Map6z6 & Jo8nv6));
assign Fm8nv6 = (!Wk8nv6);
assign W9p6z6 = (Yw06z6 ^ Uap6z6);
assign Uap6z6 = (!Ce4nv6);
assign Yw06z6 = (!Jkl7z6[12]);
assign I0p6z6 = (Cbp6z6 & Kbp6z6);
assign Kbp6z6 = (Sbp6z6 & Acp6z6);
assign Acp6z6 = (Icp6z6 & Qcp6z6);
assign Qcp6z6 = (~(Ycp6z6 & Wk8nv6));
assign Wk8nv6 = (~(G58nv6 & Gdp6z6));
assign Gdp6z6 = (~(C3p6z6 & Map6z6));
assign G58nv6 = (!Lp8nv6);
assign Ycp6z6 = (Sz06z6 ^ Odp6z6);
assign Odp6z6 = (!Cl4nv6);
assign Sz06z6 = (!Jkl7z6[11]);
assign Icp6z6 = (~(Wdp6z6 & Lp8nv6));
assign Lp8nv6 = (~(Uc8nv6 & Eep6z6));
assign Eep6z6 = (~(Mep6z6 & Jo8nv6));
assign Uc8nv6 = (!W116z6);
assign Wdp6z6 = (Q016z6 ^ Uep6z6);
assign Uep6z6 = (!H64nv6);
assign Q016z6 = (!Jkl7z6[10]);
assign Sbp6z6 = (Cfp6z6 & Kfp6z6);
assign Kfp6z6 = (~(Sfp6z6 & W116z6));
assign W116z6 = (~(Agp6z6 & V19nv6));
assign V19nv6 = (!Ik8nv6);
assign Agp6z6 = (~(Mep6z6 & C3p6z6));
assign C3p6z6 = (Igp6z6 & Jo8nv6);
assign Sfp6z6 = (M216z6 ^ Qgp6z6);
assign Qgp6z6 = (!Hd4nv6);
assign M216z6 = (!Jkl7z6[9]);
assign Cfp6z6 = (~(Ik8nv6 & Ygp6z6));
assign Ygp6z6 = (C316z6 ^ Ghp6z6);
assign C316z6 = (!Jkl7z6[8]);
assign Ik8nv6 = (S3p6z6 & Jo8nv6);
assign Cbp6z6 = (Ohp6z6 & Whp6z6);
assign Whp6z6 = (~(Eip6z6 & Vg8nv6));
assign Eip6z6 = (Ph4nv6 ^ I416z6);
assign I416z6 = (!Jkl7z6[29]);
assign Ph4nv6 = (!Ico6z6);
assign Ohp6z6 = (Mip6z6 & Uip6z6);
assign Uip6z6 = (~(Cjp6z6 & T18nv6));
assign T18nv6 = (!Pr8nv6);
assign Pr8nv6 = (Zw8nv6 & Kjp6z6);
assign Cjp6z6 = (O516z6 ^ W34nv6);
assign O516z6 = (!Jkl7z6[31]);
assign Mip6z6 = (~(Sjp6z6 & H98nv6));
assign H98nv6 = (!Zw8nv6);
assign Zw8nv6 = (J29nv6 & Akp6z6);
assign J29nv6 = (!Vg8nv6);
assign Vg8nv6 = (~(M18nv6 & Ikp6z6));
assign Ikp6z6 = (~(K3p6z6 & Igp6z6));
assign Sjp6z6 = (E616z6 ^ Pa4nv6);
assign E616z6 = (!Jkl7z6[30]);
assign Szo6z6 = (Qkp6z6 & Ykp6z6);
assign Ykp6z6 = (Glp6z6 & Olp6z6);
assign Olp6z6 = (Wlp6z6 & Emp6z6);
assign Emp6z6 = (Mmp6z6 & Ump6z6);
assign Ump6z6 = (~(Cnp6z6 & G916z6));
assign G916z6 = (!M18nv6);
assign M18nv6 = (Xgl7z6[3] & A98nv6);
assign A98nv6 = (!Jv8nv6);
assign Cnp6z6 = (O916z6 ^ Knp6z6);
assign Knp6z6 = (!U24nv6);
assign O916z6 = (!Jkl7z6[28]);
assign Mmp6z6 = (~(Snp6z6 & Jv8nv6));
assign Jv8nv6 = (~(Og8nv6 & Aop6z6));
assign Aop6z6 = (~(Map6z6 & Igp6z6));
assign Snp6z6 = (Ea16z6 ^ Iop6z6);
assign Iop6z6 = (!U94nv6);
assign Ea16z6 = (!Jkl7z6[27]);
assign Wlp6z6 = (Qop6z6 & Yop6z6);
assign Yop6z6 = (~(Gpp6z6 & Q29nv6));
assign Q29nv6 = (!Og8nv6);
assign Og8nv6 = (A28nv6 & Opp6z6);
assign Opp6z6 = (!Mep6z6);
assign A28nv6 = (!Q38nv6);
assign Gpp6z6 = (Kb16z6 ^ Ng4nv6);
assign Kb16z6 = (!Jkl7z6[26]);
assign Qop6z6 = (~(Wpp6z6 & Q38nv6));
assign Q38nv6 = (~(O98nv6 & Eqp6z6));
assign Eqp6z6 = (~(Mep6z6 & Igp6z6));
assign Wpp6z6 = (Ac16z6 ^ B34nv6);
assign Ac16z6 = (!Jkl7z6[25]);
assign Glp6z6 = (Mqp6z6 & Uqp6z6);
assign Uqp6z6 = (~(Crp6z6 & Co8nv6));
assign Crp6z6 = (Gd16z6 ^ Krp6z6);
assign Krp6z6 = (!Y44nv6);
assign Gd16z6 = (!Jkl7z6[22]);
assign Mqp6z6 = (Srp6z6 & Asp6z6);
assign Asp6z6 = (~(Isp6z6 & Eb8nv6));
assign Eb8nv6 = (!O98nv6);
assign O98nv6 = (Ch8nv6 & Qsp6z6);
assign Isp6z6 = (Me16z6 ^ Ysp6z6);
assign Me16z6 = (!Jkl7z6[24]);
assign Srp6z6 = (~(Gtp6z6 & Si8nv6));
assign Si8nv6 = (!Ch8nv6);
assign Ch8nv6 = (~(Co8nv6 | Otp6z6));
assign Co8nv6 = (~(Xa8nv6 & Wtp6z6));
assign Wtp6z6 = (~(K3p6z6 & S3p6z6));
assign Xa8nv6 = (!Mt8nv6);
assign Gtp6z6 = (Cf16z6 ^ Gg4nv6);
assign Cf16z6 = (!Jkl7z6[23]);
assign Qkp6z6 = (Eup6z6 & Mup6z6);
assign Mup6z6 = (Uup6z6 & Cvp6z6);
assign Cvp6z6 = (Kvp6z6 & Svp6z6);
assign Svp6z6 = (~(Awp6z6 & Mt8nv6));
assign Mt8nv6 = (~(Li8nv6 & Iwp6z6));
assign Iwp6z6 = (~(Otp6z6 & K3p6z6));
assign Li8nv6 = (!M09nv6);
assign Awp6z6 = (Oh16z6 ^ Kb4nv6);
assign Oh16z6 = (!Jkl7z6[21]);
assign Kvp6z6 = (~(Qwp6z6 & M09nv6));
assign M09nv6 = (~(X38nv6 & Ywp6z6));
assign Ywp6z6 = (~(Map6z6 & S3p6z6));
assign X38nv6 = (!W68nv6);
assign Qwp6z6 = (Ei16z6 ^ Ri4nv6);
assign Ei16z6 = (!Jkl7z6[20]);
assign Uup6z6 = (Gxp6z6 & Oxp6z6);
assign Oxp6z6 = (~(Wxp6z6 & W68nv6));
assign W68nv6 = (~(Lb8nv6 & Eyp6z6));
assign Eyp6z6 = (~(Otp6z6 & Map6z6));
assign Lb8nv6 = (!Ke8nv6);
assign Wxp6z6 = (Sj16z6 ^ Myp6z6);
assign Myp6z6 = (!R44nv6);
assign Sj16z6 = (!Jkl7z6[19]);
assign Gxp6z6 = (~(Uyp6z6 & Ke8nv6));
assign Ke8nv6 = (~(Zi8nv6 & Czp6z6));
assign Czp6z6 = (~(Mep6z6 & S3p6z6));
assign Zi8nv6 = (!Yl8nv6);
assign Uyp6z6 = (Qk16z6 ^ Kzp6z6);
assign Kzp6z6 = (!Rb4nv6);
assign Qk16z6 = (!Jkl7z6[18]);
assign Eup6z6 = (Szp6z6 & Gl16z6);
assign Szp6z6 = (A0q6z6 & I0q6z6);
assign I0q6z6 = (~(Q0q6z6 & Yl8nv6));
assign Yl8nv6 = (~(P68nv6 & Y0q6z6));
assign Y0q6z6 = (~(Otp6z6 & Mep6z6));
assign Mep6z6 = (K3p6z6 & Map6z6);
assign K3p6z6 = (!Akp6z6);
assign Akp6z6 = (Xgl7z6[2] & Gl16z6);
assign Otp6z6 = (Igp6z6 & S3p6z6);
assign S3p6z6 = (!Qsp6z6);
assign Qsp6z6 = (Xgl7z6[4] & Gl16z6);
assign Igp6z6 = (!Kjp6z6);
assign Kjp6z6 = (Xgl7z6[1] & Gl16z6);
assign Q0q6z6 = (Um16z6 ^ Ki4nv6);
assign Um16z6 = (!Jkl7z6[17]);
assign A0q6z6 = (~(G1q6z6 & Jo8nv6));
assign Jo8nv6 = (!P68nv6);
assign P68nv6 = (Xgl7z6[5] & Gl16z6);
assign Gl16z6 = (O1q6z6 & Xgl7z6[0]);
assign O1q6z6 = (Sjy5z6 & W1q6z6);
assign W1q6z6 = (~(Dd9nv6 & Map6z6));
assign Map6z6 = (!Xgl7z6[3]);
assign Dd9nv6 = (E2q6z6 & M2q6z6);
assign M2q6z6 = (!Xgl7z6[5]);
assign E2q6z6 = (!Xgl7z6[4]);
assign G1q6z6 = (Kn16z6 ^ J74nv6);
assign Kn16z6 = (!Jkl7z6[16]);
assign Uyo6z6 = (~(W9n6z6 & U2q6z6));
assign U2q6z6 = (Man6z6 ? K3q6z6 : C3q6z6);
assign Man6z6 = (~(S3q6z6 & A4q6z6));
assign A4q6z6 = (I4q6z6 & Q4q6z6);
assign Q4q6z6 = (Y4q6z6 & G5q6z6);
assign G5q6z6 = (O5q6z6 & W5q6z6);
assign W5q6z6 = (~(Celet6 | E6q6z6));
assign E6q6z6 = (M6q6z6 & Lr6nv6);
assign Lr6nv6 = (!Df7nv6);
assign M6q6z6 = (Pa4nv6 ^ Ag87z6);
assign O5q6z6 = (U6q6z6 & C7q6z6);
assign C7q6z6 = (~(K7q6z6 & Q426z6));
assign Q426z6 = (!Qj6nv6);
assign K7q6z6 = (U24nv6 ^ V2diw6);
assign V2diw6 = (!Kf87z6);
assign U6q6z6 = (~(S7q6z6 & Bl7nv6));
assign Bl7nv6 = (!Sy6nv6);
assign S7q6z6 = (Ng4nv6 ^ Ue87z6);
assign Y4q6z6 = (A8q6z6 & I8q6z6);
assign I8q6z6 = (Q8q6z6 & Y8q6z6);
assign Y8q6z6 = (~(G9q6z6 & Ul6nv6));
assign G9q6z6 = (B34nv6 ^ Me87z6);
assign Q8q6z6 = (~(O9q6z6 & It6nv6));
assign It6nv6 = (!Sr6nv6);
assign O9q6z6 = (I826z6 ^ Ysp6z6);
assign I826z6 = (!Rul7z6[24]);
assign A8q6z6 = (W9q6z6 & Eaq6z6);
assign Eaq6z6 = (~(Maq6z6 & Qb7nv6));
assign Maq6z6 = (Kb4nv6 ^ Od87z6);
assign W9q6z6 = (~(Uaq6z6 & Ap6nv6));
assign Uaq6z6 = (R44nv6 ^ Nkciw6);
assign Nkciw6 = (!Qc87z6);
assign I4q6z6 = (Cbq6z6 & Kbq6z6);
assign Kbq6z6 = (Sbq6z6 & Acq6z6);
assign Acq6z6 = (Icq6z6 & Qcq6z6);
assign Qcq6z6 = (~(Ycq6z6 & Ow6nv6));
assign Ycq6z6 = (Rb4nv6 ^ Xiciw6);
assign Xiciw6 = (!Yc87z6);
assign Icq6z6 = (~(Gdq6z6 & C47nv6));
assign Gdq6z6 = (Ki4nv6 ^ Gd87z6);
assign Sbq6z6 = (Odq6z6 & Wdq6z6);
assign Wdq6z6 = (~(Eeq6z6 & Ah7nv6));
assign Eeq6z6 = (Jl4nv6 ^ Vaciw6);
assign Vaciw6 = (!Sb87z6);
assign Odq6z6 = (~(Meq6z6 & Fv6nv6));
assign Meq6z6 = (Ce4nv6 ^ I7ciw6);
assign I7ciw6 = (!Ea87z6);
assign Cbq6z6 = (Ueq6z6 & Cfq6z6);
assign Cfq6z6 = (~(Kfq6z6 & Mv6nv6));
assign Kfq6z6 = (Kv5nv6 ^ Apbiw6);
assign Apbiw6 = (!W987z6);
assign Ueq6z6 = (Sfq6z6 & Agq6z6);
assign Agq6z6 = (~(Igq6z6 & P77nv6));
assign Igq6z6 = (H64nv6 ^ P0ciw6);
assign P0ciw6 = (!Ua87z6);
assign Sfq6z6 = (~(M27nv6 & Qgq6z6));
assign Qgq6z6 = (Kz16z6 ^ Ghp6z6);
assign Kz16z6 = (!Rul7z6[8]);
assign S3q6z6 = (Ygq6z6 & Ghq6z6);
assign Ghq6z6 = (Ohq6z6 & Whq6z6);
assign Whq6z6 = (Eiq6z6 & Miq6z6);
assign Miq6z6 = (Uiq6z6 & Cjq6z6);
assign Cjq6z6 = (~(Kjq6z6 & Nd7nv6));
assign Kjq6z6 = (U94nv6 ^ Y0diw6);
assign Y0diw6 = (!Cf87z6);
assign Uiq6z6 = (~(Sjq6z6 & Zy6nv6));
assign Sjq6z6 = (S4diw6 ^ Ico6z6);
assign S4diw6 = (!Sf87z6);
assign Eiq6z6 = (Akq6z6 & Ikq6z6);
assign Ikq6z6 = (~(Qkq6z6 & Ej7nv6));
assign Qkq6z6 = (Ri4nv6 ^ Ic87z6);
assign Akq6z6 = (~(Ykq6z6 & G67nv6));
assign Ykq6z6 = (Y44nv6 ^ Eqciw6);
assign Eqciw6 = (!Wd87z6);
assign Ohq6z6 = (Glq6z6 & Olq6z6);
assign Olq6z6 = (~(Wlq6z6 & Xb7nv6));
assign Xb7nv6 = (Ah7nv6 | Emq6z6);
assign Ah7nv6 = (~(Hp6nv6 & Mmq6z6));
assign Mmq6z6 = (~(Umq6z6 & N67nv6));
assign Hp6nv6 = (!Rn6nv6);
assign Wlq6z6 = (Je4nv6 ^ Zcciw6);
assign Zcciw6 = (!Ac87z6);
assign Glq6z6 = (Cnq6z6 & Knq6z6);
assign Knq6z6 = (~(Snq6z6 & W07nv6));
assign W07nv6 = (!Gz6nv6);
assign Snq6z6 = (Gg4nv6 ^ Ol77z6);
assign Cnq6z6 = (~(Aoq6z6 & Rn6nv6));
assign Rn6nv6 = (~(Vw6nv6 & Ioq6z6));
assign Ioq6z6 = (~(Emq6z6 & Umq6z6));
assign Vw6nv6 = (!Fv6nv6);
assign Fv6nv6 = (~(J47nv6 & Qoq6z6));
assign Qoq6z6 = (~(Yoq6z6 & N67nv6));
assign J47nv6 = (!A37nv6);
assign Aoq6z6 = (Q74nv6 ^ F9ciw6);
assign F9ciw6 = (!Kb87z6);
assign Ygq6z6 = (Gpq6z6 & Opq6z6);
assign Opq6z6 = (Wpq6z6 & Eqq6z6);
assign Eqq6z6 = (Mqq6z6 & Uqq6z6);
assign Uqq6z6 = (~(Crq6z6 & Uy16z6));
assign Crq6z6 = (Hd4nv6 ^ Zybiw6);
assign Zybiw6 = (!Cb87z6);
assign Mqq6z6 = (~(Krq6z6 & T27nv6));
assign T27nv6 = (Srq6z6 & Emq6z6);
assign Srq6z6 = (Asq6z6 & Umq6z6);
assign Krq6z6 = (Ak4nv6 ^ Uq16z6);
assign Uq16z6 = (!Rul7z6[5]);
assign Wpq6z6 = (Isq6z6 & Qsq6z6);
assign Qsq6z6 = (~(Ysq6z6 & Yn6nv6));
assign Yn6nv6 = (Gtq6z6 | Mv6nv6);
assign Mv6nv6 = (M27nv6 & Umq6z6);
assign Gtq6z6 = (Emq6z6 & Asq6z6);
assign Ysq6z6 = (Tp5nv6 ^ Gsbiw6);
assign Gsbiw6 = (!O987z6);
assign Isq6z6 = (~(Otq6z6 & A37nv6));
assign A37nv6 = (~(Kn6nv6 & Wtq6z6));
assign Wtq6z6 = (~(Emq6z6 & Yoq6z6));
assign Kn6nv6 = (!P77nv6);
assign P77nv6 = (~(Yu6nv6 & Euq6z6));
assign Euq6z6 = (~(Muq6z6 & N67nv6));
assign Yu6nv6 = (!Uy16z6);
assign Uy16z6 = (~(Uuq6z6 & Ji7nv6));
assign Ji7nv6 = (!M27nv6);
assign M27nv6 = (N67nv6 & Asq6z6);
assign Uuq6z6 = (~(Emq6z6 & Muq6z6));
assign Emq6z6 = (N67nv6 & Cvq6z6);
assign Otq6z6 = (Cl4nv6 ^ V3ciw6);
assign V3ciw6 = (!Ma87z6);
assign Gpq6z6 = (Kvq6z6 & Yc26z6);
assign Kvq6z6 = (Svq6z6 & Awq6z6);
assign Awq6z6 = (~(Iwq6z6 & Xj6nv6));
assign Xj6nv6 = (!T97nv6);
assign T97nv6 = (Df7nv6 & Qwq6z6);
assign Df7nv6 = (Uk7nv6 & Ywq6z6);
assign Uk7nv6 = (!Zy6nv6);
assign Zy6nv6 = (~(Qj6nv6 & Gxq6z6));
assign Gxq6z6 = (~(Umq6z6 & Cvq6z6));
assign Qj6nv6 = (Frl7z6[3] & Er6nv6);
assign Er6nv6 = (!Nd7nv6);
assign Nd7nv6 = (~(Sy6nv6 & Oxq6z6));
assign Oxq6z6 = (~(Yoq6z6 & Cvq6z6));
assign Sy6nv6 = (Ek6nv6 & Wxq6z6);
assign Wxq6z6 = (!Muq6z6);
assign Ek6nv6 = (!Ul6nv6);
assign Ul6nv6 = (~(Sr6nv6 & Eyq6z6));
assign Eyq6z6 = (~(Muq6z6 & Cvq6z6));
assign Sr6nv6 = (Gz6nv6 & Myq6z6);
assign Gz6nv6 = (~(G67nv6 | Uyq6z6));
assign G67nv6 = (~(Bt6nv6 & Czq6z6));
assign Czq6z6 = (~(Umq6z6 & Asq6z6));
assign Bt6nv6 = (!Qb7nv6);
assign Qb7nv6 = (~(P07nv6 & Kzq6z6));
assign Kzq6z6 = (~(Uyq6z6 & Umq6z6));
assign P07nv6 = (!Ej7nv6);
assign Ej7nv6 = (~(Bm6nv6 & Szq6z6));
assign Szq6z6 = (~(Yoq6z6 & Asq6z6));
assign Bm6nv6 = (!Ap6nv6);
assign Ap6nv6 = (~(Pt6nv6 & A0r6z6));
assign A0r6z6 = (~(Uyq6z6 & Yoq6z6));
assign Pt6nv6 = (!Ow6nv6);
assign Ow6nv6 = (~(D17nv6 & I0r6z6));
assign I0r6z6 = (~(Muq6z6 & Asq6z6));
assign D17nv6 = (!C47nv6);
assign C47nv6 = (~(To6nv6 & Q0r6z6));
assign Q0r6z6 = (~(Uyq6z6 & Muq6z6));
assign Muq6z6 = (Umq6z6 & Yoq6z6);
assign Umq6z6 = (!Ywq6z6);
assign Ywq6z6 = (Frl7z6[2] & Yc26z6);
assign Uyq6z6 = (Cvq6z6 & Asq6z6);
assign Asq6z6 = (!Myq6z6);
assign Myq6z6 = (Frl7z6[4] & Yc26z6);
assign Cvq6z6 = (!Qwq6z6);
assign Qwq6z6 = (Frl7z6[1] & Yc26z6);
assign Iwq6z6 = (W34nv6 ^ Ee87z6);
assign Svq6z6 = (~(Y0r6z6 & N67nv6));
assign N67nv6 = (!To6nv6);
assign To6nv6 = (Frl7z6[5] & Yc26z6);
assign Yc26z6 = (G1r6z6 & Frl7z6[0]);
assign G1r6z6 = (Sjy5z6 & O1r6z6);
assign O1r6z6 = (~(Ov7nv6 & Yoq6z6));
assign Yoq6z6 = (!Frl7z6[3]);
assign Ov7nv6 = (W1r6z6 & E2r6z6);
assign E2r6z6 = (!Frl7z6[5]);
assign W1r6z6 = (!Frl7z6[4]);
assign Y0r6z6 = (Me26z6 ^ J74nv6);
assign Me26z6 = (!Rul7z6[16]);
assign K3q6z6 = (M2r6z6 | U2r6z6);
assign U2r6z6 = (C3r6z6 & Xgl7z6[22]);
assign C3r6z6 = (Ysn6z6 & K3r6z6);
assign K3r6z6 = (Xgl7z6[20] | Xgl7z6[21]);
assign M2r6z6 = (Xgl7z6[20] ? A4r6z6 : S3r6z6);
assign A4r6z6 = (~(Glm6z6 | Xgl7z6[21]));
assign S3r6z6 = (!I4r6z6);
assign I4r6z6 = (Xgl7z6[21] ? Wtn6z6 : Xgl7z6[22]);
assign C3q6z6 = (Q4r6z6 | Y4r6z6);
assign Y4r6z6 = (G5r6z6 & Frl7z6[22]);
assign G5r6z6 = (Ysn6z6 & O5r6z6);
assign O5r6z6 = (Frl7z6[20] | Frl7z6[21]);
assign Q4r6z6 = (Frl7z6[20] ? E6r6z6 : W5r6z6);
assign E6r6z6 = (~(Glm6z6 | Frl7z6[21]));
assign W5r6z6 = (!M6r6z6);
assign M6r6z6 = (Frl7z6[21] ? Wtn6z6 : Frl7z6[22]);
assign W9n6z6 = (~(U6r6z6 | Aga6z6));
assign Myo6z6 = (~(Kvo6z6 & C7r6z6));
assign C7r6z6 = (Qcn6z6 ? S7r6z6 : K7r6z6);
assign Qcn6z6 = (A8r6z6 & I8r6z6);
assign I8r6z6 = (Q8r6z6 & Y8r6z6);
assign Y8r6z6 = (G9r6z6 & O9r6z6);
assign O9r6z6 = (W9r6z6 & Ear6z6);
assign Ear6z6 = (~(Caiet6 | Mar6z6));
assign Mar6z6 = (Uar6z6 & Mpcnv6);
assign Mpcnv6 = (!Eddnv6);
assign Uar6z6 = (Pa4nv6 ^ Um87z6);
assign W9r6z6 = (Cbr6z6 & Kbr6z6);
assign Kbr6z6 = (~(Sbr6z6 & Sv26z6));
assign Sv26z6 = (!Rhcnv6);
assign Sbr6z6 = (U24nv6 ^ A2diw6);
assign A2diw6 = (!Em87z6);
assign Cbr6z6 = (~(Acr6z6 & Vidnv6));
assign Vidnv6 = (!Twcnv6);
assign Acr6z6 = (Ng4nv6 ^ Ol87z6);
assign G9r6z6 = (Icr6z6 & Qcr6z6);
assign Qcr6z6 = (Ycr6z6 & Gdr6z6);
assign Gdr6z6 = (~(Odr6z6 & Vjcnv6));
assign Odr6z6 = (B34nv6 ^ Gl87z6);
assign Ycr6z6 = (~(Wdr6z6 & Jrcnv6));
assign Jrcnv6 = (!Tpcnv6);
assign Wdr6z6 = (Kz26z6 ^ Ysp6z6);
assign Kz26z6 = (!Lpk7z6[24]);
assign Icr6z6 = (Eer6z6 & Mer6z6);
assign Mer6z6 = (~(Uer6z6 & R9dnv6));
assign Uer6z6 = (Kb4nv6 ^ Ik87z6);
assign Eer6z6 = (~(Cfr6z6 & Bncnv6));
assign Cfr6z6 = (R44nv6 ^ Sjciw6);
assign Sjciw6 = (!Kj87z6);
assign Q8r6z6 = (Kfr6z6 & Sfr6z6);
assign Sfr6z6 = (Agr6z6 & Igr6z6);
assign Igr6z6 = (Qgr6z6 & Ygr6z6);
assign Ygr6z6 = (~(Ghr6z6 & Pucnv6));
assign Ghr6z6 = (Rb4nv6 ^ Ciciw6);
assign Ciciw6 = (!Sj87z6);
assign Qgr6z6 = (~(Ohr6z6 & D2dnv6));
assign Ohr6z6 = (Ki4nv6 ^ Ak87z6);
assign Agr6z6 = (Whr6z6 & Eir6z6);
assign Eir6z6 = (~(Mir6z6 & Bfdnv6));
assign Mir6z6 = (Jl4nv6 ^ Aaciw6);
assign Aaciw6 = (!Mi87z6);
assign Whr6z6 = (~(Uir6z6 & Gtcnv6));
assign Uir6z6 = (Ce4nv6 ^ L5ciw6);
assign L5ciw6 = (!Yg87z6);
assign Kfr6z6 = (Cjr6z6 & Kjr6z6);
assign Kjr6z6 = (~(Sjr6z6 & Ntcnv6));
assign Sjr6z6 = (Kv5nv6 ^ Fobiw6);
assign Fobiw6 = (!Qg87z6);
assign Cjr6z6 = (Akr6z6 & Ikr6z6);
assign Ikr6z6 = (~(Qkr6z6 & Q5dnv6));
assign Qkr6z6 = (H64nv6 ^ Uzbiw6);
assign Uzbiw6 = (!Oh87z6);
assign Akr6z6 = (~(N0dnv6 & Ykr6z6));
assign Ykr6z6 = (Mq26z6 ^ Ghp6z6);
assign Mq26z6 = (!Lpk7z6[8]);
assign A8r6z6 = (Glr6z6 & Olr6z6);
assign Olr6z6 = (Wlr6z6 & Emr6z6);
assign Emr6z6 = (Mmr6z6 & Umr6z6);
assign Umr6z6 = (Cnr6z6 & Knr6z6);
assign Knr6z6 = (~(Snr6z6 & Obdnv6));
assign Snr6z6 = (U94nv6 ^ D0diw6);
assign D0diw6 = (!Wl87z6);
assign Cnr6z6 = (~(Aor6z6 & Axcnv6));
assign Aor6z6 = (X3diw6 ^ Ico6z6);
assign X3diw6 = (!Mm87z6);
assign Mmr6z6 = (Ior6z6 & Qor6z6);
assign Qor6z6 = (~(Yor6z6 & Rgdnv6));
assign Yor6z6 = (Ri4nv6 ^ Cj87z6);
assign Ior6z6 = (~(Gpr6z6 & H4dnv6));
assign Gpr6z6 = (Y44nv6 ^ Jpciw6);
assign Jpciw6 = (!Qk87z6);
assign Wlr6z6 = (Opr6z6 & Wpr6z6);
assign Wpr6z6 = (~(Eqr6z6 & Y9dnv6));
assign Y9dnv6 = (Bfdnv6 | Mqr6z6);
assign Bfdnv6 = (~(Incnv6 & Uqr6z6));
assign Uqr6z6 = (~(Crr6z6 & O4dnv6));
assign Incnv6 = (!Slcnv6);
assign Eqr6z6 = (Je4nv6 ^ Xbciw6);
assign Xbciw6 = (!Ui87z6);
assign Opr6z6 = (Krr6z6 & Srr6z6);
assign Srr6z6 = (~(Asr6z6 & Xycnv6));
assign Xycnv6 = (!Hxcnv6);
assign Asr6z6 = (Gg4nv6 ^ Mm77z6);
assign Krr6z6 = (~(Isr6z6 & Slcnv6));
assign Slcnv6 = (~(Wucnv6 & Qsr6z6));
assign Qsr6z6 = (~(Mqr6z6 & Crr6z6));
assign Wucnv6 = (!Gtcnv6);
assign Gtcnv6 = (~(K2dnv6 & Ysr6z6));
assign Ysr6z6 = (~(Gtr6z6 & O4dnv6));
assign K2dnv6 = (!B1dnv6);
assign Isr6z6 = (Q74nv6 ^ K8ciw6);
assign K8ciw6 = (!Ei87z6);
assign Glr6z6 = (Otr6z6 & Wtr6z6);
assign Wtr6z6 = (Eur6z6 & Mur6z6);
assign Mur6z6 = (Uur6z6 & Cvr6z6);
assign Cvr6z6 = (~(Kvr6z6 & Wp26z6));
assign Kvr6z6 = (Hd4nv6 ^ Eybiw6);
assign Eybiw6 = (!Wh87z6);
assign Uur6z6 = (~(Svr6z6 & U0dnv6));
assign U0dnv6 = (Awr6z6 & Mqr6z6);
assign Awr6z6 = (Iwr6z6 & Crr6z6);
assign Svr6z6 = (Ak4nv6 ^ Wh26z6);
assign Wh26z6 = (!Lpk7z6[5]);
assign Eur6z6 = (Qwr6z6 & Ywr6z6);
assign Ywr6z6 = (~(Gxr6z6 & Zlcnv6));
assign Zlcnv6 = (Oxr6z6 | Ntcnv6);
assign Ntcnv6 = (N0dnv6 & Crr6z6);
assign Oxr6z6 = (Mqr6z6 & Iwr6z6);
assign Gxr6z6 = (Tp5nv6 ^ Jqbiw6);
assign Jqbiw6 = (!Ig87z6);
assign Qwr6z6 = (~(Wxr6z6 & B1dnv6));
assign B1dnv6 = (~(Llcnv6 & Eyr6z6));
assign Eyr6z6 = (~(Mqr6z6 & Gtr6z6));
assign Llcnv6 = (!Q5dnv6);
assign Q5dnv6 = (~(Zscnv6 & Myr6z6));
assign Myr6z6 = (~(Uyr6z6 & O4dnv6));
assign Zscnv6 = (!Wp26z6);
assign Wp26z6 = (~(Czr6z6 & Aidnv6));
assign Aidnv6 = (!N0dnv6);
assign N0dnv6 = (O4dnv6 & Iwr6z6);
assign Czr6z6 = (~(Mqr6z6 & Uyr6z6));
assign Mqr6z6 = (O4dnv6 & Kzr6z6);
assign Wxr6z6 = (Cl4nv6 ^ Y1ciw6);
assign Y1ciw6 = (!Gh87z6);
assign Otr6z6 = (Szr6z6 & A436z6);
assign Szr6z6 = (A0s6z6 & I0s6z6);
assign I0s6z6 = (~(Q0s6z6 & Yhcnv6));
assign Yhcnv6 = (!U7dnv6);
assign U7dnv6 = (Eddnv6 & Y0s6z6);
assign Eddnv6 = (Oidnv6 & G1s6z6);
assign Oidnv6 = (!Axcnv6);
assign Axcnv6 = (~(Rhcnv6 & O1s6z6));
assign O1s6z6 = (~(Crr6z6 & Kzr6z6));
assign Rhcnv6 = (Zlk7z6[3] & Fpcnv6);
assign Fpcnv6 = (!Obdnv6);
assign Obdnv6 = (~(Twcnv6 & W1s6z6));
assign W1s6z6 = (~(Gtr6z6 & Kzr6z6));
assign Twcnv6 = (Ficnv6 & E2s6z6);
assign E2s6z6 = (!Uyr6z6);
assign Ficnv6 = (!Vjcnv6);
assign Vjcnv6 = (~(Tpcnv6 & M2s6z6));
assign M2s6z6 = (~(Uyr6z6 & Kzr6z6));
assign Tpcnv6 = (Hxcnv6 & U2s6z6);
assign Hxcnv6 = (~(H4dnv6 | C3s6z6));
assign H4dnv6 = (~(Crcnv6 & K3s6z6));
assign K3s6z6 = (~(Crr6z6 & Iwr6z6));
assign Crcnv6 = (!R9dnv6);
assign R9dnv6 = (~(Qycnv6 & S3s6z6));
assign S3s6z6 = (~(C3s6z6 & Crr6z6));
assign Qycnv6 = (!Rgdnv6);
assign Rgdnv6 = (~(Ckcnv6 & A4s6z6));
assign A4s6z6 = (~(Gtr6z6 & Iwr6z6));
assign Ckcnv6 = (!Bncnv6);
assign Bncnv6 = (~(Qrcnv6 & I4s6z6));
assign I4s6z6 = (~(C3s6z6 & Gtr6z6));
assign Qrcnv6 = (!Pucnv6);
assign Pucnv6 = (~(Ezcnv6 & Q4s6z6));
assign Q4s6z6 = (~(Uyr6z6 & Iwr6z6));
assign Ezcnv6 = (!D2dnv6);
assign D2dnv6 = (~(Umcnv6 & Y4s6z6));
assign Y4s6z6 = (~(C3s6z6 & Uyr6z6));
assign Uyr6z6 = (Crr6z6 & Gtr6z6);
assign Crr6z6 = (!G1s6z6);
assign G1s6z6 = (Zlk7z6[2] & A436z6);
assign C3s6z6 = (Kzr6z6 & Iwr6z6);
assign Iwr6z6 = (!U2s6z6);
assign U2s6z6 = (Zlk7z6[4] & A436z6);
assign Kzr6z6 = (!Y0s6z6);
assign Y0s6z6 = (Zlk7z6[1] & A436z6);
assign Q0s6z6 = (W34nv6 ^ Yk87z6);
assign A0s6z6 = (~(G5s6z6 & O4dnv6));
assign O4dnv6 = (!Umcnv6);
assign Umcnv6 = (Zlk7z6[5] & A436z6);
assign A436z6 = (O5s6z6 & Zlk7z6[0]);
assign O5s6z6 = (Sjy5z6 & W5s6z6);
assign W5s6z6 = (~(Itdnv6 & Gtr6z6));
assign Gtr6z6 = (!Zlk7z6[3]);
assign Itdnv6 = (E6s6z6 & M6s6z6);
assign M6s6z6 = (!Zlk7z6[5]);
assign E6s6z6 = (!Zlk7z6[4]);
assign G5s6z6 = (O536z6 ^ J74nv6);
assign O536z6 = (!Lpk7z6[16]);
assign S7r6z6 = (U6s6z6 | C7s6z6);
assign C7s6z6 = (K7s6z6 & Zlk7z6[22]);
assign K7s6z6 = (Ysn6z6 & S7s6z6);
assign S7s6z6 = (Zlk7z6[20] | Zlk7z6[21]);
assign U6s6z6 = (Zlk7z6[20] ? I8s6z6 : A8s6z6);
assign I8s6z6 = (~(Glm6z6 | Zlk7z6[21]));
assign A8s6z6 = (!Q8s6z6);
assign Q8s6z6 = (Zlk7z6[21] ? Wtn6z6 : Zlk7z6[22]);
assign K7r6z6 = (Y8s6z6 | G9s6z6);
assign G9s6z6 = (O9s6z6 & Rbk7z6[22]);
assign O9s6z6 = (Ysn6z6 & W9s6z6);
assign W9s6z6 = (Rbk7z6[20] | Rbk7z6[21]);
assign Y8s6z6 = (Rbk7z6[20] ? Mas6z6 : Eas6z6);
assign Mas6z6 = (~(Glm6z6 | Rbk7z6[21]));
assign Eas6z6 = (!Uas6z6);
assign Uas6z6 = (Rbk7z6[21] ? Wtn6z6 : Rbk7z6[22]);
assign Kvo6z6 = (~(Cvn6z6 | Cbs6z6));
assign Cbs6z6 = (Kbs6z6 & Sbs6z6);
assign Sbs6z6 = (Acs6z6 & Ics6z6);
assign Ics6z6 = (Qcs6z6 & Ycs6z6);
assign Ycs6z6 = (Gds6z6 & Ods6z6);
assign Ods6z6 = (~(C2jet6 | Wds6z6));
assign Wds6z6 = (Ees6z6 & Mjbnv6);
assign Mjbnv6 = (Mes6z6 & Ues6z6);
assign Mes6z6 = (Cfs6z6 & Kfs6z6);
assign Ees6z6 = (Ak4nv6 ^ Kz36z6);
assign Kz36z6 = (!Tzk7z6[5]);
assign Gds6z6 = (Sfs6z6 & Ags6z6);
assign Ags6z6 = (~(Igs6z6 & R4bnv6));
assign R4bnv6 = (Qgs6z6 | Fcbnv6);
assign Qgs6z6 = (Ues6z6 & Kfs6z6);
assign Igs6z6 = (Tp5nv6 ^ Xqbiw6);
assign Xqbiw6 = (!Cn87z6);
assign Sfs6z6 = (~(Ygs6z6 & Fcbnv6));
assign Fcbnv6 = (Fjbnv6 & Cfs6z6);
assign Ygs6z6 = (Kv5nv6 ^ Mobiw6);
assign Mobiw6 = (!Kn87z6);
assign Qcs6z6 = (Ghs6z6 & Ohs6z6);
assign Ohs6z6 = (Whs6z6 & Eis6z6);
assign Eis6z6 = (~(Mis6z6 & Qsbnv6));
assign Qsbnv6 = (Txbnv6 | Ues6z6);
assign Mis6z6 = (Je4nv6 ^ Ecciw6);
assign Ecciw6 = (!Op87z6);
assign Whs6z6 = (~(Uis6z6 & Txbnv6));
assign Txbnv6 = (~(A6bnv6 & Cjs6z6));
assign Cjs6z6 = (~(Cfs6z6 & Gnbnv6));
assign A6bnv6 = (!K4bnv6);
assign Uis6z6 = (Jl4nv6 ^ Haciw6);
assign Haciw6 = (!Gp87z6);
assign Ghs6z6 = (Kjs6z6 & Sjs6z6);
assign Sjs6z6 = (~(Aks6z6 & K4bnv6));
assign K4bnv6 = (~(Odbnv6 & Iks6z6));
assign Iks6z6 = (~(Ues6z6 & Cfs6z6));
assign Odbnv6 = (!Ybbnv6);
assign Aks6z6 = (Q74nv6 ^ R8ciw6);
assign R8ciw6 = (!Yo87z6);
assign Kjs6z6 = (~(Qks6z6 & Ybbnv6));
assign Ybbnv6 = (~(Clbnv6 & Yks6z6));
assign Yks6z6 = (~(Gls6z6 & Gnbnv6));
assign Clbnv6 = (!Tjbnv6);
assign Qks6z6 = (Ce4nv6 ^ Z5ciw6);
assign Z5ciw6 = (!Sn87z6);
assign Acs6z6 = (Ols6z6 & Wls6z6);
assign Wls6z6 = (Ems6z6 & Mms6z6);
assign Mms6z6 = (Ums6z6 & Cns6z6);
assign Cns6z6 = (~(Kns6z6 & Tjbnv6));
assign Tjbnv6 = (~(D4bnv6 & Sns6z6));
assign Sns6z6 = (~(Ues6z6 & Gls6z6));
assign D4bnv6 = (!Iobnv6);
assign Kns6z6 = (Cl4nv6 ^ M2ciw6);
assign M2ciw6 = (!Ao87z6);
assign Ums6z6 = (~(Aos6z6 & Iobnv6));
assign Iobnv6 = (~(Rbbnv6 & Ios6z6));
assign Ios6z6 = (~(Qos6z6 & Gnbnv6));
assign Rbbnv6 = (!K746z6);
assign Aos6z6 = (H64nv6 ^ B0ciw6);
assign B0ciw6 = (!Io87z6);
assign Ems6z6 = (Yos6z6 & Gps6z6);
assign Gps6z6 = (~(Ops6z6 & K746z6));
assign K746z6 = (~(Wps6z6 & S0cnv6));
assign S0cnv6 = (!Fjbnv6);
assign Wps6z6 = (~(Qos6z6 & Ues6z6));
assign Ues6z6 = (Eqs6z6 & Gnbnv6);
assign Ops6z6 = (Hd4nv6 ^ Lybiw6);
assign Lybiw6 = (!Qo87z6);
assign Yos6z6 = (~(Fjbnv6 & Mqs6z6));
assign Mqs6z6 = (A846z6 ^ Ghp6z6);
assign A846z6 = (!Tzk7z6[8]);
assign Fjbnv6 = (Kfs6z6 & Gnbnv6);
assign Ols6z6 = (Uqs6z6 & Crs6z6);
assign Crs6z6 = (~(Krs6z6 & Sfbnv6));
assign Krs6z6 = (E4diw6 ^ Ico6z6);
assign E4diw6 = (!Gt87z6);
assign Uqs6z6 = (Srs6z6 & Ass6z6);
assign Ass6z6 = (~(Iss6z6 & Q0bnv6));
assign Q0bnv6 = (!Mqbnv6);
assign Mqbnv6 = (Wvbnv6 & Qss6z6);
assign Iss6z6 = (W34nv6 ^ Sr87z6);
assign Srs6z6 = (~(Yss6z6 & E8bnv6));
assign E8bnv6 = (!Wvbnv6);
assign Wvbnv6 = (G1cnv6 & Gts6z6);
assign G1cnv6 = (!Sfbnv6);
assign Sfbnv6 = (~(J0bnv6 & Ots6z6));
assign Ots6z6 = (~(Cfs6z6 & Eqs6z6));
assign Yss6z6 = (Pa4nv6 ^ Ot87z6);
assign Kbs6z6 = (Wts6z6 & Eus6z6);
assign Eus6z6 = (Mus6z6 & Uus6z6);
assign Uus6z6 = (Cvs6z6 & Kvs6z6);
assign Kvs6z6 = (Svs6z6 & Aws6z6);
assign Aws6z6 = (~(Iws6z6 & Gd46z6));
assign Gd46z6 = (!J0bnv6);
assign J0bnv6 = (Hwk7z6[3] & X7bnv6);
assign X7bnv6 = (!Gubnv6);
assign Iws6z6 = (U24nv6 ^ H2diw6);
assign H2diw6 = (!Ys87z6);
assign Svs6z6 = (~(Qws6z6 & Gubnv6));
assign Gubnv6 = (~(Lfbnv6 & Yws6z6));
assign Yws6z6 = (~(Gls6z6 & Eqs6z6));
assign Qws6z6 = (U94nv6 ^ K0diw6);
assign K0diw6 = (!Qs87z6);
assign Cvs6z6 = (Gxs6z6 & Oxs6z6);
assign Oxs6z6 = (~(Wxs6z6 & N1cnv6));
assign N1cnv6 = (!Lfbnv6);
assign Lfbnv6 = (X0bnv6 & Eys6z6);
assign Eys6z6 = (!Qos6z6);
assign X0bnv6 = (!N2bnv6);
assign Wxs6z6 = (Ng4nv6 ^ Is87z6);
assign Gxs6z6 = (~(Mys6z6 & N2bnv6));
assign N2bnv6 = (~(L8bnv6 & Uys6z6));
assign Uys6z6 = (~(Qos6z6 & Eqs6z6));
assign Mys6z6 = (B34nv6 ^ As87z6);
assign Mus6z6 = (Czs6z6 & Kzs6z6);
assign Kzs6z6 = (~(Szs6z6 & Zmbnv6));
assign Szs6z6 = (Y44nv6 ^ Qpciw6);
assign Qpciw6 = (!Kr87z6);
assign Czs6z6 = (A0t6z6 & I0t6z6);
assign I0t6z6 = (~(Q0t6z6 & Babnv6));
assign Babnv6 = (!L8bnv6);
assign L8bnv6 = (Zfbnv6 & Y0t6z6);
assign Q0t6z6 = (Yg46z6 ^ Ysp6z6);
assign Yg46z6 = (!Tzk7z6[24]);
assign A0t6z6 = (~(G1t6z6 & Phbnv6));
assign Phbnv6 = (!Zfbnv6);
assign Zfbnv6 = (~(Zmbnv6 | O1t6z6));
assign Zmbnv6 = (~(U9bnv6 & W1t6z6));
assign W1t6z6 = (~(Cfs6z6 & Kfs6z6));
assign U9bnv6 = (!Jsbnv6);
assign G1t6z6 = (Gg4nv6 ^ Em77z6);
assign Wts6z6 = (E2t6z6 & M2t6z6);
assign M2t6z6 = (U2t6z6 & C3t6z6);
assign C3t6z6 = (K3t6z6 & S3t6z6);
assign S3t6z6 = (~(A4t6z6 & Jsbnv6));
assign Jsbnv6 = (~(Ihbnv6 & I4t6z6));
assign I4t6z6 = (~(O1t6z6 & Cfs6z6));
assign Ihbnv6 = (!Jzbnv6);
assign A4t6z6 = (Kb4nv6 ^ Cr87z6);
assign K3t6z6 = (~(Q4t6z6 & Jzbnv6));
assign Jzbnv6 = (~(U2bnv6 & Y4t6z6));
assign Y4t6z6 = (~(Gls6z6 & Kfs6z6));
assign U2bnv6 = (!T5bnv6);
assign Q4t6z6 = (Ri4nv6 ^ Wp87z6);
assign U2t6z6 = (G5t6z6 & O5t6z6);
assign O5t6z6 = (~(W5t6z6 & T5bnv6));
assign T5bnv6 = (~(Iabnv6 & E6t6z6));
assign E6t6z6 = (~(O1t6z6 & Gls6z6));
assign Iabnv6 = (!Hdbnv6);
assign W5t6z6 = (R44nv6 ^ Zjciw6);
assign Zjciw6 = (!Eq87z6);
assign G5t6z6 = (~(M6t6z6 & Hdbnv6));
assign Hdbnv6 = (~(Whbnv6 & U6t6z6));
assign U6t6z6 = (~(Qos6z6 & Kfs6z6));
assign Whbnv6 = (!Vkbnv6);
assign M6t6z6 = (Rb4nv6 ^ Jiciw6);
assign Jiciw6 = (!Mq87z6);
assign E2t6z6 = (C7t6z6 & Ol46z6);
assign C7t6z6 = (K7t6z6 & S7t6z6);
assign S7t6z6 = (~(A8t6z6 & Vkbnv6));
assign Vkbnv6 = (~(M5bnv6 & I8t6z6));
assign I8t6z6 = (~(O1t6z6 & Qos6z6));
assign Qos6z6 = (Cfs6z6 & Gls6z6);
assign Cfs6z6 = (!Gts6z6);
assign Gts6z6 = (Hwk7z6[2] & Ol46z6);
assign O1t6z6 = (Eqs6z6 & Kfs6z6);
assign Kfs6z6 = (!Y0t6z6);
assign Y0t6z6 = (Hwk7z6[4] & Ol46z6);
assign Eqs6z6 = (!Qss6z6);
assign Qss6z6 = (Hwk7z6[1] & Ol46z6);
assign A8t6z6 = (Ki4nv6 ^ Uq87z6);
assign K7t6z6 = (~(Q8t6z6 & Gnbnv6));
assign Gnbnv6 = (!M5bnv6);
assign M5bnv6 = (Hwk7z6[5] & Ol46z6);
assign Ol46z6 = (Y8t6z6 & Hwk7z6[0]);
assign Y8t6z6 = (Sjy5z6 & G9t6z6);
assign G9t6z6 = (~(Accnv6 & Gls6z6));
assign Gls6z6 = (!Hwk7z6[3]);
assign Accnv6 = (O9t6z6 & W9t6z6);
assign W9t6z6 = (!Hwk7z6[5]);
assign O9t6z6 = (!Hwk7z6[4]);
assign Q8t6z6 = (Cn46z6 ^ J74nv6);
assign Cn46z6 = (!Tzk7z6[16]);
assign Cvn6z6 = (Eat6z6 & Mat6z6);
assign Mat6z6 = (Uat6z6 & Cbt6z6);
assign Cbt6z6 = (Kbt6z6 & Sbt6z6);
assign Sbt6z6 = (Act6z6 & Ict6z6);
assign Ict6z6 = (~(Cujet6 | Qct6z6));
assign Qct6z6 = (Yct6z6 & Pq9nv6);
assign Pq9nv6 = (!Heanv6);
assign Yct6z6 = (Pa4nv6 ^ I097z6);
assign Act6z6 = (Gdt6z6 & Odt6z6);
assign Odt6z6 = (~(Wdt6z6 & Um36z6));
assign Um36z6 = (!Ui9nv6);
assign Wdt6z6 = (U24nv6 ^ O2diw6);
assign O2diw6 = (!Sz87z6);
assign Gdt6z6 = (~(Eet6z6 & Yjanv6));
assign Yjanv6 = (!Wx9nv6);
assign Eet6z6 = (Ng4nv6 ^ Cz87z6);
assign Kbt6z6 = (Met6z6 & Uet6z6);
assign Uet6z6 = (Cft6z6 & Kft6z6);
assign Kft6z6 = (~(Sft6z6 & Yk9nv6));
assign Sft6z6 = (B34nv6 ^ Uy87z6);
assign Cft6z6 = (~(Agt6z6 & Ms9nv6));
assign Ms9nv6 = (!Wq9nv6);
assign Agt6z6 = (Bal7z6[24] ^ N94nv6);
assign Met6z6 = (Igt6z6 & Qgt6z6);
assign Qgt6z6 = (~(Ygt6z6 & Uaanv6));
assign Ygt6z6 = (Kb4nv6 ^ Wx87z6);
assign Igt6z6 = (~(Ght6z6 & Eo9nv6));
assign Ght6z6 = (R44nv6 ^ Gkciw6);
assign Gkciw6 = (!Yw87z6);
assign Uat6z6 = (Oht6z6 & Wht6z6);
assign Wht6z6 = (Eit6z6 & Mit6z6);
assign Mit6z6 = (Uit6z6 & Cjt6z6);
assign Cjt6z6 = (~(Kjt6z6 & Sv9nv6));
assign Kjt6z6 = (Rb4nv6 ^ Qiciw6);
assign Qiciw6 = (!Gx87z6);
assign Uit6z6 = (~(Sjt6z6 & G3anv6));
assign Sjt6z6 = (Ki4nv6 ^ Ox87z6);
assign Eit6z6 = (Akt6z6 & Ikt6z6);
assign Ikt6z6 = (~(Qkt6z6 & Eganv6));
assign Qkt6z6 = (Jl4nv6 ^ Oaciw6);
assign Oaciw6 = (!Aw87z6);
assign Akt6z6 = (~(Ykt6z6 & Ju9nv6));
assign Ykt6z6 = (Ce4nv6 ^ N6ciw6);
assign N6ciw6 = (!Mu87z6);
assign Oht6z6 = (Glt6z6 & Olt6z6);
assign Olt6z6 = (~(Wlt6z6 & Qu9nv6));
assign Wlt6z6 = (Kv5nv6 ^ Tobiw6);
assign Tobiw6 = (!Eu87z6);
assign Glt6z6 = (Emt6z6 & Mmt6z6);
assign Mmt6z6 = (~(Umt6z6 & T6anv6));
assign Umt6z6 = (H64nv6 ^ I0ciw6);
assign I0ciw6 = (!Cv87z6);
assign Emt6z6 = (~(Q1anv6 & Cnt6z6));
assign Cnt6z6 = (Bal7z6[8] ^ Hk4nv6);
assign Eat6z6 = (Knt6z6 & Snt6z6);
assign Snt6z6 = (Aot6z6 & Iot6z6);
assign Iot6z6 = (Qot6z6 & Yot6z6);
assign Yot6z6 = (Gpt6z6 & Opt6z6);
assign Opt6z6 = (~(Wpt6z6 & Rcanv6));
assign Wpt6z6 = (U94nv6 ^ R0diw6);
assign R0diw6 = (!Kz87z6);
assign Gpt6z6 = (~(Eqt6z6 & Dy9nv6));
assign Eqt6z6 = (L4diw6 ^ Ico6z6);
assign L4diw6 = (!A097z6);
assign Qot6z6 = (Mqt6z6 & Uqt6z6);
assign Uqt6z6 = (~(Crt6z6 & Uhanv6));
assign Crt6z6 = (Ri4nv6 ^ Qw87z6);
assign Mqt6z6 = (~(Krt6z6 & K5anv6));
assign Krt6z6 = (Y44nv6 ^ Xpciw6);
assign Xpciw6 = (!Ey87z6);
assign Aot6z6 = (Srt6z6 & Ast6z6);
assign Ast6z6 = (~(Ist6z6 & Bbanv6));
assign Bbanv6 = (Eganv6 | Qst6z6);
assign Eganv6 = (~(Lo9nv6 & Yst6z6));
assign Yst6z6 = (~(Gtt6z6 & R5anv6));
assign Lo9nv6 = (!Vm9nv6);
assign Ist6z6 = (Je4nv6 ^ Lcciw6);
assign Lcciw6 = (!Iw87z6);
assign Srt6z6 = (Ott6z6 & Wtt6z6);
assign Wtt6z6 = (~(Eut6z6 & A0anv6));
assign A0anv6 = (!Ky9nv6);
assign Eut6z6 = (Gg4nv6 ^ Wl77z6);
assign Ott6z6 = (~(Mut6z6 & Vm9nv6));
assign Vm9nv6 = (~(Zv9nv6 & Uut6z6));
assign Uut6z6 = (~(Qst6z6 & Gtt6z6));
assign Zv9nv6 = (!Ju9nv6);
assign Ju9nv6 = (~(N3anv6 & Cvt6z6));
assign Cvt6z6 = (~(Kvt6z6 & R5anv6));
assign N3anv6 = (!E2anv6);
assign Mut6z6 = (Q74nv6 ^ Y8ciw6);
assign Y8ciw6 = (!Sv87z6);
assign Knt6z6 = (Svt6z6 & Awt6z6);
assign Awt6z6 = (Iwt6z6 & Qwt6z6);
assign Qwt6z6 = (Ywt6z6 & Gxt6z6);
assign Gxt6z6 = (~(Oxt6z6 & Gh36z6));
assign Oxt6z6 = (Hd4nv6 ^ Sybiw6);
assign Sybiw6 = (!Kv87z6);
assign Ywt6z6 = (~(Wxt6z6 & X1anv6));
assign X1anv6 = (Eyt6z6 & Qst6z6);
assign Eyt6z6 = (Myt6z6 & Gtt6z6);
assign Wxt6z6 = (Ak4nv6 ^ G936z6);
assign G936z6 = (!Bal7z6[5]);
assign Iwt6z6 = (Uyt6z6 & Czt6z6);
assign Czt6z6 = (~(Kzt6z6 & Cn9nv6));
assign Cn9nv6 = (Szt6z6 | Qu9nv6);
assign Qu9nv6 = (Q1anv6 & Gtt6z6);
assign Szt6z6 = (Qst6z6 & Myt6z6);
assign Kzt6z6 = (Tp5nv6 ^ Lrbiw6);
assign Lrbiw6 = (!Wt87z6);
assign Uyt6z6 = (~(A0u6z6 & E2anv6));
assign E2anv6 = (~(Om9nv6 & I0u6z6));
assign I0u6z6 = (~(Qst6z6 & Kvt6z6));
assign Om9nv6 = (!T6anv6);
assign T6anv6 = (~(Cu9nv6 & Q0u6z6));
assign Q0u6z6 = (~(Y0u6z6 & R5anv6));
assign Cu9nv6 = (!Gh36z6);
assign Gh36z6 = (~(G1u6z6 & Djanv6));
assign Djanv6 = (!Q1anv6);
assign Q1anv6 = (R5anv6 & Myt6z6);
assign G1u6z6 = (~(Qst6z6 & Y0u6z6));
assign Qst6z6 = (R5anv6 & O1u6z6);
assign A0u6z6 = (Cl4nv6 ^ A3ciw6);
assign A3ciw6 = (!Uu87z6);
assign Svt6z6 = (W1u6z6 & Uu36z6);
assign W1u6z6 = (E2u6z6 & M2u6z6);
assign M2u6z6 = (~(U2u6z6 & Bj9nv6));
assign Bj9nv6 = (!X8anv6);
assign X8anv6 = (Heanv6 & C3u6z6);
assign Heanv6 = (Rjanv6 & K3u6z6);
assign Rjanv6 = (!Dy9nv6);
assign Dy9nv6 = (~(Ui9nv6 & S3u6z6));
assign S3u6z6 = (~(Gtt6z6 & O1u6z6));
assign Ui9nv6 = (P6l7z6[3] & Iq9nv6);
assign Iq9nv6 = (!Rcanv6);
assign Rcanv6 = (~(Wx9nv6 & A4u6z6));
assign A4u6z6 = (~(Kvt6z6 & O1u6z6));
assign Wx9nv6 = (Ij9nv6 & I4u6z6);
assign I4u6z6 = (!Y0u6z6);
assign Ij9nv6 = (!Yk9nv6);
assign Yk9nv6 = (~(Wq9nv6 & Q4u6z6));
assign Q4u6z6 = (~(Y0u6z6 & O1u6z6));
assign Wq9nv6 = (Ky9nv6 & Y4u6z6);
assign Ky9nv6 = (~(K5anv6 | G5u6z6));
assign K5anv6 = (~(Fs9nv6 & O5u6z6));
assign O5u6z6 = (~(Gtt6z6 & Myt6z6));
assign Fs9nv6 = (!Uaanv6);
assign Uaanv6 = (~(Tz9nv6 & W5u6z6));
assign W5u6z6 = (~(G5u6z6 & Gtt6z6));
assign Tz9nv6 = (!Uhanv6);
assign Uhanv6 = (~(Fl9nv6 & E6u6z6));
assign E6u6z6 = (~(Kvt6z6 & Myt6z6));
assign Fl9nv6 = (!Eo9nv6);
assign Eo9nv6 = (~(Ts9nv6 & M6u6z6));
assign M6u6z6 = (~(G5u6z6 & Kvt6z6));
assign Ts9nv6 = (!Sv9nv6);
assign Sv9nv6 = (~(H0anv6 & U6u6z6));
assign U6u6z6 = (~(Y0u6z6 & Myt6z6));
assign H0anv6 = (!G3anv6);
assign G3anv6 = (~(Xn9nv6 & C7u6z6));
assign C7u6z6 = (~(G5u6z6 & Y0u6z6));
assign Y0u6z6 = (Gtt6z6 & Kvt6z6);
assign Gtt6z6 = (!K3u6z6);
assign K3u6z6 = (P6l7z6[2] & Uu36z6);
assign G5u6z6 = (O1u6z6 & Myt6z6);
assign Myt6z6 = (!Y4u6z6);
assign Y4u6z6 = (P6l7z6[4] & Uu36z6);
assign O1u6z6 = (!C3u6z6);
assign C3u6z6 = (P6l7z6[1] & Uu36z6);
assign U2u6z6 = (W34nv6 ^ My87z6);
assign E2u6z6 = (~(K7u6z6 & R5anv6));
assign R5anv6 = (!Xn9nv6);
assign Xn9nv6 = (P6l7z6[5] & Uu36z6);
assign Uu36z6 = (S7u6z6 & P6l7z6[0]);
assign S7u6z6 = (Sjy5z6 & A8u6z6);
assign A8u6z6 = (~(Luanv6 & Kvt6z6));
assign Kvt6z6 = (!P6l7z6[3]);
assign Luanv6 = (I8u6z6 & Q8u6z6);
assign Q8u6z6 = (!P6l7z6[5]);
assign I8u6z6 = (!P6l7z6[4]);
assign K7u6z6 = (~(Bal7z6[16] ^ J74nv6));
assign Wxo6z6 = (Y8u6z6 & G9u6z6);
assign G9u6z6 = (~(Mea6z6 & O9u6z6));
assign O9u6z6 = (~(W9u6z6 & Eau6z6));
assign Eau6z6 = (N1m7z6[22] ? Uau6z6 : Mau6z6);
assign Uau6z6 = (~(Ysn6z6 & Mau6z6));
assign Mau6z6 = (N1m7z6[21] | N1m7z6[20]);
assign W9u6z6 = (N1m7z6[21] ? Kbu6z6 : Cbu6z6);
assign Kbu6z6 = (Wtn6z6 | N1m7z6[20]);
assign Cbu6z6 = (~(N1m7z6[20] & Eun6z6));
assign Mea6z6 = (U6r6z6 & Sbu6z6);
assign U6r6z6 = (Acu6z6 & Icu6z6);
assign Icu6z6 = (Qcu6z6 & Ycu6z6);
assign Ycu6z6 = (Gdu6z6 & Odu6z6);
assign Odu6z6 = (Wdu6z6 & Eeu6z6);
assign Eeu6z6 = (~(C6met6 | Meu6z6));
assign Meu6z6 = (Ueu6z6 & Xk5nv6);
assign Xk5nv6 = (Cfu6z6 & Kfu6z6);
assign Cfu6z6 = (Sfu6z6 & Agu6z6);
assign Ueu6z6 = (Ak4nv6 ^ Wxz5z6);
assign Wxz5z6 = (!Z4m7z6[5]);
assign Wdu6z6 = (Igu6z6 & Qgu6z6);
assign Qgu6z6 = (~(Ygu6z6 & C65nv6));
assign C65nv6 = (Ghu6z6 | Qd5nv6);
assign Ghu6z6 = (Kfu6z6 & Agu6z6);
assign Ygu6z6 = (Tp5nv6 ^ Usbiw6);
assign Usbiw6 = (!U287z6);
assign Igu6z6 = (~(Ohu6z6 & Qd5nv6));
assign Qd5nv6 = (Qk5nv6 & Sfu6z6);
assign Ohu6z6 = (Kv5nv6 ^ Hpbiw6);
assign Hpbiw6 = (!C387z6);
assign Gdu6z6 = (Whu6z6 & Eiu6z6);
assign Eiu6z6 = (Miu6z6 & Uiu6z6);
assign Uiu6z6 = (~(Cju6z6 & Iu5nv6));
assign Iu5nv6 = (Sz5nv6 | Kfu6z6);
assign Cju6z6 = (Je4nv6 ^ Ndciw6);
assign Ndciw6 = (!G587z6);
assign Miu6z6 = (~(Kju6z6 & Sz5nv6));
assign Sz5nv6 = (~(L75nv6 & Sju6z6));
assign Sju6z6 = (~(Sfu6z6 & Ro5nv6));
assign L75nv6 = (!V55nv6);
assign Kju6z6 = (Jl4nv6 ^ Cbciw6);
assign Cbciw6 = (!Y487z6);
assign Whu6z6 = (Aku6z6 & Iku6z6);
assign Iku6z6 = (~(Qku6z6 & V55nv6));
assign V55nv6 = (~(Ze5nv6 & Yku6z6));
assign Yku6z6 = (~(Kfu6z6 & Sfu6z6));
assign Ze5nv6 = (!Jd5nv6);
assign Qku6z6 = (Q74nv6 ^ M9ciw6);
assign M9ciw6 = (!Q487z6);
assign Aku6z6 = (~(Glu6z6 & Jd5nv6));
assign Jd5nv6 = (~(Nm5nv6 & Olu6z6));
assign Olu6z6 = (~(Wlu6z6 & Ro5nv6));
assign Nm5nv6 = (!El5nv6);
assign Glu6z6 = (Ce4nv6 ^ P7ciw6);
assign P7ciw6 = (!K387z6);
assign Qcu6z6 = (Emu6z6 & Mmu6z6);
assign Mmu6z6 = (Umu6z6 & Cnu6z6);
assign Cnu6z6 = (Knu6z6 & Snu6z6);
assign Snu6z6 = (~(Aou6z6 & El5nv6));
assign El5nv6 = (~(O55nv6 & Iou6z6));
assign Iou6z6 = (~(Kfu6z6 & Wlu6z6));
assign O55nv6 = (!Aq5nv6);
assign Aou6z6 = (Cl4nv6 ^ Q4ciw6);
assign Q4ciw6 = (!S387z6);
assign Knu6z6 = (~(Qou6z6 & Aq5nv6));
assign Aq5nv6 = (~(Cd5nv6 & You6z6));
assign You6z6 = (~(Gpu6z6 & Ro5nv6));
assign Cd5nv6 = (!W506z6);
assign Qou6z6 = (H64nv6 ^ W0ciw6);
assign W0ciw6 = (!A487z6);
assign Umu6z6 = (Opu6z6 & Wpu6z6);
assign Wpu6z6 = (~(Equ6z6 & W506z6));
assign W506z6 = (~(Mqu6z6 & R26nv6));
assign R26nv6 = (!Qk5nv6);
assign Mqu6z6 = (~(Gpu6z6 & Kfu6z6));
assign Kfu6z6 = (Uqu6z6 & Ro5nv6);
assign Equ6z6 = (Hd4nv6 ^ Gzbiw6);
assign Gzbiw6 = (!I487z6);
assign Opu6z6 = (~(Qk5nv6 & Cru6z6));
assign Cru6z6 = (U606z6 ^ Ghp6z6);
assign U606z6 = (!Z4m7z6[8]);
assign Qk5nv6 = (Agu6z6 & Ro5nv6);
assign Emu6z6 = (Kru6z6 & Sru6z6);
assign Sru6z6 = (~(Asu6z6 & Dh5nv6));
assign Asu6z6 = (Z4diw6 ^ Ico6z6);
assign Z4diw6 = (!Y887z6);
assign Kru6z6 = (Isu6z6 & Qsu6z6);
assign Qsu6z6 = (~(Ysu6z6 & B25nv6));
assign B25nv6 = (!Es5nv6);
assign Es5nv6 = (Vx5nv6 & Gtu6z6);
assign Ysu6z6 = (W34nv6 ^ K787z6);
assign Isu6z6 = (~(Otu6z6 & P95nv6));
assign P95nv6 = (!Vx5nv6);
assign Vx5nv6 = (F36nv6 & Wtu6z6);
assign F36nv6 = (!Dh5nv6);
assign Dh5nv6 = (~(U15nv6 & Euu6z6));
assign Euu6z6 = (~(Sfu6z6 & Uqu6z6));
assign Otu6z6 = (Pa4nv6 ^ G987z6);
assign Acu6z6 = (Muu6z6 & Uuu6z6);
assign Uuu6z6 = (Cvu6z6 & Kvu6z6);
assign Kvu6z6 = (Svu6z6 & Awu6z6);
assign Awu6z6 = (Iwu6z6 & Qwu6z6);
assign Qwu6z6 = (~(Ywu6z6 & Ac06z6));
assign Ac06z6 = (!U15nv6);
assign U15nv6 = (N1m7z6[3] & I95nv6);
assign I95nv6 = (!Fw5nv6);
assign Ywu6z6 = (U24nv6 ^ J3diw6);
assign J3diw6 = (!Q887z6);
assign Iwu6z6 = (~(Gxu6z6 & Fw5nv6));
assign Fw5nv6 = (~(Wg5nv6 & Oxu6z6));
assign Oxu6z6 = (~(Wlu6z6 & Uqu6z6));
assign Gxu6z6 = (U94nv6 ^ F1diw6);
assign F1diw6 = (!I887z6);
assign Svu6z6 = (Wxu6z6 & Eyu6z6);
assign Eyu6z6 = (~(Myu6z6 & M36nv6));
assign M36nv6 = (!Wg5nv6);
assign Wg5nv6 = (I25nv6 & Uyu6z6);
assign Uyu6z6 = (!Gpu6z6);
assign I25nv6 = (!Y35nv6);
assign Myu6z6 = (Ng4nv6 ^ A887z6);
assign Wxu6z6 = (~(Czu6z6 & Y35nv6));
assign Y35nv6 = (~(W95nv6 & Kzu6z6));
assign Kzu6z6 = (~(Gpu6z6 & Uqu6z6));
assign Czu6z6 = (B34nv6 ^ S787z6);
assign Cvu6z6 = (Szu6z6 & A0v6z6);
assign A0v6z6 = (~(I0v6z6 & Ko5nv6));
assign I0v6z6 = (Y44nv6 ^ Lqciw6);
assign Lqciw6 = (!C787z6);
assign Szu6z6 = (Q0v6z6 & Y0v6z6);
assign Y0v6z6 = (~(G1v6z6 & Mb5nv6));
assign Mb5nv6 = (!W95nv6);
assign W95nv6 = (Kh5nv6 & O1v6z6);
assign G1v6z6 = (Sf06z6 ^ Ysp6z6);
assign Ysp6z6 = (!N94nv6);
assign Sf06z6 = (!Z4m7z6[24]);
assign Q0v6z6 = (~(W1v6z6 & Aj5nv6));
assign Aj5nv6 = (!Kh5nv6);
assign Kh5nv6 = (~(Ko5nv6 | E2v6z6));
assign Ko5nv6 = (~(Fb5nv6 & M2v6z6));
assign M2v6z6 = (~(Sfu6z6 & Agu6z6));
assign Fb5nv6 = (!Bu5nv6);
assign W1v6z6 = (Gg4nv6 ^ Gl77z6);
assign Muu6z6 = (U2v6z6 & C3v6z6);
assign C3v6z6 = (K3v6z6 & S3v6z6);
assign S3v6z6 = (A4v6z6 & I4v6z6);
assign I4v6z6 = (~(Q4v6z6 & Bu5nv6));
assign Bu5nv6 = (~(Ti5nv6 & Y4v6z6));
assign Y4v6z6 = (~(E2v6z6 & Sfu6z6));
assign Ti5nv6 = (!I16nv6);
assign Q4v6z6 = (Kb4nv6 ^ U687z6);
assign A4v6z6 = (~(G5v6z6 & I16nv6));
assign I16nv6 = (~(F45nv6 & O5v6z6));
assign O5v6z6 = (~(Wlu6z6 & Agu6z6));
assign F45nv6 = (!E75nv6);
assign G5v6z6 = (Ri4nv6 ^ O587z6);
assign K3v6z6 = (W5v6z6 & E6v6z6);
assign E6v6z6 = (~(M6v6z6 & E75nv6));
assign E75nv6 = (~(Tb5nv6 & U6v6z6));
assign U6v6z6 = (~(E2v6z6 & Wlu6z6));
assign Tb5nv6 = (!Se5nv6);
assign M6v6z6 = (R44nv6 ^ Ukciw6);
assign Ukciw6 = (!W587z6);
assign W5v6z6 = (~(C7v6z6 & Se5nv6));
assign Se5nv6 = (~(Hj5nv6 & K7v6z6));
assign K7v6z6 = (~(Gpu6z6 & Agu6z6));
assign Hj5nv6 = (!Gm5nv6);
assign C7v6z6 = (Rb4nv6 ^ Ejciw6);
assign Ejciw6 = (!E687z6);
assign U2v6z6 = (S7v6z6 & Ik06z6);
assign S7v6z6 = (A8v6z6 & I8v6z6);
assign I8v6z6 = (~(Q8v6z6 & Gm5nv6));
assign Gm5nv6 = (~(X65nv6 & Y8v6z6));
assign Y8v6z6 = (~(E2v6z6 & Gpu6z6));
assign Gpu6z6 = (Sfu6z6 & Wlu6z6);
assign Sfu6z6 = (!Wtu6z6);
assign Wtu6z6 = (N1m7z6[2] & Ik06z6);
assign E2v6z6 = (Uqu6z6 & Agu6z6);
assign Agu6z6 = (!O1v6z6);
assign O1v6z6 = (N1m7z6[4] & Ik06z6);
assign Uqu6z6 = (!Gtu6z6);
assign Gtu6z6 = (N1m7z6[1] & Ik06z6);
assign Q8v6z6 = (Ki4nv6 ^ M687z6);
assign A8v6z6 = (~(G9v6z6 & Ro5nv6));
assign Ro5nv6 = (!X65nv6);
assign X65nv6 = (N1m7z6[5] & Ik06z6);
assign Ik06z6 = (O9v6z6 & N1m7z6[0]);
assign O9v6z6 = (Sjy5z6 & W9v6z6);
assign W9v6z6 = (~(Zd6nv6 & Wlu6z6));
assign Wlu6z6 = (!N1m7z6[3]);
assign Zd6nv6 = (Eav6z6 & Mav6z6);
assign Mav6z6 = (!N1m7z6[5]);
assign Eav6z6 = (!N1m7z6[4]);
assign G9v6z6 = (Em06z6 ^ J74nv6);
assign Em06z6 = (!Z4m7z6[16]);
assign Y8u6z6 = (~(Aga6z6 & Uav6z6));
assign Uav6z6 = (~(Cbv6z6 & Kbv6z6));
assign Kbv6z6 = (Vbm7z6[22] ? Acv6z6 : Sbv6z6);
assign Acv6z6 = (~(Ysn6z6 & Sbv6z6));
assign Sbv6z6 = (Vbm7z6[21] | Vbm7z6[20]);
assign Cbv6z6 = (Vbm7z6[21] ? Qcv6z6 : Icv6z6);
assign Qcv6z6 = (Wtn6z6 | Vbm7z6[20]);
assign Wtn6z6 = (~(Eun6z6 & Ysn6z6));
assign Ysn6z6 = (I4a6z6 ? Lhmov6 : Qwget6);
assign Lhmov6 = (~(Ycv6z6 & Gdv6z6));
assign Gdv6z6 = (Odv6z6 & Wdv6z6);
assign Wdv6z6 = (Hjphw6 & J1a7x6);
assign Hjphw6 = (!Wxi6z6);
assign Odv6z6 = (X3yxx6 & Gwsiw6);
assign Gwsiw6 = (L8hhw6 | Dwb7z6[0]);
assign L8hhw6 = (~(Uakiy6 & Bwvnv6));
assign Ycv6z6 = (Eev6z6 & Mev6z6);
assign Mev6z6 = (Uev6z6 & Cfv6z6);
assign Uev6z6 = (Kfv6z6 | X4eet6);
assign Eev6z6 = (Sfv6z6 & Agv6z6);
assign Agv6z6 = (~(U6hiy6 & Dwb7z6[1]));
assign Sfv6z6 = (~(Ii9ov6 & Igv6z6));
assign Igv6z6 = (~(Qgv6z6 & Ygv6z6));
assign Qgv6z6 = (Ghv6z6 & Twphw6);
assign Ghv6z6 = (~(Ohv6z6 & Doihw6));
assign Ohv6z6 = (Dwb7z6[1] & Uvvnv6);
assign Icv6z6 = (~(Vbm7z6[20] & Eun6z6));
assign Eun6z6 = (!Glm6z6);
assign Glm6z6 = (P1het6 ? Dzget6 : Hjqnv6);
assign Hjqnv6 = (~(Whv6z6 & Eiv6z6));
assign Eiv6z6 = (~(N99iw6 & Miv6z6));
assign Miv6z6 = (Uiv6z6 | A0ghw6);
assign A0ghw6 = (!Ecc7z6[12]);
assign Uiv6z6 = (~(Tlmov6 & Pbadt6));
assign N99iw6 = (!Gbo6x6);
assign Gbo6x6 = (J2cdt6 & Tkbdt6);
assign Whv6z6 = (~(H7wxx6 & Gvvnv6));
assign Aga6z6 = (!Sbu6z6);
assign Sbu6z6 = (~(Cjv6z6 & Kjv6z6));
assign Kjv6z6 = (Sjv6z6 & Akv6z6);
assign Akv6z6 = (Ikv6z6 & Qkv6z6);
assign Qkv6z6 = (Ykv6z6 & Glv6z6);
assign Glv6z6 = (~(Cymet6 | Olv6z6));
assign Olv6z6 = (Wlv6z6 & En3nv6);
assign Wlv6z6 = (Pa4nv6 ^ Ey77z6);
assign Pa4nv6 = (P1het6 ? E6a6z6 : Yygnv6);
assign E6a6z6 = (!V5k7z6[30]);
assign Ykv6z6 = (Emv6z6 & Mmv6z6);
assign Mmv6z6 = (~(Umv6z6 & Ma66z6));
assign Ma66z6 = (!Oe3nv6);
assign Umv6z6 = (U24nv6 ^ Q3diw6);
assign Q3diw6 = (!Ox77z6);
assign U24nv6 = (P1het6 ? V5k7z6[28] : Cmm7z6[28]);
assign Emv6z6 = (~(Cnv6z6 & Su3nv6));
assign Cnv6z6 = (Ng4nv6 ^ Yw77z6);
assign Ng4nv6 = (P1het6 ? U297z6 : V0hnv6);
assign Ikv6z6 = (Knv6z6 & Snv6z6);
assign Snv6z6 = (Aov6z6 & Iov6z6);
assign Iov6z6 = (~(Qov6z6 & Jf3nv6));
assign Qov6z6 = (Kn66z6 ^ B34nv6);
assign B34nv6 = (P1het6 ? Knn6z6 : C1hnv6);
assign Knn6z6 = (!V5k7z6[25]);
assign Kn66z6 = (!Hfm7z6[25]);
assign Aov6z6 = (~(Yov6z6 & Bp3nv6));
assign Bp3nv6 = (!Xm3nv6);
assign Yov6z6 = (~(N94nv6 ^ Qw77z6));
assign N94nv6 = (P1het6 ? V5k7z6[24] : Cmm7z6[24]);
assign Knv6z6 = (Gpv6z6 & Opv6z6);
assign Opv6z6 = (~(Wpv6z6 & U676z6));
assign U676z6 = (!Uo3nv6);
assign Wpv6z6 = (Kb4nv6 ^ E287z6);
assign Kb4nv6 = (P1het6 ? Aon6z6 : E2hnv6);
assign Aon6z6 = (!V5k7z6[21]);
assign Gpv6z6 = (~(Eqv6z6 & Mk3nv6));
assign Eqv6z6 = (R44nv6 ^ Blciw6);
assign Blciw6 = (!O187z6);
assign R44nv6 = (P1het6 ? V5k7z6[19] : Cmm7z6[19]);
assign Sjv6z6 = (Mqv6z6 & Uqv6z6);
assign Uqv6z6 = (Crv6z6 & Krv6z6);
assign Krv6z6 = (Srv6z6 & Asv6z6);
assign Asv6z6 = (~(Isv6z6 & Vs3nv6));
assign Isv6z6 = (Rb4nv6 ^ Ljciw6);
assign Ljciw6 = (!O597z6);
assign Rb4nv6 = (P1het6 ? V5k7z6[18] : Cmm7z6[18]);
assign Srv6z6 = (~(Qsv6z6 & X04nv6));
assign Qsv6z6 = (Ki4nv6 ^ W187z6);
assign Ki4nv6 = (P1het6 ? Ui77z6 : I4hnv6);
assign I4hnv6 = (!Cmm7z6[17]);
assign Crv6z6 = (Ysv6z6 & Gtv6z6);
assign Gtv6z6 = (~(Otv6z6 & J04nv6));
assign Otv6z6 = (Jl4nv6 ^ Jbciw6);
assign Jbciw6 = (!Q087z6);
assign Jl4nv6 = (P1het6 ? V5k7z6[14] : Cmm7z6[14]);
assign Ysv6z6 = (~(Wtv6z6 & Mr3nv6));
assign Wtv6z6 = (Ce4nv6 ^ D8ciw6);
assign D8ciw6 = (!Cz77z6);
assign Ce4nv6 = (P1het6 ? V5k7z6[12] : Cmm7z6[12]);
assign Mqv6z6 = (Euv6z6 & Muv6z6);
assign Muv6z6 = (~(Uuv6z6 & Fr3nv6));
assign Uuv6z6 = (Kv5nv6 ^ Opbiw6);
assign Opbiw6 = (!Uy77z6);
assign Kv5nv6 = (P1het6 ? V5k7z6[6] : Cmm7z6[6]);
assign Euv6z6 = (Cvv6z6 & Kvv6z6);
assign Kvv6z6 = (~(Svv6z6 & Is56z6));
assign Is56z6 = (!Pi3nv6);
assign Svv6z6 = (H64nv6 ^ D1ciw6);
assign D1ciw6 = (!Sz77z6);
assign H64nv6 = (P1het6 ? V5k7z6[10] : Cmm7z6[10]);
assign Cvv6z6 = (~(Ty3nv6 & Awv6z6));
assign Awv6z6 = (G166z6 ^ Ghp6z6);
assign Ghp6z6 = (!Hk4nv6);
assign Hk4nv6 = (P1het6 ? V5k7z6[8] : Cmm7z6[8]);
assign G166z6 = (!Hfm7z6[8]);
assign Cjv6z6 = (Iwv6z6 & Qwv6z6);
assign Qwv6z6 = (Ywv6z6 & Gxv6z6);
assign Gxv6z6 = (Oxv6z6 & Wxv6z6);
assign Wxv6z6 = (Eyv6z6 & Myv6z6);
assign Myv6z6 = (~(Uyv6z6 & Qm3nv6));
assign Uyv6z6 = (U94nv6 ^ M1diw6);
assign M1diw6 = (!Gx77z6);
assign U94nv6 = (P1het6 ? V5k7z6[27] : Cmm7z6[27]);
assign Eyv6z6 = (~(Czv6z6 & Gv3nv6));
assign Czv6z6 = (G5diw6 ^ Ico6z6);
assign Ico6z6 = (~(M6a6z6 & Kzv6z6));
assign Kzv6z6 = (~(Cmm7z6[29] & I4a6z6));
assign I4a6z6 = (!P1het6);
assign M6a6z6 = (~(V5k7z6[29] & P1het6));
assign G5diw6 = (!Wx77z6);
assign Oxv6z6 = (Szv6z6 & A0w6z6);
assign A0w6z6 = (~(I0w6z6 & Ww3nv6));
assign I0w6z6 = (Ri4nv6 ^ G187z6);
assign Ri4nv6 = (P1het6 ? Cj77z6 : L2hnv6);
assign Szv6z6 = (~(Q0w6z6 & Zg3nv6));
assign Q0w6z6 = (Y44nv6 ^ Sqciw6);
assign Sqciw6 = (!M287z6);
assign Y44nv6 = (P1het6 ? V5k7z6[22] : Cmm7z6[22]);
assign Ywv6z6 = (Y0w6z6 & G1w6z6);
assign G1w6z6 = (~(O1w6z6 & Hs3nv6));
assign Hs3nv6 = (J04nv6 | W1w6z6);
assign J04nv6 = (~(Tk3nv6 & E2w6z6));
assign E2w6z6 = (~(M2w6z6 & Ys76z6));
assign Tk3nv6 = (!Wi3nv6);
assign O1w6z6 = (Je4nv6 ^ Udciw6);
assign Udciw6 = (!Y087z6);
assign Je4nv6 = (P1het6 ? V5k7z6[15] : Cmm7z6[15]);
assign Y0w6z6 = (U2w6z6 & C3w6z6);
assign C3w6z6 = (~(K3w6z6 & Kx3nv6));
assign Kx3nv6 = (!Zu3nv6);
assign K3w6z6 = (Gg4nv6 ^ Yk77z6);
assign Gg4nv6 = (P1het6 ? Kj77z6 : Q1hnv6);
assign U2w6z6 = (~(S3w6z6 & Wi3nv6));
assign Wi3nv6 = (~(Os3nv6 & A4w6z6));
assign A4w6z6 = (~(W1w6z6 & M2w6z6));
assign Os3nv6 = (!Mr3nv6);
assign Mr3nv6 = (~(Q04nv6 & I4w6z6));
assign I4w6z6 = (~(Q4w6z6 & Ys76z6));
assign Q04nv6 = (!Oz3nv6);
assign S3w6z6 = (Q74nv6 ^ T9ciw6);
assign T9ciw6 = (!I087z6);
assign Q74nv6 = (P1het6 ? V5k7z6[13] : Cmm7z6[13]);
assign Iwv6z6 = (Y4w6z6 & G5w6z6);
assign G5w6z6 = (O5w6z6 & W5w6z6);
assign W5w6z6 = (E6w6z6 & M6w6z6);
assign M6w6z6 = (~(U6w6z6 & Rq3nv6));
assign U6w6z6 = (Hd4nv6 ^ Nzbiw6);
assign Nzbiw6 = (!A087z6);
assign Hd4nv6 = (P1het6 ? V5k7z6[9] : Cmm7z6[9]);
assign E6w6z6 = (~(C7w6z6 & Hz3nv6));
assign Hz3nv6 = (K7w6z6 & W1w6z6);
assign K7w6z6 = (S7w6z6 & M2w6z6);
assign C7w6z6 = (Ak4nv6 ^ Mq46z6);
assign Mq46z6 = (!Hfm7z6[5]);
assign Ak4nv6 = (!Ci7nv6);
assign Ci7nv6 = (P1het6 ? V5k7z6[5] : Cmm7z6[5]);
assign O5w6z6 = (A8w6z6 & I8w6z6);
assign I8w6z6 = (~(Q8w6z6 & Dj3nv6));
assign Dj3nv6 = (Y8w6z6 | Fr3nv6);
assign Fr3nv6 = (Ty3nv6 & M2w6z6);
assign Y8w6z6 = (W1w6z6 & S7w6z6);
assign Q8w6z6 = (Tp5nv6 ^ Btbiw6);
assign Btbiw6 = (!My77z6);
assign Tp5nv6 = (P1het6 ? V5k7z6[7] : Cmm7z6[7]);
assign A8w6z6 = (~(G9w6z6 & Oz3nv6));
assign Oz3nv6 = (~(Pi3nv6 & O9w6z6));
assign O9w6z6 = (~(W1w6z6 & Q4w6z6));
assign Pi3nv6 = (~(Rq3nv6 | W9w6z6));
assign W9w6z6 = (Eaw6z6 & Ys76z6);
assign Rq3nv6 = (Maw6z6 | Ty3nv6);
assign Ty3nv6 = (Ys76z6 & S7w6z6);
assign Maw6z6 = (W1w6z6 & Eaw6z6);
assign W1w6z6 = (Ys76z6 & Uaw6z6);
assign G9w6z6 = (Cl4nv6 ^ X4ciw6);
assign X4ciw6 = (!Kz77z6);
assign Cl4nv6 = (P1het6 ? V5k7z6[11] : Cmm7z6[11]);
assign Y4w6z6 = (Cbw6z6 & Sn76z6);
assign Cbw6z6 = (Kbw6z6 & Sbw6z6);
assign Sbw6z6 = (~(Acw6z6 & Ve3nv6));
assign Ve3nv6 = (En3nv6 | Uaw6z6);
assign En3nv6 = (Gv3nv6 | M2w6z6);
assign Gv3nv6 = (~(Oe3nv6 & Icw6z6));
assign Icw6z6 = (~(M2w6z6 & Uaw6z6));
assign Oe3nv6 = (~(Q4w6z6 | Qm3nv6));
assign Qm3nv6 = (Su3nv6 | Qcw6z6);
assign Qcw6z6 = (~(Vbm7z6[3] | Ycw6z6));
assign Su3nv6 = (Jf3nv6 | Eaw6z6);
assign Jf3nv6 = (~(Xm3nv6 & Gdw6z6));
assign Gdw6z6 = (~(Eaw6z6 & Uaw6z6));
assign Xm3nv6 = (Zu3nv6 & Odw6z6);
assign Zu3nv6 = (~(Zg3nv6 | Wdw6z6));
assign Zg3nv6 = (~(Uo3nv6 & Eew6z6));
assign Eew6z6 = (~(M2w6z6 & S7w6z6));
assign Uo3nv6 = (~(Ww3nv6 | Mew6z6));
assign Mew6z6 = (Wdw6z6 & M2w6z6);
assign Ww3nv6 = (~(Gh3nv6 & Uew6z6));
assign Uew6z6 = (~(Q4w6z6 & S7w6z6));
assign Gh3nv6 = (!Mk3nv6);
assign Mk3nv6 = (~(Ip3nv6 & Cfw6z6));
assign Cfw6z6 = (~(Wdw6z6 & Q4w6z6));
assign Ip3nv6 = (!Vs3nv6);
assign Vs3nv6 = (~(Dx3nv6 & Kfw6z6));
assign Kfw6z6 = (~(Eaw6z6 & S7w6z6));
assign Dx3nv6 = (!X04nv6);
assign X04nv6 = (~(Fk3nv6 & Sfw6z6));
assign Sfw6z6 = (~(Wdw6z6 & Eaw6z6));
assign Eaw6z6 = (M2w6z6 & Q4w6z6);
assign M2w6z6 = (~(Vbm7z6[2] & Sn76z6));
assign Wdw6z6 = (Uaw6z6 & S7w6z6);
assign S7w6z6 = (!Odw6z6);
assign Odw6z6 = (Vbm7z6[4] & Sn76z6);
assign Uaw6z6 = (!Ycw6z6);
assign Ycw6z6 = (Vbm7z6[1] & Sn76z6);
assign Acw6z6 = (W34nv6 ^ Iw77z6);
assign W34nv6 = (!Agw6z6);
assign Agw6z6 = (P1het6 ? V5k7z6[31] : Cmm7z6[31]);
assign Kbw6z6 = (~(Igw6z6 & Ys76z6));
assign Ys76z6 = (!Fk3nv6);
assign Fk3nv6 = (Vbm7z6[5] & Sn76z6);
assign Sn76z6 = (Qgw6z6 & Vbm7z6[0]);
assign Qgw6z6 = (Sjy5z6 & Ygw6z6);
assign Ygw6z6 = (~(Wv4nv6 & Q4w6z6));
assign Q4w6z6 = (!Vbm7z6[3]);
assign Wv4nv6 = (Ghw6z6 & Ohw6z6);
assign Ohw6z6 = (!Vbm7z6[5]);
assign Ghw6z6 = (!Vbm7z6[4]);
assign Igw6z6 = (Gt76z6 ^ J74nv6);
assign J74nv6 = (P1het6 ? Snm6z6 : P4hnv6);
assign Snm6z6 = (!V5k7z6[16]);
assign P4hnv6 = (!Cmm7z6[16]);
assign Gt76z6 = (!Hfm7z6[16]);
assign Sjy5z6 = (Phget6 & Whw6z6);
assign Whw6z6 = (Weget6 | Etinv6);
assign Etinv6 = (Dxgov6 & Ev2nv6);
assign Ev2nv6 = (!Fjadt6);
assign Dxgov6 = (S34jy6 & Cn2nv6);
assign Cn2nv6 = (!X3get6);
assign S34jy6 = (!Inadt6);
assign Ein6z6 = (~(Zmnyx6 & L3bdt6));
assign HMASTERS[0] = (~(Eiw6z6 & Miw6z6));
assign Miw6z6 = (~(Uiw6z6 & Cjw6z6));
assign Uiw6z6 = (K6uet6 & J0jxx6);
assign Eiw6z6 = (~(Fk9ov6 & T52iw6));
assign HMASTERD[0] = (~(Kjw6z6 & Sjw6z6));
assign Sjw6z6 = (~(Akw6z6 & Cjw6z6));
assign Cjw6z6 = (Ikw6z6 & Ewyet6);
assign Akw6z6 = (K6uet6 & Jn1ov6);
assign Kjw6z6 = (~(Vm1ov6 & T52iw6));
assign T52iw6 = (Zn0ft6 | Lq0ft6);
assign HBURSTS[0] = (~(Qkw6z6 & Ykw6z6));
assign Ykw6z6 = (~(J0jxx6 & Glw6z6));
assign Glw6z6 = (Vugxx6 | Jinyx6);
assign Qkw6z6 = (En9ov6 & Cfonv6);
assign HBURSTD[0] = (~(Ibonv6 & Jfonv6));
assign HADDRS[9] = (~(Olw6z6 & Wlw6z6));
assign Wlw6z6 = (Emw6z6 & Mmw6z6);
assign Mmw6z6 = (~(S7m6z6 & Cmm7z6[14]));
assign Emw6z6 = (Umw6z6 & Cnw6z6);
assign Cnw6z6 = (~(Mma6z6 & Fvb7z6[9]));
assign Umw6z6 = (~(Zmnyx6 & Fvb7z6[14]));
assign Olw6z6 = (Knw6z6 & Snw6z6);
assign Snw6z6 = (~(Aoa6z6 & Cmm7z6[9]));
assign Knw6z6 = (~(Onret6 & J0jxx6));
assign HADDRS[8] = (~(Aow6z6 & Iow6z6));
assign Iow6z6 = (Qow6z6 & Yow6z6);
assign Yow6z6 = (~(S7m6z6 & Cmm7z6[13]));
assign Qow6z6 = (Gpw6z6 & Opw6z6);
assign Opw6z6 = (~(Mma6z6 & Fvb7z6[8]));
assign Gpw6z6 = (~(Zmnyx6 & Fvb7z6[13]));
assign Aow6z6 = (Wpw6z6 & Eqw6z6);
assign Eqw6z6 = (~(Aoa6z6 & Cmm7z6[8]));
assign Wpw6z6 = (~(Ppret6 & J0jxx6));
assign HADDRS[7] = (~(Mqw6z6 & Uqw6z6));
assign Uqw6z6 = (Crw6z6 & Krw6z6);
assign Krw6z6 = (~(S7m6z6 & Cmm7z6[12]));
assign Crw6z6 = (Srw6z6 & Asw6z6);
assign Asw6z6 = (~(Mma6z6 & Fvb7z6[7]));
assign Srw6z6 = (~(Zmnyx6 & Fvb7z6[12]));
assign Mqw6z6 = (Isw6z6 & Qsw6z6);
assign Qsw6z6 = (~(Aoa6z6 & Cmm7z6[7]));
assign Isw6z6 = (~(Qrret6 & J0jxx6));
assign HADDRS[6] = (~(Ysw6z6 & Gtw6z6));
assign Gtw6z6 = (Otw6z6 & Wtw6z6);
assign Wtw6z6 = (~(S7m6z6 & Cmm7z6[11]));
assign Otw6z6 = (Euw6z6 & Muw6z6);
assign Muw6z6 = (~(Mma6z6 & Fvb7z6[6]));
assign Euw6z6 = (~(Zmnyx6 & Fvb7z6[11]));
assign Ysw6z6 = (Uuw6z6 & Cvw6z6);
assign Cvw6z6 = (~(Aoa6z6 & Cmm7z6[6]));
assign Uuw6z6 = (~(Rtret6 & J0jxx6));
assign HADDRS[5] = (~(Kvw6z6 & Svw6z6));
assign Svw6z6 = (Aww6z6 & Iww6z6);
assign Iww6z6 = (~(S7m6z6 & Cmm7z6[10]));
assign Aww6z6 = (Qww6z6 & Yww6z6);
assign Yww6z6 = (~(Mma6z6 & Fvb7z6[5]));
assign Qww6z6 = (~(Zmnyx6 & Fvb7z6[10]));
assign Kvw6z6 = (Gxw6z6 & Oxw6z6);
assign Oxw6z6 = (~(Aoa6z6 & Cmm7z6[5]));
assign Gxw6z6 = (~(Svret6 & J0jxx6));
assign HADDRS[4] = (~(Wxw6z6 & Eyw6z6));
assign Eyw6z6 = (Myw6z6 & Uyw6z6);
assign Uyw6z6 = (~(S7m6z6 & Cmm7z6[9]));
assign Myw6z6 = (Czw6z6 & Kzw6z6);
assign Kzw6z6 = (~(Mma6z6 & Fvb7z6[4]));
assign Czw6z6 = (~(Zmnyx6 & Fvb7z6[9]));
assign Wxw6z6 = (Szw6z6 & A0x6z6);
assign A0x6z6 = (~(Aoa6z6 & Cmm7z6[4]));
assign Szw6z6 = (~(Txret6 & J0jxx6));
assign HADDRS[3] = (~(I0x6z6 & Q0x6z6));
assign Q0x6z6 = (Y0x6z6 & G1x6z6);
assign G1x6z6 = (~(S7m6z6 & Cmm7z6[8]));
assign Y0x6z6 = (O1x6z6 & W1x6z6);
assign W1x6z6 = (~(Mma6z6 & Fvb7z6[3]));
assign O1x6z6 = (~(Zmnyx6 & Fvb7z6[8]));
assign I0x6z6 = (E2x6z6 & M2x6z6);
assign M2x6z6 = (~(Aoa6z6 & Cmm7z6[3]));
assign E2x6z6 = (~(Uzret6 & J0jxx6));
assign HADDRS[31] = (~(U2x6z6 & C3x6z6));
assign C3x6z6 = (~(Seqet6 & J0jxx6));
assign U2x6z6 = (K3x6z6 & S3x6z6);
assign S3x6z6 = (~(Fk9ov6 & Fvb7z6[31]));
assign K3x6z6 = (~(Rj9ov6 & Cmm7z6[31]));
assign HADDRS[30] = (~(A4x6z6 & I4x6z6));
assign I4x6z6 = (~(Tgqet6 & J0jxx6));
assign A4x6z6 = (Q4x6z6 & Y4x6z6);
assign Y4x6z6 = (~(Fk9ov6 & Fvb7z6[30]));
assign Q4x6z6 = (~(Rj9ov6 & Cmm7z6[30]));
assign HADDRS[2] = (~(G5x6z6 & O5x6z6));
assign O5x6z6 = (W5x6z6 & E6x6z6);
assign E6x6z6 = (~(S7m6z6 & Cmm7z6[7]));
assign W5x6z6 = (M6x6z6 & U6x6z6);
assign U6x6z6 = (~(Mma6z6 & Fvb7z6[2]));
assign M6x6z6 = (~(Zmnyx6 & Fvb7z6[7]));
assign G5x6z6 = (C7x6z6 & K7x6z6);
assign K7x6z6 = (~(Aoa6z6 & Yefnv6));
assign C7x6z6 = (~(V1set6 & J0jxx6));
assign HADDRS[29] = (~(S7x6z6 & A8x6z6));
assign A8x6z6 = (~(Uiqet6 & J0jxx6));
assign S7x6z6 = (I8x6z6 & Q8x6z6);
assign Q8x6z6 = (~(Fk9ov6 & Fvb7z6[29]));
assign I8x6z6 = (~(Rj9ov6 & Cmm7z6[29]));
assign HADDRS[28] = (~(Y8x6z6 & G9x6z6));
assign G9x6z6 = (~(Vkqet6 & J0jxx6));
assign Y8x6z6 = (O9x6z6 & W9x6z6);
assign W9x6z6 = (~(Fvb7z6[28] & Fk9ov6));
assign O9x6z6 = (~(Rj9ov6 & Cmm7z6[28]));
assign HADDRS[27] = (~(Eax6z6 & Max6z6));
assign Max6z6 = (~(Wmqet6 & J0jxx6));
assign Eax6z6 = (Uax6z6 & Cbx6z6);
assign Cbx6z6 = (~(Mma6z6 & Fvb7z6[27]));
assign Uax6z6 = (~(Aoa6z6 & Cmm7z6[27]));
assign HADDRS[26] = (~(Kbx6z6 & Sbx6z6));
assign Sbx6z6 = (~(Xoqet6 & J0jxx6));
assign Kbx6z6 = (Acx6z6 & Icx6z6);
assign Icx6z6 = (~(Mma6z6 & Fvb7z6[26]));
assign Acx6z6 = (~(Aoa6z6 & Cmm7z6[26]));
assign HADDRS[25] = (~(Qcx6z6 & Ycx6z6));
assign Ycx6z6 = (~(Yqqet6 & J0jxx6));
assign Qcx6z6 = (Gdx6z6 & Odx6z6);
assign Odx6z6 = (~(Mma6z6 & Fvb7z6[25]));
assign Gdx6z6 = (~(Aoa6z6 & Cmm7z6[25]));
assign HADDRS[24] = (~(Wdx6z6 & Eex6z6));
assign Eex6z6 = (~(Zsqet6 & J0jxx6));
assign Wdx6z6 = (Mex6z6 & Uex6z6);
assign Uex6z6 = (~(Mma6z6 & Fvb7z6[24]));
assign Mex6z6 = (~(Aoa6z6 & Cmm7z6[24]));
assign HADDRS[23] = (~(Cfx6z6 & Kfx6z6));
assign Kfx6z6 = (~(Avqet6 & J0jxx6));
assign Cfx6z6 = (Sfx6z6 & Agx6z6);
assign Agx6z6 = (~(Mma6z6 & Fvb7z6[23]));
assign Sfx6z6 = (~(Aoa6z6 & Cmm7z6[23]));
assign HADDRS[22] = (~(Igx6z6 & Qgx6z6));
assign Qgx6z6 = (~(Bxqet6 & J0jxx6));
assign Igx6z6 = (Ygx6z6 & Ghx6z6);
assign Ghx6z6 = (~(Mma6z6 & Fvb7z6[22]));
assign Ygx6z6 = (~(Aoa6z6 & Cmm7z6[22]));
assign HADDRS[21] = (~(Ohx6z6 & Whx6z6));
assign Whx6z6 = (~(Czqet6 & J0jxx6));
assign Ohx6z6 = (Eix6z6 & Mix6z6);
assign Mix6z6 = (~(Mma6z6 & Fvb7z6[21]));
assign Eix6z6 = (~(Aoa6z6 & Cmm7z6[21]));
assign HADDRS[20] = (~(Uix6z6 & Cjx6z6));
assign Cjx6z6 = (~(D1ret6 & J0jxx6));
assign Uix6z6 = (Kjx6z6 & Sjx6z6);
assign Sjx6z6 = (~(Mma6z6 & Fvb7z6[20]));
assign Kjx6z6 = (~(Aoa6z6 & Cmm7z6[20]));
assign HADDRS[1] = (~(Akx6z6 & Ikx6z6));
assign Ikx6z6 = (Qkx6z6 & Ykx6z6);
assign Ykx6z6 = (~(Mma6z6 & Stpnv6));
assign Qkx6z6 = (Glx6z6 & Olx6z6);
assign Olx6z6 = (~(Wlx6z6 & S7m6z6));
assign Wlx6z6 = (Cmm7z6[6] & Emx6z6);
assign Emx6z6 = (~(Anehw6 & Ta4iw6));
assign Glx6z6 = (~(Mmx6z6 & Zmnyx6));
assign Mmx6z6 = (Fvb7z6[6] & Ohe7x6);
assign Ohe7x6 = (Jie7x6 | Hub7z6[0]);
assign Akx6z6 = (Umx6z6 & Cnx6z6);
assign Cnx6z6 = (~(Aoa6z6 & Cmm7z6[1]));
assign Umx6z6 = (~(W3set6 & J0jxx6));
assign HADDRS[19] = (~(Knx6z6 & Snx6z6));
assign Snx6z6 = (Aox6z6 & Iox6z6);
assign Iox6z6 = (~(S7m6z6 & Cmm7z6[24]));
assign Aox6z6 = (Qox6z6 & Yox6z6);
assign Yox6z6 = (~(Mma6z6 & Fvb7z6[19]));
assign Qox6z6 = (~(Zmnyx6 & Fvb7z6[24]));
assign Knx6z6 = (Gpx6z6 & Opx6z6);
assign Opx6z6 = (~(Aoa6z6 & Cmm7z6[19]));
assign Gpx6z6 = (~(E3ret6 & J0jxx6));
assign HADDRS[18] = (~(Wpx6z6 & Eqx6z6));
assign Eqx6z6 = (Mqx6z6 & Uqx6z6);
assign Uqx6z6 = (~(S7m6z6 & Cmm7z6[23]));
assign Mqx6z6 = (Crx6z6 & Krx6z6);
assign Krx6z6 = (~(Mma6z6 & Fvb7z6[18]));
assign Crx6z6 = (~(Zmnyx6 & Fvb7z6[23]));
assign Wpx6z6 = (Srx6z6 & Asx6z6);
assign Asx6z6 = (~(Aoa6z6 & Cmm7z6[18]));
assign Srx6z6 = (~(F5ret6 & J0jxx6));
assign HADDRS[17] = (~(Isx6z6 & Qsx6z6));
assign Qsx6z6 = (Ysx6z6 & Gtx6z6);
assign Gtx6z6 = (~(S7m6z6 & Cmm7z6[22]));
assign Ysx6z6 = (Otx6z6 & Wtx6z6);
assign Wtx6z6 = (~(Mma6z6 & Fvb7z6[17]));
assign Otx6z6 = (~(Zmnyx6 & Fvb7z6[22]));
assign Isx6z6 = (Eux6z6 & Mux6z6);
assign Mux6z6 = (~(Aoa6z6 & Cmm7z6[17]));
assign Eux6z6 = (~(G7ret6 & J0jxx6));
assign HADDRS[16] = (~(Uux6z6 & Cvx6z6));
assign Cvx6z6 = (Kvx6z6 & Svx6z6);
assign Svx6z6 = (~(S7m6z6 & Cmm7z6[21]));
assign Kvx6z6 = (Awx6z6 & Iwx6z6);
assign Iwx6z6 = (~(Mma6z6 & Fvb7z6[16]));
assign Awx6z6 = (~(Zmnyx6 & Fvb7z6[21]));
assign Uux6z6 = (Qwx6z6 & Ywx6z6);
assign Ywx6z6 = (~(Aoa6z6 & Cmm7z6[16]));
assign Qwx6z6 = (~(H9ret6 & J0jxx6));
assign HADDRS[15] = (~(Gxx6z6 & Oxx6z6));
assign Oxx6z6 = (Wxx6z6 & Eyx6z6);
assign Eyx6z6 = (~(S7m6z6 & Cmm7z6[20]));
assign Wxx6z6 = (Myx6z6 & Uyx6z6);
assign Uyx6z6 = (~(Mma6z6 & Fvb7z6[15]));
assign Myx6z6 = (~(Zmnyx6 & Fvb7z6[20]));
assign Gxx6z6 = (Czx6z6 & Kzx6z6);
assign Kzx6z6 = (~(Aoa6z6 & Cmm7z6[15]));
assign Czx6z6 = (~(Ibret6 & J0jxx6));
assign HADDRS[14] = (~(Szx6z6 & A0y6z6));
assign A0y6z6 = (I0y6z6 & Q0y6z6);
assign Q0y6z6 = (~(S7m6z6 & Cmm7z6[19]));
assign I0y6z6 = (Y0y6z6 & G1y6z6);
assign G1y6z6 = (~(Mma6z6 & Fvb7z6[14]));
assign Y0y6z6 = (~(Zmnyx6 & Fvb7z6[19]));
assign Szx6z6 = (O1y6z6 & W1y6z6);
assign W1y6z6 = (~(Aoa6z6 & Cmm7z6[14]));
assign O1y6z6 = (~(Jdret6 & J0jxx6));
assign HADDRS[13] = (~(E2y6z6 & M2y6z6));
assign M2y6z6 = (U2y6z6 & C3y6z6);
assign C3y6z6 = (~(S7m6z6 & Cmm7z6[18]));
assign U2y6z6 = (K3y6z6 & S3y6z6);
assign S3y6z6 = (~(Mma6z6 & Fvb7z6[13]));
assign K3y6z6 = (~(Zmnyx6 & Fvb7z6[18]));
assign E2y6z6 = (A4y6z6 & I4y6z6);
assign I4y6z6 = (~(Aoa6z6 & Cmm7z6[13]));
assign A4y6z6 = (~(Kfret6 & J0jxx6));
assign HADDRS[12] = (~(Q4y6z6 & Y4y6z6));
assign Y4y6z6 = (G5y6z6 & O5y6z6);
assign O5y6z6 = (~(S7m6z6 & Cmm7z6[17]));
assign G5y6z6 = (W5y6z6 & E6y6z6);
assign E6y6z6 = (~(Mma6z6 & Fvb7z6[12]));
assign W5y6z6 = (~(Zmnyx6 & Fvb7z6[17]));
assign Q4y6z6 = (M6y6z6 & U6y6z6);
assign U6y6z6 = (~(Aoa6z6 & Cmm7z6[12]));
assign M6y6z6 = (~(Lhret6 & J0jxx6));
assign HADDRS[11] = (~(C7y6z6 & K7y6z6));
assign K7y6z6 = (S7y6z6 & A8y6z6);
assign A8y6z6 = (~(S7m6z6 & Cmm7z6[16]));
assign S7y6z6 = (I8y6z6 & Q8y6z6);
assign Q8y6z6 = (~(Mma6z6 & Fvb7z6[11]));
assign I8y6z6 = (~(Zmnyx6 & Fvb7z6[16]));
assign C7y6z6 = (Y8y6z6 & G9y6z6);
assign G9y6z6 = (~(Aoa6z6 & Cmm7z6[11]));
assign Y8y6z6 = (~(Mjret6 & J0jxx6));
assign HADDRS[10] = (~(O9y6z6 & W9y6z6));
assign W9y6z6 = (Eay6z6 & May6z6);
assign May6z6 = (~(S7m6z6 & Cmm7z6[15]));
assign Eay6z6 = (Uay6z6 & Cby6z6);
assign Cby6z6 = (~(Mma6z6 & Fvb7z6[10]));
assign Uay6z6 = (~(Zmnyx6 & Fvb7z6[15]));
assign O9y6z6 = (Kby6z6 & Sby6z6);
assign Sby6z6 = (~(Aoa6z6 & Cmm7z6[10]));
assign Kby6z6 = (~(Nlret6 & J0jxx6));
assign HADDRS[0] = (~(Acy6z6 & Icy6z6));
assign Icy6z6 = (Qcy6z6 & Ycy6z6);
assign Ycy6z6 = (~(Mma6z6 & Mbqnv6));
assign Mma6z6 = (Fk9ov6 & E2ziy6);
assign Fk9ov6 = (!Zn9ov6);
assign Qcy6z6 = (Gdy6z6 & Ody6z6);
assign Ody6z6 = (~(Wdy6z6 & Eey6z6));
assign Eey6z6 = (M6giy6 & Jie7x6);
assign Jie7x6 = (!Hub7z6[1]);
assign M6giy6 = (!Hub7z6[0]);
assign Wdy6z6 = (Zmnyx6 & Fvb7z6[5]);
assign Zmnyx6 = (!En9ov6);
assign En9ov6 = (Zn9ov6 | E2ziy6);
assign Zn9ov6 = (~(Mey6z6 & Uey6z6));
assign Uey6z6 = (Cfy6z6 & Kfy6z6);
assign Cfy6z6 = (Oz1iw6 & Uaonv6);
assign Oz1iw6 = (~(Sfy6z6 & Agy6z6));
assign Agy6z6 = (Igy6z6 & Qgy6z6);
assign Qgy6z6 = (Ygy6z6 & Ghy6z6);
assign Ygy6z6 = (~(Fvb7z6[27] | Fvb7z6[28]));
assign Igy6z6 = (~(Ohy6z6 | Fvb7z6[23]));
assign Ohy6z6 = (Fvb7z6[24] | Fvb7z6[25]);
assign Sfy6z6 = (Why6z6 & Eiy6z6);
assign Eiy6z6 = (~(Miy6z6 | Fvb7z6[20]));
assign Miy6z6 = (Fvb7z6[21] | Fvb7z6[22]);
assign Why6z6 = (Uiy6z6 & Fvb7z6[31]);
assign Uiy6z6 = (Fvb7z6[29] & Fvb7z6[30]);
assign Mey6z6 = (Cjy6z6 & Hz1iw6);
assign Hz1iw6 = (K4bdt6 & Kjy6z6);
assign Cjy6z6 = (Sjy6z6 & Aky6z6);
assign Aky6z6 = (~(Gazet6 & Iky6z6));
assign Iky6z6 = (Kyn7z6[0] | Kyn7z6[2]);
assign Sjy6z6 = (~(Qky6z6 & Yky6z6));
assign Yky6z6 = (~(Gly6z6 & Oly6z6));
assign Oly6z6 = (Wly6z6 & Dhnyx6);
assign Wly6z6 = (~(Aoyiy6 | Khoet6));
assign Gly6z6 = (Emy6z6 & Mmy6z6);
assign Mmy6z6 = (~(Ewyet6 & Qln7z6[0]));
assign Gdy6z6 = (~(Umy6z6 & Cny6z6));
assign Cny6z6 = (Cmm7z6[5] & Ta4iw6);
assign Umy6z6 = (S7m6z6 & Pbhnv6);
assign Pbhnv6 = (!Anehw6);
assign S7m6z6 = (!U2m6z6);
assign U2m6z6 = (Sgonv6 | Cfonv6);
assign Cfonv6 = (!Rj9ov6);
assign Acy6z6 = (Kny6z6 & Sny6z6);
assign Sny6z6 = (~(Aoa6z6 & Cmm7z6[0]));
assign Aoa6z6 = (!G5m6z6);
assign G5m6z6 = (~(Rj9ov6 & Sgonv6));
assign Kny6z6 = (~(X5set6 & J0jxx6));
assign HADDRI[4] = (Lhmyx6 ? X0d7z6[4] : Dvc7z6[4]);
assign X0d7z6[4] = (~(Aoy6z6 & Ioy6z6));
assign Ioy6z6 = (Qoy6z6 & Yoy6z6);
assign Yoy6z6 = (~(Pic7z6[4] & Ir0ov6));
assign Qoy6z6 = (Gpy6z6 & Opy6z6);
assign Opy6z6 = (Qs46z6 | Li0ov6);
assign Li0ov6 = (Wpy6z6 & Eqy6z6);
assign Eqy6z6 = (~(Wkd7z6[4] & Ddmhw6));
assign Wpy6z6 = (Mqy6z6 & Uqy6z6);
assign Uqy6z6 = (~(Xhd7z6[4] & Eu46z6));
assign Mqy6z6 = (~(Vnd7z6[4] & Jamnv6));
assign Gpy6z6 = (~(Pdc7z6[4] & Mu46z6));
assign Aoy6z6 = (Cry6z6 & Kry6z6);
assign Kry6z6 = (~(Znnov6 & P2j7z6[2]));
assign Cry6z6 = (~(Qdcdt6 & E3c7z6[4]));
assign HADDRI[3] = (Lhmyx6 ? X0d7z6[3] : Dvc7z6[3]);
assign X0d7z6[3] = (~(Sry6z6 & Asy6z6));
assign Asy6z6 = (Isy6z6 & Qsy6z6);
assign Qsy6z6 = (~(Pic7z6[3] & Ir0ov6));
assign Isy6z6 = (Ysy6z6 & Gty6z6);
assign Gty6z6 = (Qs46z6 | Mm0ov6);
assign Mm0ov6 = (Oty6z6 & Wty6z6);
assign Wty6z6 = (~(Wkd7z6[3] & Ddmhw6));
assign Oty6z6 = (Euy6z6 & Muy6z6);
assign Muy6z6 = (~(Xhd7z6[3] & Eu46z6));
assign Euy6z6 = (~(Vnd7z6[3] & Jamnv6));
assign Ysy6z6 = (~(Pdc7z6[3] & Mu46z6));
assign Sry6z6 = (Uuy6z6 & Cvy6z6);
assign Cvy6z6 = (~(Znnov6 & P2j7z6[1]));
assign Uuy6z6 = (~(Qdcdt6 & E3c7z6[3]));
assign HADDRI[2] = (Lhmyx6 ? X0d7z6[2] : Dvc7z6[2]);
assign Lhmyx6 = (!Crcdt6);
assign X0d7z6[2] = (~(Kvy6z6 & Svy6z6));
assign Svy6z6 = (Awy6z6 & Iwy6z6);
assign Iwy6z6 = (~(Pdc7z6[2] & Mu46z6));
assign Awy6z6 = (Qwy6z6 & R537x6);
assign Qwy6z6 = (Qs46z6 | Rs0ov6);
assign Rs0ov6 = (Ywy6z6 & Gxy6z6);
assign Gxy6z6 = (~(Wkd7z6[2] & Ddmhw6));
assign Ywy6z6 = (Oxy6z6 & Wxy6z6);
assign Wxy6z6 = (~(Xhd7z6[2] & Eu46z6));
assign Eu46z6 = (~(Jamnv6 | Ddmhw6));
assign Oxy6z6 = (~(Vnd7z6[2] & Jamnv6));
assign Qs46z6 = (~(Eyy6z6 & Au0ov6));
assign Au0ov6 = (Pcmhw6 & E2k6z6);
assign E2k6z6 = (!Qdcdt6);
assign Eyy6z6 = (~(Emoov6 | Mu46z6));
assign Mu46z6 = (~(Myy6z6 & Uyy6z6));
assign Uyy6z6 = (E31ov6 | Znnov6);
assign E31ov6 = (~(Czy6z6 | Geddt6));
assign Czy6z6 = (T8ddt6 | Nbddt6);
assign Myy6z6 = (Iooov6 & Qsoov6);
assign Qsoov6 = (Z8oov6 | Cgc7z6[2]);
assign Z8oov6 = (!Oznov6);
assign Oznov6 = (I51ov6 & Cgc7z6[1]);
assign Iooov6 = (~(Qmnov6 & P1piw6));
assign Qmnov6 = (I51ov6 & Cgc7z6[2]);
assign Emoov6 = (~(Bwnov6 & Nx0ov6));
assign Nx0ov6 = (!N9oov6);
assign N9oov6 = (E6piw6 & V4jhw6);
assign E6piw6 = (!W51ov6);
assign W51ov6 = (~(Kzy6z6 & Cgc7z6[0]));
assign Bwnov6 = (R537x6 & X6xnv6);
assign R537x6 = (!Ipnov6);
assign Ipnov6 = (K3k6z6 & V4jhw6);
assign V4jhw6 = (!Cgc7z6[3]);
assign K3k6z6 = (B51ov6 & O4jhw6);
assign B51ov6 = (Cgc7z6[1] & A4jhw6);
assign Kvy6z6 = (Szy6z6 & A0z6z6);
assign A0z6z6 = (~(Qdcdt6 & E3c7z6[2]));
assign Szy6z6 = (I0z6z6 & Q0z6z6);
assign Q0z6z6 = (~(Pic7z6[2] & Ir0ov6));
assign I0z6z6 = (~(Znnov6 & P2j7z6[0]));
assign Znnov6 = (!X6xnv6);
assign HADDRD[9] = (~(Y0z6z6 & G1z6z6));
assign G1z6z6 = (~(Onret6 & Jn1ov6));
assign Y0z6z6 = (O1z6z6 & W1z6z6);
assign W1z6z6 = (~(Fvb7z6[9] & Vm1ov6));
assign O1z6z6 = (~(Cmm7z6[9] & Hm1ov6));
assign HADDRD[8] = (~(E2z6z6 & M2z6z6));
assign M2z6z6 = (~(Ppret6 & Jn1ov6));
assign E2z6z6 = (U2z6z6 & C3z6z6);
assign C3z6z6 = (~(Fvb7z6[8] & Vm1ov6));
assign U2z6z6 = (~(Cmm7z6[8] & Hm1ov6));
assign HADDRD[7] = (~(K3z6z6 & S3z6z6));
assign S3z6z6 = (~(Qrret6 & Jn1ov6));
assign K3z6z6 = (A4z6z6 & I4z6z6);
assign I4z6z6 = (~(Fvb7z6[7] & Vm1ov6));
assign A4z6z6 = (~(Cmm7z6[7] & Hm1ov6));
assign HADDRD[6] = (~(Q4z6z6 & Y4z6z6));
assign Y4z6z6 = (~(Rtret6 & Jn1ov6));
assign Q4z6z6 = (G5z6z6 & O5z6z6);
assign O5z6z6 = (~(Fvb7z6[6] & Vm1ov6));
assign G5z6z6 = (~(Cmm7z6[6] & Hm1ov6));
assign HADDRD[5] = (~(W5z6z6 & E6z6z6));
assign E6z6z6 = (~(Svret6 & Jn1ov6));
assign W5z6z6 = (M6z6z6 & U6z6z6);
assign U6z6z6 = (~(Fvb7z6[5] & Vm1ov6));
assign M6z6z6 = (~(Cmm7z6[5] & Hm1ov6));
assign HADDRD[4] = (~(C7z6z6 & K7z6z6));
assign K7z6z6 = (~(Txret6 & Jn1ov6));
assign C7z6z6 = (S7z6z6 & A8z6z6);
assign A8z6z6 = (~(Fvb7z6[4] & Vm1ov6));
assign S7z6z6 = (~(Cmm7z6[4] & Hm1ov6));
assign HADDRD[3] = (~(I8z6z6 & Q8z6z6));
assign Q8z6z6 = (~(Uzret6 & Jn1ov6));
assign I8z6z6 = (Y8z6z6 & G9z6z6);
assign G9z6z6 = (~(Fvb7z6[3] & Vm1ov6));
assign Y8z6z6 = (~(Cmm7z6[3] & Hm1ov6));
assign HADDRD[2] = (~(O9z6z6 & W9z6z6));
assign W9z6z6 = (~(V1set6 & Jn1ov6));
assign O9z6z6 = (Eaz6z6 & Maz6z6);
assign Maz6z6 = (~(Yefnv6 & Hm1ov6));
assign Yefnv6 = (!I1c8x6);
assign I1c8x6 = (~(Xz7et6 & U28et6));
assign Eaz6z6 = (~(Fvb7z6[2] & Vm1ov6));
assign HADDRD[28] = (~(Uaz6z6 & Cbz6z6));
assign Cbz6z6 = (~(Vkqet6 & Jn1ov6));
assign Uaz6z6 = (Kbz6z6 & Sbz6z6);
assign Sbz6z6 = (~(Fvb7z6[28] & Vm1ov6));
assign Kbz6z6 = (~(Cmm7z6[28] & Hm1ov6));
assign HADDRD[27] = (~(Acz6z6 & Icz6z6));
assign Icz6z6 = (~(Wmqet6 & Jn1ov6));
assign Acz6z6 = (Qcz6z6 & Ycz6z6);
assign Ycz6z6 = (~(Fvb7z6[27] & Vm1ov6));
assign Qcz6z6 = (~(Cmm7z6[27] & Hm1ov6));
assign HADDRD[26] = (~(Gdz6z6 & Odz6z6));
assign Odz6z6 = (~(Xoqet6 & Jn1ov6));
assign Gdz6z6 = (Wdz6z6 & Eez6z6);
assign Eez6z6 = (~(Fvb7z6[26] & Vm1ov6));
assign Wdz6z6 = (~(Cmm7z6[26] & Hm1ov6));
assign HADDRD[25] = (~(Mez6z6 & Uez6z6));
assign Uez6z6 = (~(Yqqet6 & Jn1ov6));
assign Mez6z6 = (Cfz6z6 & Kfz6z6);
assign Kfz6z6 = (~(Vm1ov6 & Fvb7z6[25]));
assign Cfz6z6 = (~(Hm1ov6 & Cmm7z6[25]));
assign HADDRD[24] = (~(Sfz6z6 & Agz6z6));
assign Agz6z6 = (~(Zsqet6 & Jn1ov6));
assign Sfz6z6 = (Igz6z6 & Qgz6z6);
assign Qgz6z6 = (~(Fvb7z6[24] & Vm1ov6));
assign Igz6z6 = (~(Cmm7z6[24] & Hm1ov6));
assign HADDRD[23] = (~(Ygz6z6 & Ghz6z6));
assign Ghz6z6 = (~(Avqet6 & Jn1ov6));
assign Ygz6z6 = (Ohz6z6 & Whz6z6);
assign Whz6z6 = (~(Fvb7z6[23] & Vm1ov6));
assign Ohz6z6 = (~(Cmm7z6[23] & Hm1ov6));
assign HADDRD[22] = (~(Eiz6z6 & Miz6z6));
assign Miz6z6 = (~(Bxqet6 & Jn1ov6));
assign Eiz6z6 = (Uiz6z6 & Cjz6z6);
assign Cjz6z6 = (~(Fvb7z6[22] & Vm1ov6));
assign Uiz6z6 = (~(Cmm7z6[22] & Hm1ov6));
assign HADDRD[21] = (~(Kjz6z6 & Sjz6z6));
assign Sjz6z6 = (~(Czqet6 & Jn1ov6));
assign Kjz6z6 = (Akz6z6 & Ikz6z6);
assign Ikz6z6 = (~(Fvb7z6[21] & Vm1ov6));
assign Akz6z6 = (~(Cmm7z6[21] & Hm1ov6));
assign HADDRD[20] = (~(Qkz6z6 & Ykz6z6));
assign Ykz6z6 = (~(D1ret6 & Jn1ov6));
assign Qkz6z6 = (Glz6z6 & Olz6z6);
assign Olz6z6 = (~(Fvb7z6[20] & Vm1ov6));
assign Glz6z6 = (~(Cmm7z6[20] & Hm1ov6));
assign HADDRD[1] = (~(Wlz6z6 & Emz6z6));
assign Emz6z6 = (~(W3set6 & Jn1ov6));
assign Wlz6z6 = (Mmz6z6 & Umz6z6);
assign Umz6z6 = (~(Vm1ov6 & Stpnv6));
assign Mmz6z6 = (~(Hm1ov6 & Cmm7z6[1]));
assign HADDRD[19] = (~(Cnz6z6 & Knz6z6));
assign Knz6z6 = (~(E3ret6 & Jn1ov6));
assign Cnz6z6 = (Snz6z6 & Aoz6z6);
assign Aoz6z6 = (~(Fvb7z6[19] & Vm1ov6));
assign Snz6z6 = (~(Cmm7z6[19] & Hm1ov6));
assign HADDRD[18] = (~(Ioz6z6 & Qoz6z6));
assign Qoz6z6 = (~(F5ret6 & Jn1ov6));
assign Ioz6z6 = (Yoz6z6 & Gpz6z6);
assign Gpz6z6 = (~(Fvb7z6[18] & Vm1ov6));
assign Yoz6z6 = (~(Cmm7z6[18] & Hm1ov6));
assign HADDRD[17] = (~(Opz6z6 & Wpz6z6));
assign Wpz6z6 = (~(G7ret6 & Jn1ov6));
assign Opz6z6 = (Eqz6z6 & Mqz6z6);
assign Mqz6z6 = (~(Fvb7z6[17] & Vm1ov6));
assign Eqz6z6 = (~(Cmm7z6[17] & Hm1ov6));
assign HADDRD[16] = (~(Uqz6z6 & Crz6z6));
assign Crz6z6 = (~(H9ret6 & Jn1ov6));
assign Uqz6z6 = (Krz6z6 & Srz6z6);
assign Srz6z6 = (~(Fvb7z6[16] & Vm1ov6));
assign Krz6z6 = (~(Cmm7z6[16] & Hm1ov6));
assign HADDRD[15] = (~(Asz6z6 & Isz6z6));
assign Isz6z6 = (~(Ibret6 & Jn1ov6));
assign Asz6z6 = (Qsz6z6 & Ysz6z6);
assign Ysz6z6 = (~(Fvb7z6[15] & Vm1ov6));
assign Qsz6z6 = (~(Cmm7z6[15] & Hm1ov6));
assign HADDRD[14] = (~(Gtz6z6 & Otz6z6));
assign Otz6z6 = (~(Jdret6 & Jn1ov6));
assign Gtz6z6 = (Wtz6z6 & Euz6z6);
assign Euz6z6 = (~(Fvb7z6[14] & Vm1ov6));
assign Wtz6z6 = (~(Cmm7z6[14] & Hm1ov6));
assign HADDRD[13] = (~(Muz6z6 & Uuz6z6));
assign Uuz6z6 = (~(Kfret6 & Jn1ov6));
assign Muz6z6 = (Cvz6z6 & Kvz6z6);
assign Kvz6z6 = (~(Fvb7z6[13] & Vm1ov6));
assign Cvz6z6 = (~(Cmm7z6[13] & Hm1ov6));
assign HADDRD[12] = (~(Svz6z6 & Awz6z6));
assign Awz6z6 = (~(Lhret6 & Jn1ov6));
assign Svz6z6 = (Iwz6z6 & Qwz6z6);
assign Qwz6z6 = (~(Fvb7z6[12] & Vm1ov6));
assign Iwz6z6 = (~(Cmm7z6[12] & Hm1ov6));
assign HADDRD[11] = (~(Ywz6z6 & Gxz6z6));
assign Gxz6z6 = (~(Mjret6 & Jn1ov6));
assign Ywz6z6 = (Oxz6z6 & Wxz6z6);
assign Wxz6z6 = (~(Fvb7z6[11] & Vm1ov6));
assign Oxz6z6 = (~(Cmm7z6[11] & Hm1ov6));
assign HADDRD[10] = (~(Eyz6z6 & Myz6z6));
assign Myz6z6 = (~(Nlret6 & Jn1ov6));
assign Eyz6z6 = (Uyz6z6 & Czz6z6);
assign Czz6z6 = (~(Fvb7z6[10] & Vm1ov6));
assign Uyz6z6 = (~(Cmm7z6[10] & Hm1ov6));
assign HADDRD[0] = (~(Kzz6z6 & Szz6z6));
assign Szz6z6 = (~(X5set6 & Jn1ov6));
assign Kzz6z6 = (A007z6 & I007z6);
assign I007z6 = (~(Vm1ov6 & Mbqnv6));
assign Vm1ov6 = (!V4myx6);
assign V4myx6 = (~(Q007z6 & Y007z6));
assign Y007z6 = (G107z6 & O107z6);
assign O107z6 = (~(Jn1ov6 | U4zet6));
assign G107z6 = (W107z6 & E207z6);
assign Q007z6 = (Yx1iw6 & M207z6);
assign M207z6 = (U207z6 & C307z6);
assign U207z6 = (~(K307z6 & S307z6));
assign S307z6 = (~(A407z6 & I407z6));
assign I407z6 = (~(Aoyiy6 | Wmoet6));
assign Aoyiy6 = (Ewyet6 & Kb0jy6);
assign Kb0jy6 = (~(Xvgxx6 | Benyx6));
assign A407z6 = (Emy6z6 & Q407z6);
assign Q407z6 = (~(Ewyet6 & Qln7z6[1]));
assign Emy6z6 = (~(Ekoet6 | Y407z6));
assign Y407z6 = (Q086z6 & G507z6);
assign G507z6 = (~(O507z6 & Ikw6z6));
assign Ikw6z6 = (U6y5z6 & Tbqnv6);
assign U6y5z6 = (!Xnnet6);
assign O507z6 = (W507z6 & Ag0jy6);
assign Ag0jy6 = (~(E607z6 & P6u6x6));
assign P6u6x6 = (M607z6 & A9gxx6);
assign A9gxx6 = (Benyx6 & Rxixx6);
assign Benyx6 = (!Znn7z6[0]);
assign M607z6 = (~(Eq0jy6 | U607z6));
assign Eq0jy6 = (!Qakiw6);
assign Qakiw6 = (Vugxx6 & Xvgxx6);
assign E607z6 = (C707z6 & Knh7v6);
assign C707z6 = (Dkm7z6[0] | Dkm7z6[1]);
assign W507z6 = (I086z6 | U607z6);
assign I086z6 = (~(Wcmov6 & K707z6));
assign Yx1iw6 = (~(K7giy6 | Kjy6z6));
assign Kjy6z6 = (S707z6 | Fvb7z6[29]);
assign S707z6 = (Fvb7z6[30] | Fvb7z6[31]);
assign K7giy6 = (!K4bdt6);
assign A007z6 = (~(Hm1ov6 & Cmm7z6[0]));
assign GATEHCLK = (A807z6 & I807z6);
assign I807z6 = (~(ISOLATEn & Bq5yx6));
assign Bq5yx6 = (!Bnhiw6);
assign Bnhiw6 = (SLEEPING | Gwj8v6);
assign SLEEPING = (Q807z6 & Y807z6);
assign Q807z6 = (~(Crcdt6 | Ztcdt6));
assign A807z6 = (T1zhw6 & D9h7v6);
assign T1zhw6 = (!Kr97z6);
assign EXREQS = (~(G907z6 & O907z6));
assign O907z6 = (~(J0jxx6 & W907z6));
assign W907z6 = (~(Ea07z6 & Ma07z6));
assign Ma07z6 = (~(Ua07z6 & Ozadt6));
assign Ea07z6 = (~(H7nyx6 & E1uet6));
assign H7nyx6 = (!Luixx6);
assign Luixx6 = (~(Q0j6z6 & Qo8iy6));
assign Q0j6z6 = (Znn7z6[0] & Rxixx6);
assign G907z6 = (~(Cyphw6 & Rj9ov6));
assign Rj9ov6 = (~(Kfy6z6 | J0jxx6));
assign J0jxx6 = (!Uaonv6);
assign Uaonv6 = (~(Cb07z6 & U2v5z6));
assign U2v5z6 = (Kb07z6 & Qln7z6[1]);
assign Kb07z6 = (Znn7z6[0] & Sb07z6);
assign Sb07z6 = (~(Ac07z6 & Cakiw6));
assign Ac07z6 = (Rxixx6 ? Xvgxx6 : Znn7z6[2]);
assign Cb07z6 = (Ic07z6 & Qky6z6);
assign Ic07z6 = (~(Kyn7z6[0] & Gazet6));
assign Kfy6z6 = (~(Sjwiy6 & Wcmov6));
assign Sjwiy6 = (Qc07z6 & Yc07z6);
assign Yc07z6 = (Gd07z6 & Lxjiw6);
assign Lxjiw6 = (Lgonv6 & Szphw6);
assign Szphw6 = (!Ysdiw6);
assign Lgonv6 = (~(Od07z6 & Wd07z6));
assign Wd07z6 = (Ee07z6 & Me07z6);
assign Me07z6 = (Ue07z6 & V0hnv6);
assign Ue07z6 = (O0hnv6 & H0hnv6);
assign Ee07z6 = (Cf07z6 & Q1hnv6);
assign Q1hnv6 = (!Cmm7z6[23]);
assign Cf07z6 = (J1hnv6 & C1hnv6);
assign C1hnv6 = (!Cmm7z6[25]);
assign J1hnv6 = (!Cmm7z6[24]);
assign Od07z6 = (Kf07z6 & Sf07z6);
assign Sf07z6 = (Ag07z6 & L2hnv6);
assign L2hnv6 = (!Cmm7z6[20]);
assign Ag07z6 = (E2hnv6 & X1hnv6);
assign X1hnv6 = (!Cmm7z6[22]);
assign E2hnv6 = (!Cmm7z6[21]);
assign Kf07z6 = (~(Rygnv6 | Ig07z6));
assign Gd07z6 = (Dhnyx6 & Qky6z6);
assign Dhnyx6 = (~(Qg07z6 & Qo8iy6));
assign Qo8iy6 = (~(Vugxx6 | Xvgxx6));
assign Qg07z6 = (Znn7z6[1] & Znn7z6[0]);
assign Qc07z6 = (Yg07z6 & Cryiy6);
assign Cryiy6 = (Y497z6 & Gh07z6);
assign Gh07z6 = (W186z6 | Tbqnv6);
assign Tbqnv6 = (!Styet6);
assign W186z6 = (!Qln7z6[0]);
assign Yg07z6 = (Oh07z6 & Wh07z6);
assign Wh07z6 = (~(Kyn7z6[2] & Gazet6));
assign EXREQD = (Cyphw6 & Hm1ov6);
assign Hm1ov6 = (!Jfonv6);
assign Jfonv6 = (C307z6 | Jn1ov6);
assign Jn1ov6 = (!Ibonv6);
assign Ibonv6 = (~(Ei07z6 & Mi07z6));
assign Mi07z6 = (E207z6 & K307z6);
assign E207z6 = (~(Ysn7z6[0] & N7zet6));
assign Ei07z6 = (Qln7z6[0] & Djonv6);
assign Djonv6 = (Ozixx6 & Znn7z6[0]);
assign Ozixx6 = (~(Xvgxx6 | Znn7z6[2]));
assign C307z6 = (~(Wcmov6 & Whwiy6));
assign Whwiy6 = (Ui07z6 & Cj07z6);
assign Cj07z6 = (Kj07z6 & Sj07z6);
assign Sj07z6 = (~(Qboet6 | U4zet6));
assign Kj07z6 = (Uqyiy6 & K307z6);
assign Uqyiy6 = (~(Qln7z6[1] & Styet6));
assign Ui07z6 = (Ak07z6 & Ysdiw6);
assign Ysdiw6 = (Ohm6z6 & Rygnv6);
assign Ak07z6 = (Oh07z6 & W107z6);
assign W107z6 = (~(Ysn7z6[2] & N7zet6));
assign Oh07z6 = (Ik07z6 & Qk07z6);
assign Qk07z6 = (~(Bzjiw6 | U8oet6));
assign Bzjiw6 = (Yk07z6 & Y0m6z6);
assign Y0m6z6 = (Cakiw6 & Gl07z6);
assign Gl07z6 = (~(Rxixx6 & Xvgxx6));
assign Rxixx6 = (!Znn7z6[1]);
assign Cakiw6 = (Vugxx6 | Znn7z6[3]);
assign Vugxx6 = (!Znn7z6[2]);
assign Yk07z6 = (Styet6 & Znn7z6[0]);
assign Ik07z6 = (Kryiy6 & Ol07z6);
assign Ol07z6 = (~(K707z6 & Wl07z6));
assign Wl07z6 = (Em07z6 | U607z6);
assign U607z6 = (Mm07z6 & Q086z6);
assign Q086z6 = (~(Go9ov6 & E2ziy6));
assign E2ziy6 = (~(Um07z6 & Cn07z6));
assign Cn07z6 = (~(Kn07z6 | Fvb7z6[27]));
assign Kn07z6 = (Fvb7z6[28] | Fvb7z6[31]);
assign Um07z6 = (Sn07z6 & Fvb7z6[25]);
assign Sn07z6 = (Ao07z6 & Ghy6z6);
assign Ghy6z6 = (!Fvb7z6[26]);
assign Ao07z6 = (Fvb7z6[30] ^ Fvb7z6[29]);
assign Go9ov6 = (Jvdiw6 & Sbm6z6);
assign Sbm6z6 = (!Zwdiw6);
assign Zwdiw6 = (~(Io07z6 & Qo07z6));
assign Qo07z6 = (~(Hub7z6[0] & Mbqnv6));
assign Io07z6 = (~(Yo07z6 & Stpnv6));
assign Jvdiw6 = (~(Yo07z6 | Gp07z6));
assign Gp07z6 = (!Rzdiw6);
assign Rzdiw6 = (~(Op07z6 & Hub7z6[1]));
assign Op07z6 = (Stpnv6 & Wp07z6);
assign Stpnv6 = (~(Xie7x6 | A6wnv6));
assign Xie7x6 = (!Ugo7z6[1]);
assign Yo07z6 = (Mbqnv6 & Hub7z6[1]);
assign Mbqnv6 = (!Wp07z6);
assign Wp07z6 = (Qie7x6 | A6wnv6);
assign A6wnv6 = (~(Ejo7z6[1] & C7wnv6));
assign C7wnv6 = (!Ejo7z6[0]);
assign Qie7x6 = (!Ugo7z6[0]);
assign Mm07z6 = (~(Qky6z6 & K307z6));
assign K307z6 = (~(N7zet6 & Ysn7z6[1]));
assign Qky6z6 = (~(Gazet6 & Kyn7z6[1]));
assign Em07z6 = (Xnnet6 | Ewyet6);
assign K707z6 = (~(Zblov6 & Sgonv6));
assign Sgonv6 = (~(Eq07z6 & Mq07z6));
assign Mq07z6 = (Uq07z6 & Cr07z6);
assign Cr07z6 = (H0hnv6 & Rygnv6);
assign Rygnv6 = (!Cmm7z6[31]);
assign H0hnv6 = (!Cmm7z6[28]);
assign Uq07z6 = (V0hnv6 & O0hnv6);
assign O0hnv6 = (!Cmm7z6[27]);
assign V0hnv6 = (!Cmm7z6[26]);
assign Eq07z6 = (Kr07z6 & Cmm7z6[25]);
assign Kr07z6 = (Ig07z6 & Iom6z6);
assign Iom6z6 = (!Ohm6z6);
assign Ohm6z6 = (A0hnv6 & Yygnv6);
assign Yygnv6 = (!Cmm7z6[30]);
assign A0hnv6 = (!Cmm7z6[29]);
assign Ig07z6 = (~(Cmm7z6[30] & Cmm7z6[29]));
assign Zblov6 = (Srhiy6 & Nxdiw6);
assign Nxdiw6 = (~(Cmm7z6[0] & Sr07z6));
assign Sr07z6 = (~(Ta4iw6 & As07z6));
assign Ta4iw6 = (~(I0c7z6[0] & Is07z6));
assign Srhiy6 = (!Qvdiw6);
assign Qvdiw6 = (~(As07z6 & Qs07z6));
assign Qs07z6 = (~(Cmm7z6[0] & Anehw6));
assign As07z6 = (!Mam6z6);
assign Mam6z6 = (Cmm7z6[1] & Anehw6);
assign Anehw6 = (~(Ys07z6 & Gt07z6));
assign Gt07z6 = (Ot07z6 & Wt07z6);
assign Wt07z6 = (Eu07z6 & Kfoiy6);
assign Kfoiy6 = (~(Beyxx6 & Dwb7z6[1]));
assign Eu07z6 = (Srknv6 & Z2yxx6);
assign Z2yxx6 = (!Uakiy6);
assign Srknv6 = (!Hulov6);
assign Ot07z6 = (Cfv6z6 & Vcyxx6);
assign Cfv6z6 = (~(Mu07z6 & Ytlnv6));
assign Mu07z6 = (Kioov6 & Sna7x6);
assign Ys07z6 = (Uu07z6 & Cv07z6);
assign Cv07z6 = (Kv07z6 & Inphw6);
assign Inphw6 = (~(Sv07z6 & Vqihw6));
assign Sv07z6 = (Dwb7z6[4] & Dwb7z6[2]);
assign Kv07z6 = (Aw07z6 & Iw07z6);
assign Iw07z6 = (~(Qw07z6 & Eekiy6));
assign Qw07z6 = (Gonov6 & Dwb7z6[2]);
assign Aw07z6 = (~(I0c7z6[1] & Is07z6));
assign Is07z6 = (~(Ygv6z6 & Yw07z6));
assign Yw07z6 = (~(Gx07z6 & Doihw6));
assign Gx07z6 = (Ox07z6 & Zna7x6);
assign Ox07z6 = (Uvvnv6 ^ Bwvnv6);
assign Ygv6z6 = (Oxpiy6 & Wx07z6);
assign Wx07z6 = (~(S2a7x6 & C7jxx6));
assign Oxpiy6 = (~(Ey07z6 & Ywaov6));
assign Ey07z6 = (Fulnv6 & C7jxx6);
assign Uu07z6 = (My07z6 & Kfv6z6);
assign Kfv6z6 = (~(G5kiy6 & Luvnv6));
assign My07z6 = (~(Tiphw6 & Mpihw6));
assign Tiphw6 = (~(Gvvnv6 | Uvvnv6));
assign Kryiy6 = (~(Ua07z6 | Hryet6));
assign Ua07z6 = (!Lblov6);
assign Lblov6 = (Jinyx6 | Znn7z6[2]);
assign Jinyx6 = (~(Uy07z6 & Znn7z6[1]));
assign Uy07z6 = (Znn7z6[0] & Xvgxx6);
assign Xvgxx6 = (!Znn7z6[3]);
assign Wcmov6 = (~(Nsr7x6 | K6adt6));
assign Nsr7x6 = (!Vb4iw6);
assign Vb4iw6 = (~(Cz07z6 & Kz07z6));
assign Kz07z6 = (Sz07z6 & A017z6);
assign A017z6 = (Vcyxx6 & Fsxxx6);
assign Fsxxx6 = (!H7wxx6);
assign H7wxx6 = (Fulnv6 & G5kiy6);
assign Vcyxx6 = (~(I017z6 & K3jnv6));
assign I017z6 = (~(Xxknv6 | Tnzdt6));
assign Xxknv6 = (~(Ywaov6 & Kioov6));
assign Sz07z6 = (Iwjiy6 & Q017z6);
assign Q017z6 = (~(Y017z6 & Eekiy6));
assign Eekiy6 = (Bhoov6 & Fulnv6);
assign Y017z6 = (Dwb7z6[2] & Rgo7v6);
assign Rgo7v6 = (~(Venov6 | Aiadt6));
assign Venov6 = (!Gonov6);
assign Gonov6 = (~(Tnzdt6 | Kkadt6));
assign Iwjiy6 = (Eminv6 | Cubdt6);
assign Eminv6 = (~(U6hiy6 & Kioov6));
assign Cz07z6 = (G117z6 & O117z6);
assign O117z6 = (W117z6 & E217z6);
assign E217z6 = (~(M217z6 & Lxydt6));
assign M217z6 = (~(U217z6 & C317z6));
assign C317z6 = (K317z6 & S317z6);
assign S317z6 = (~(A417z6 & Vglhw6));
assign Vglhw6 = (~(Iqmov6 & Mulnv6));
assign Mulnv6 = (!Pi9ov6);
assign Pi9ov6 = (Ltvxx6 & Dwb7z6[1]);
assign Iqmov6 = (Gha7x6 | Mpihw6);
assign Mpihw6 = (!Fulnv6);
assign Gha7x6 = (!Rb9iw6);
assign Rb9iw6 = (Ywaov6 & Ytlnv6);
assign Ywaov6 = (~(Gvvnv6 | Sna7x6));
assign A417z6 = (~(I417z6 & Bi9ov6));
assign I417z6 = (Ii9ov6 & F5jxx6);
assign F5jxx6 = (!S7xdt6);
assign Ii9ov6 = (!Zzihw6);
assign Zzihw6 = (Ecc7z6[6] & Pbadt6);
assign K317z6 = (~(Dihhw6 | Hulov6));
assign Dihhw6 = (Uakiy6 & Fxaov6);
assign U217z6 = (P3yxx6 & Q417z6);
assign Q417z6 = (~(Ruxxx6 & Kioov6));
assign P3yxx6 = (Ojphw6 & Rja7x6);
assign Rja7x6 = (~(Cwlnv6 | U2wnv6));
assign U2wnv6 = (Sv97x6 & Dwb7z6[2]);
assign Sv97x6 = (!Tulnv6);
assign Tulnv6 = (~(Y417z6 & Doihw6));
assign Y417z6 = (Fxaov6 & Uvvnv6);
assign Cwlnv6 = (S2a7x6 & Xfa7x6);
assign S2a7x6 = (~(Xvxxx6 | Euvnv6));
assign Xvxxx6 = (!Vqihw6);
assign Ojphw6 = (L0bov6 & Eyi6z6);
assign Eyi6z6 = (~(Ltvxx6 & Kioov6));
assign Ltvxx6 = (Ytlnv6 & Doihw6);
assign L0bov6 = (J1a7x6 | Dwb7z6[5]);
assign J1a7x6 = (~(G517z6 & Dwb7z6[4]));
assign G517z6 = (Kioov6 & Nvvnv6);
assign W117z6 = (~(O517z6 & M43et6));
assign O517z6 = (K73et6 & Hulov6);
assign Hulov6 = (Ggoov6 & Fulnv6);
assign Ggoov6 = (Bhoov6 & Ytlnv6);
assign Bhoov6 = (~(Sna7x6 | Dwb7z6[4]));
assign G117z6 = (A8k6z6 & G9k6z6);
assign G9k6z6 = (T1yxx6 | Iga7z6);
assign T1yxx6 = (~(Wxi6z6 | Rioov6));
assign Rioov6 = (!Yihhw6);
assign Yihhw6 = (Ajphw6 | Dwb7z6[3]);
assign Ajphw6 = (~(Fxaov6 & Beyxx6));
assign Beyxx6 = (~(Pnxxx6 | Dwb7z6[2]));
assign Wxi6z6 = (W517z6 & Vqihw6);
assign W517z6 = (Dioov6 & Dwb7z6[4]);
assign A8k6z6 = (E617z6 & M617z6);
assign M617z6 = (~(U617z6 & Bfo7v6));
assign U617z6 = (~(M6hiy6 & Qsaov6));
assign Qsaov6 = (~(U6hiy6 & Vqihw6));
assign U6hiy6 = (~(Mmriy6 | Pnxxx6));
assign Pnxxx6 = (!Lpwxx6);
assign Lpwxx6 = (Dwb7z6[4] & Sna7x6);
assign Mmriy6 = (!Ytlnv6);
assign Ytlnv6 = (C7jxx6 & Uvvnv6);
assign M6hiy6 = (~(Uakiy6 & Fulnv6));
assign E617z6 = (C717z6 & K717z6);
assign K717z6 = (~(S717z6 & Sj77z6));
assign S717z6 = (~(Vovxx6 | Twphw6));
assign Twphw6 = (!Clhhw6);
assign Clhhw6 = (Ruxxx6 & Fulnv6);
assign Fulnv6 = (Luvnv6 & Bwvnv6);
assign Ruxxx6 = (~(Euvnv6 | Isjiy6));
assign Euvnv6 = (!Doihw6);
assign Vovxx6 = (!Lsphw6);
assign Lsphw6 = (Lxydt6 & Hjihw6);
assign Hjihw6 = (!Wfxdt6);
assign C717z6 = (~(A817z6 & Lxydt6));
assign Lxydt6 = (Bfo7v6 & Qg2nv6);
assign Bfo7v6 = (!Iga7z6);
assign Iga7z6 = (~(I817z6 & Tr8iw6));
assign Tr8iw6 = (~(Ez2et6 & I2jnv6));
assign I2jnv6 = (!U1jnv6);
assign U1jnv6 = (~(Q817z6 & Y817z6));
assign Y817z6 = (G917z6 | Tfh7z6[1]);
assign G917z6 = (Tfh7z6[0] & Cmm7z6[0]);
assign Q817z6 = (~(D94iw6 & Xc4iw6));
assign Xc4iw6 = (!Cmm7z6[1]);
assign D94iw6 = (!Cmm7z6[0]);
assign I817z6 = (Ijmov6 & Ftlov6);
assign Ftlov6 = (!M43et6);
assign Ijmov6 = (!Uebdt6);
assign A817z6 = (~(O917z6 & W917z6));
assign W917z6 = (Ea17z6 & X3yxx6);
assign X3yxx6 = (~(Fxaov6 & G5kiy6));
assign G5kiy6 = (~(Sna7x6 | Isjiy6));
assign Isjiy6 = (!Nvvnv6);
assign Ea17z6 = (~(B2yxx6 | Ot97x6));
assign Ot97x6 = (Vqihw6 & Mahiy6);
assign Mahiy6 = (Doihw6 & Dioov6);
assign Dioov6 = (Dwb7z6[2] & Uvvnv6);
assign Uvvnv6 = (!Dwb7z6[3]);
assign Doihw6 = (Gvvnv6 & Sna7x6);
assign Sna7x6 = (!Dwb7z6[5]);
assign Gvvnv6 = (!Dwb7z6[4]);
assign B2yxx6 = (Dophw6 & Fxaov6);
assign Fxaov6 = (Dwb7z6[1] & Luvnv6);
assign Luvnv6 = (!Dwb7z6[0]);
assign Dophw6 = (Dwb7z6[4] & Nvvnv6);
assign Nvvnv6 = (Dwb7z6[3] & Dwb7z6[2]);
assign O917z6 = (Ma17z6 & Ua17z6);
assign Ua17z6 = (~(Rmwxx6 & Dwb7z6[4]));
assign Rmwxx6 = (~(Zna7x6 | Bqvxx6));
assign Bqvxx6 = (!Kioov6);
assign Kioov6 = (Dwb7z6[0] & Bwvnv6);
assign Bwvnv6 = (!Dwb7z6[1]);
assign Zna7x6 = (!Xfa7x6);
assign Ma17z6 = (~(Uakiy6 & Vqihw6));
assign Vqihw6 = (Dwb7z6[1] & Dwb7z6[0]);
assign Uakiy6 = (Xfa7x6 & Dwb7z6[4]);
assign Xfa7x6 = (Dwb7z6[3] & C7jxx6);
assign C7jxx6 = (!Dwb7z6[2]);
assign Cyphw6 = (Cb17z6 & Tlmov6);
assign Tlmov6 = (~(Oe2et6 | Ldbdt6));
assign Cb17z6 = (Bi9ov6 & Ldo7v6);
assign Bi9ov6 = (Ecc7z6[13] & Pbadt6);
assign ETMINTNUM[8] = (Glh7v6 & Nob7z6[8]);
assign ETMINTNUM[7] = (Glh7v6 & Nob7z6[7]);
assign ETMINTNUM[6] = (Glh7v6 ? Nob7z6[6] : P2j7z6[6]);
assign ETMINTNUM[5] = (Glh7v6 ? Nob7z6[5] : P2j7z6[5]);
assign ETMINTNUM[4] = (Glh7v6 ? Nob7z6[4] : P2j7z6[4]);
assign ETMINTNUM[3] = (Glh7v6 ? Nob7z6[3] : P2j7z6[3]);
assign ETMINTNUM[2] = (Glh7v6 ? Nob7z6[2] : P2j7z6[2]);
assign ETMINTNUM[1] = (Glh7v6 ? Nob7z6[1] : P2j7z6[1]);
assign ETMINTNUM[0] = (Glh7v6 ? Nob7z6[0] : P2j7z6[0]);
assign CURRPRI[7] = (~(Kb17z6 & Sb17z6));
assign Sb17z6 = (Ac17z6 & Ic17z6);
assign Ic17z6 = (~(Sz3jy6 & Qc17z6));
assign Qc17z6 = (~(Yc17z6 & Gd17z6));
assign Gd17z6 = (Od17z6 & Wd17z6);
assign Wd17z6 = (Ee17z6 & Me17z6);
assign Me17z6 = (~(Ao2jy6 & Gx08x6));
assign Gx08x6 = (Ppb7z6[7] | Jm98x6);
assign Jm98x6 = (!J92nv6);
assign Ee17z6 = (~(Ffj7z6[2] & Cshov6));
assign Od17z6 = (Ue17z6 & Cf17z6);
assign Cf17z6 = (~(Zdj7z6[2] & I2oiw6));
assign Ue17z6 = (~(Tcj7z6[2] & Rphov6));
assign Yc17z6 = (Kf17z6 & Sf17z6);
assign Sf17z6 = (Ag17z6 & Ig17z6);
assign Ig17z6 = (~(Gaj7z6[2] & Hzh7x6));
assign Ag17z6 = (~(Nbj7z6[2] & L1i7x6));
assign Kf17z6 = (Qg17z6 & Yg17z6);
assign Yg17z6 = (~(Z8j7z6[2] & P3i7x6));
assign Qg17z6 = (~(T7j7z6[2] & V6i7x6));
assign Ac17z6 = (Gh17z6 & Oh17z6);
assign Oh17z6 = (~(Wtgjy6 & Wh17z6));
assign Wh17z6 = (~(Ei17z6 & Mi17z6));
assign Mi17z6 = (Ui17z6 & Cj17z6);
assign Cj17z6 = (Kj17z6 & Sj17z6);
assign Sj17z6 = (Ak17z6 & Ik17z6);
assign Ik17z6 = (~(Lgj7z6[2] & Ao2jy6));
assign Ak17z6 = (~(Lgj7z6[5] & Nuniw6));
assign Kj17z6 = (Qk17z6 & Yk17z6);
assign Yk17z6 = (~(Lgj7z6[8] & Jfmiw6));
assign Qk17z6 = (~(Lgj7z6[11] & Cn2jy6));
assign Ui17z6 = (Gl17z6 & Ol17z6);
assign Ol17z6 = (Wl17z6 & Em17z6);
assign Em17z6 = (~(Lgj7z6[14] & Cshov6));
assign Wl17z6 = (~(Lgj7z6[17] & I2oiw6));
assign Gl17z6 = (Mm17z6 & Um17z6);
assign Um17z6 = (~(Lgj7z6[20] & Rphov6));
assign Mm17z6 = (~(Lgj7z6[23] & J6oiw6));
assign Ei17z6 = (Cn17z6 & Kn17z6);
assign Kn17z6 = (Sn17z6 & Ao17z6);
assign Ao17z6 = (Io17z6 & Qo17z6);
assign Qo17z6 = (~(Lgj7z6[26] & Uy2jy6));
assign Io17z6 = (~(Lgj7z6[29] & Mbj7x6));
assign Sn17z6 = (Yo17z6 & Gp17z6);
assign Gp17z6 = (~(Lgj7z6[32] & Nfj7x6));
assign Yo17z6 = (~(Lgj7z6[35] & Hzh7x6));
assign Cn17z6 = (Op17z6 & Wp17z6);
assign Wp17z6 = (Eq17z6 & Mq17z6);
assign Mq17z6 = (~(Lgj7z6[38] & L1i7x6));
assign Eq17z6 = (~(Lgj7z6[41] & Jrj7x6));
assign Op17z6 = (Uq17z6 & Cr17z6);
assign Cr17z6 = (~(Lgj7z6[44] & P3i7x6));
assign Uq17z6 = (~(Lgj7z6[47] & V6i7x6));
assign Gh17z6 = (~(Awcjy6 & Kr17z6));
assign Kr17z6 = (~(Sr17z6 & As17z6));
assign As17z6 = (Is17z6 & Qs17z6);
assign Qs17z6 = (Ys17z6 & Gt17z6);
assign Gt17z6 = (Ot17z6 & Wt17z6);
assign Wt17z6 = (~(Lgj7z6[50] & Ao2jy6));
assign Ot17z6 = (~(Lgj7z6[53] & Nuniw6));
assign Ys17z6 = (Eu17z6 & Mu17z6);
assign Mu17z6 = (~(Lgj7z6[56] & Jfmiw6));
assign Eu17z6 = (~(Lgj7z6[59] & Cn2jy6));
assign Is17z6 = (Uu17z6 & Cv17z6);
assign Cv17z6 = (Kv17z6 & Sv17z6);
assign Sv17z6 = (~(Cshov6 & Lgj7z6[62]));
assign Kv17z6 = (~(I2oiw6 & Lgj7z6[65]));
assign Uu17z6 = (Aw17z6 & Iw17z6);
assign Iw17z6 = (~(Lgj7z6[68] & Rphov6));
assign Aw17z6 = (~(J6oiw6 & Lgj7z6[71]));
assign Sr17z6 = (Qw17z6 & Yw17z6);
assign Yw17z6 = (Gx17z6 & Ox17z6);
assign Ox17z6 = (Wx17z6 & Ey17z6);
assign Ey17z6 = (~(Lgj7z6[74] & Uy2jy6));
assign Wx17z6 = (~(Lgj7z6[77] & Mbj7x6));
assign Gx17z6 = (My17z6 & Uy17z6);
assign Uy17z6 = (~(Lgj7z6[80] & Nfj7x6));
assign My17z6 = (~(Lgj7z6[83] & Hzh7x6));
assign Qw17z6 = (Cz17z6 & Kz17z6);
assign Kz17z6 = (Sz17z6 & A027z6);
assign A027z6 = (~(Lgj7z6[86] & L1i7x6));
assign Sz17z6 = (~(Jrj7x6 & Lgj7z6[89]));
assign Cz17z6 = (I027z6 & Q027z6);
assign Q027z6 = (~(Lgj7z6[92] & P3i7x6));
assign I027z6 = (~(Lgj7z6[95] & V6i7x6));
assign Kb17z6 = (Y027z6 & G127z6);
assign G127z6 = (~(Maajy6 & O127z6));
assign O127z6 = (~(W127z6 & E227z6));
assign E227z6 = (M227z6 & U227z6);
assign U227z6 = (C327z6 & K327z6);
assign K327z6 = (S327z6 & A427z6);
assign A427z6 = (~(Lgj7z6[98] & Ao2jy6));
assign S327z6 = (~(Lgj7z6[101] & Nuniw6));
assign C327z6 = (I427z6 & Q427z6);
assign Q427z6 = (~(Lgj7z6[104] & Jfmiw6));
assign I427z6 = (~(Lgj7z6[107] & Cn2jy6));
assign M227z6 = (Y427z6 & G527z6);
assign G527z6 = (O527z6 & W527z6);
assign W527z6 = (~(Lgj7z6[110] & Cshov6));
assign O527z6 = (~(Lgj7z6[113] & I2oiw6));
assign Y427z6 = (E627z6 & M627z6);
assign M627z6 = (~(Lgj7z6[116] & Rphov6));
assign E627z6 = (~(Lgj7z6[119] & J6oiw6));
assign W127z6 = (U627z6 & C727z6);
assign C727z6 = (K727z6 & S727z6);
assign S727z6 = (A827z6 & I827z6);
assign I827z6 = (~(Lgj7z6[122] & Uy2jy6));
assign A827z6 = (~(Lgj7z6[125] & Mbj7x6));
assign K727z6 = (Q827z6 & Y827z6);
assign Y827z6 = (~(Lgj7z6[128] & Nfj7x6));
assign Q827z6 = (~(Lgj7z6[131] & Hzh7x6));
assign U627z6 = (G927z6 & O927z6);
assign O927z6 = (W927z6 & Ea27z6);
assign Ea27z6 = (~(Lgj7z6[134] & L1i7x6));
assign W927z6 = (~(Lgj7z6[137] & Jrj7x6));
assign G927z6 = (Ma27z6 & Ua27z6);
assign Ua27z6 = (~(Lgj7z6[140] & P3i7x6));
assign Ma27z6 = (~(Lgj7z6[143] & V6i7x6));
assign Y027z6 = (~(A87jy6 & Cb27z6));
assign Cb27z6 = (~(Kb27z6 & Sb27z6));
assign Sb27z6 = (Ac27z6 & Ic27z6);
assign Ic27z6 = (Qc27z6 & Yc27z6);
assign Yc27z6 = (Gd27z6 & Od27z6);
assign Od27z6 = (~(Lgj7z6[146] & Ao2jy6));
assign Gd27z6 = (~(Lgj7z6[149] & Nuniw6));
assign Qc27z6 = (Wd27z6 & Ee27z6);
assign Ee27z6 = (~(Lgj7z6[152] & Jfmiw6));
assign Wd27z6 = (~(Lgj7z6[155] & Cn2jy6));
assign Ac27z6 = (Me27z6 & Ue27z6);
assign Ue27z6 = (Cf27z6 & Kf27z6);
assign Kf27z6 = (~(Lgj7z6[158] & Cshov6));
assign Cf27z6 = (~(Lgj7z6[161] & I2oiw6));
assign Me27z6 = (Sf27z6 & Ag27z6);
assign Ag27z6 = (~(Lgj7z6[164] & Rphov6));
assign Sf27z6 = (~(Lgj7z6[167] & J6oiw6));
assign Kb27z6 = (Ig27z6 & Qg27z6);
assign Qg27z6 = (Yg27z6 & Gh27z6);
assign Gh27z6 = (Oh27z6 & Wh27z6);
assign Wh27z6 = (~(Lgj7z6[170] & Uy2jy6));
assign Oh27z6 = (~(Lgj7z6[173] & Mbj7x6));
assign Yg27z6 = (Ei27z6 & Mi27z6);
assign Mi27z6 = (~(Lgj7z6[176] & Nfj7x6));
assign Ei27z6 = (~(Lgj7z6[179] & Hzh7x6));
assign Ig27z6 = (Ui27z6 & Cj27z6);
assign Cj27z6 = (Kj27z6 & Sj27z6);
assign Sj27z6 = (~(Lgj7z6[182] & L1i7x6));
assign Kj27z6 = (~(Lgj7z6[185] & Jrj7x6));
assign Ui27z6 = (Ak27z6 & Ik27z6);
assign Ik27z6 = (~(Lgj7z6[188] & P3i7x6));
assign Ak27z6 = (~(Lgj7z6[191] & V6i7x6));
assign CURRPRI[6] = (~(Qk27z6 & Yk27z6));
assign Yk27z6 = (Gl27z6 & Ol27z6);
assign Ol27z6 = (~(Sz3jy6 & Wl27z6));
assign Wl27z6 = (~(Em27z6 & Mm27z6));
assign Mm27z6 = (Um27z6 & Cn27z6);
assign Cn27z6 = (Kn27z6 & Sn27z6);
assign Sn27z6 = (Rqmiw6 | Xg18x6);
assign Xg18x6 = (I8oiy6 & J92nv6);
assign I8oiy6 = (!Ppb7z6[6]);
assign Kn27z6 = (~(Ffj7z6[1] & Cshov6));
assign Um27z6 = (Ao27z6 & Io27z6);
assign Io27z6 = (~(Zdj7z6[1] & I2oiw6));
assign Ao27z6 = (~(Tcj7z6[1] & Rphov6));
assign Em27z6 = (Qo27z6 & Yo27z6);
assign Yo27z6 = (Gp27z6 & Op27z6);
assign Op27z6 = (~(Gaj7z6[1] & Hzh7x6));
assign Gp27z6 = (~(Nbj7z6[1] & L1i7x6));
assign Qo27z6 = (Wp27z6 & Eq27z6);
assign Eq27z6 = (~(Z8j7z6[1] & P3i7x6));
assign Wp27z6 = (~(T7j7z6[1] & V6i7x6));
assign Gl27z6 = (Mq27z6 & Uq27z6);
assign Uq27z6 = (~(Wtgjy6 & Cr27z6));
assign Cr27z6 = (~(Kr27z6 & Sr27z6));
assign Sr27z6 = (As27z6 & Is27z6);
assign Is27z6 = (Qs27z6 & Ys27z6);
assign Ys27z6 = (Gt27z6 & Ot27z6);
assign Ot27z6 = (~(Lgj7z6[1] & Ao2jy6));
assign Gt27z6 = (~(Lgj7z6[4] & Nuniw6));
assign Qs27z6 = (Wt27z6 & Eu27z6);
assign Eu27z6 = (~(Lgj7z6[7] & Jfmiw6));
assign Wt27z6 = (~(Lgj7z6[10] & Cn2jy6));
assign As27z6 = (Mu27z6 & Uu27z6);
assign Uu27z6 = (Cv27z6 & Kv27z6);
assign Kv27z6 = (~(Lgj7z6[13] & Cshov6));
assign Cv27z6 = (~(Lgj7z6[16] & I2oiw6));
assign Mu27z6 = (Sv27z6 & Aw27z6);
assign Aw27z6 = (~(Lgj7z6[19] & Rphov6));
assign Sv27z6 = (~(Lgj7z6[22] & J6oiw6));
assign Kr27z6 = (Iw27z6 & Qw27z6);
assign Qw27z6 = (Yw27z6 & Gx27z6);
assign Gx27z6 = (Ox27z6 & Wx27z6);
assign Wx27z6 = (~(Lgj7z6[25] & Uy2jy6));
assign Ox27z6 = (~(Lgj7z6[28] & Mbj7x6));
assign Yw27z6 = (Ey27z6 & My27z6);
assign My27z6 = (~(Lgj7z6[31] & Nfj7x6));
assign Ey27z6 = (~(Lgj7z6[34] & Hzh7x6));
assign Iw27z6 = (Uy27z6 & Cz27z6);
assign Cz27z6 = (Kz27z6 & Sz27z6);
assign Sz27z6 = (~(Lgj7z6[37] & L1i7x6));
assign Kz27z6 = (~(Lgj7z6[40] & Jrj7x6));
assign Uy27z6 = (A037z6 & I037z6);
assign I037z6 = (~(Lgj7z6[43] & P3i7x6));
assign A037z6 = (~(Lgj7z6[46] & V6i7x6));
assign Mq27z6 = (~(Awcjy6 & Q037z6));
assign Q037z6 = (~(Y037z6 & G137z6));
assign G137z6 = (O137z6 & W137z6);
assign W137z6 = (E237z6 & M237z6);
assign M237z6 = (U237z6 & C337z6);
assign C337z6 = (~(Lgj7z6[49] & Ao2jy6));
assign U237z6 = (~(Lgj7z6[52] & Nuniw6));
assign E237z6 = (K337z6 & S337z6);
assign S337z6 = (~(Lgj7z6[55] & Jfmiw6));
assign K337z6 = (~(Lgj7z6[58] & Cn2jy6));
assign O137z6 = (A437z6 & I437z6);
assign I437z6 = (Q437z6 & Y437z6);
assign Y437z6 = (~(Cshov6 & Lgj7z6[61]));
assign Q437z6 = (~(I2oiw6 & Lgj7z6[64]));
assign A437z6 = (G537z6 & O537z6);
assign O537z6 = (~(Lgj7z6[67] & Rphov6));
assign G537z6 = (~(J6oiw6 & Lgj7z6[70]));
assign Y037z6 = (W537z6 & E637z6);
assign E637z6 = (M637z6 & U637z6);
assign U637z6 = (C737z6 & K737z6);
assign K737z6 = (~(Lgj7z6[73] & Uy2jy6));
assign C737z6 = (~(Lgj7z6[76] & Mbj7x6));
assign M637z6 = (S737z6 & A837z6);
assign A837z6 = (~(Lgj7z6[79] & Nfj7x6));
assign S737z6 = (~(Lgj7z6[82] & Hzh7x6));
assign W537z6 = (I837z6 & Q837z6);
assign Q837z6 = (Y837z6 & G937z6);
assign G937z6 = (~(Lgj7z6[85] & L1i7x6));
assign Y837z6 = (~(Jrj7x6 & Lgj7z6[88]));
assign I837z6 = (O937z6 & W937z6);
assign W937z6 = (~(Lgj7z6[91] & P3i7x6));
assign O937z6 = (~(Lgj7z6[94] & V6i7x6));
assign Qk27z6 = (Ea37z6 & Ma37z6);
assign Ma37z6 = (~(Maajy6 & Ua37z6));
assign Ua37z6 = (~(Cb37z6 & Kb37z6));
assign Kb37z6 = (Sb37z6 & Ac37z6);
assign Ac37z6 = (Ic37z6 & Qc37z6);
assign Qc37z6 = (Yc37z6 & Gd37z6);
assign Gd37z6 = (~(Lgj7z6[97] & Ao2jy6));
assign Yc37z6 = (~(Lgj7z6[100] & Nuniw6));
assign Ic37z6 = (Od37z6 & Wd37z6);
assign Wd37z6 = (~(Lgj7z6[103] & Jfmiw6));
assign Od37z6 = (~(Lgj7z6[106] & Cn2jy6));
assign Sb37z6 = (Ee37z6 & Me37z6);
assign Me37z6 = (Ue37z6 & Cf37z6);
assign Cf37z6 = (~(Lgj7z6[109] & Cshov6));
assign Ue37z6 = (~(Lgj7z6[112] & I2oiw6));
assign Ee37z6 = (Kf37z6 & Sf37z6);
assign Sf37z6 = (~(Lgj7z6[115] & Rphov6));
assign Kf37z6 = (~(Lgj7z6[118] & J6oiw6));
assign Cb37z6 = (Ag37z6 & Ig37z6);
assign Ig37z6 = (Qg37z6 & Yg37z6);
assign Yg37z6 = (Gh37z6 & Oh37z6);
assign Oh37z6 = (~(Lgj7z6[121] & Uy2jy6));
assign Gh37z6 = (~(Lgj7z6[124] & Mbj7x6));
assign Qg37z6 = (Wh37z6 & Ei37z6);
assign Ei37z6 = (~(Lgj7z6[127] & Nfj7x6));
assign Wh37z6 = (~(Lgj7z6[130] & Hzh7x6));
assign Ag37z6 = (Mi37z6 & Ui37z6);
assign Ui37z6 = (Cj37z6 & Kj37z6);
assign Kj37z6 = (~(Lgj7z6[133] & L1i7x6));
assign Cj37z6 = (~(Lgj7z6[136] & Jrj7x6));
assign Mi37z6 = (Sj37z6 & Ak37z6);
assign Ak37z6 = (~(Lgj7z6[139] & P3i7x6));
assign Sj37z6 = (~(Lgj7z6[142] & V6i7x6));
assign Ea37z6 = (~(A87jy6 & Ik37z6));
assign Ik37z6 = (~(Qk37z6 & Yk37z6));
assign Yk37z6 = (Gl37z6 & Ol37z6);
assign Ol37z6 = (Wl37z6 & Em37z6);
assign Em37z6 = (Mm37z6 & Um37z6);
assign Um37z6 = (~(Lgj7z6[145] & Ao2jy6));
assign Mm37z6 = (~(Lgj7z6[148] & Nuniw6));
assign Wl37z6 = (Cn37z6 & Kn37z6);
assign Kn37z6 = (~(Lgj7z6[151] & Jfmiw6));
assign Cn37z6 = (~(Lgj7z6[154] & Cn2jy6));
assign Gl37z6 = (Sn37z6 & Ao37z6);
assign Ao37z6 = (Io37z6 & Qo37z6);
assign Qo37z6 = (~(Lgj7z6[157] & Cshov6));
assign Io37z6 = (~(Lgj7z6[160] & I2oiw6));
assign Sn37z6 = (Yo37z6 & Gp37z6);
assign Gp37z6 = (~(Lgj7z6[163] & Rphov6));
assign Yo37z6 = (~(Lgj7z6[166] & J6oiw6));
assign Qk37z6 = (Op37z6 & Wp37z6);
assign Wp37z6 = (Eq37z6 & Mq37z6);
assign Mq37z6 = (Uq37z6 & Cr37z6);
assign Cr37z6 = (~(Lgj7z6[169] & Uy2jy6));
assign Uq37z6 = (~(Lgj7z6[172] & Mbj7x6));
assign Eq37z6 = (Kr37z6 & Sr37z6);
assign Sr37z6 = (~(Lgj7z6[175] & Nfj7x6));
assign Kr37z6 = (~(Lgj7z6[178] & Hzh7x6));
assign Op37z6 = (As37z6 & Is37z6);
assign Is37z6 = (Qs37z6 & Ys37z6);
assign Ys37z6 = (~(Lgj7z6[181] & L1i7x6));
assign Qs37z6 = (~(Lgj7z6[184] & Jrj7x6));
assign As37z6 = (Gt37z6 & Ot37z6);
assign Ot37z6 = (~(Lgj7z6[187] & P3i7x6));
assign Gt37z6 = (~(Lgj7z6[190] & V6i7x6));
assign CURRPRI[5] = (~(Wt37z6 & Eu37z6));
assign Eu37z6 = (Mu37z6 & Uu37z6);
assign Uu37z6 = (~(Sz3jy6 & Cv37z6));
assign Cv37z6 = (~(Kv37z6 & Sv37z6));
assign Sv37z6 = (Aw37z6 & Iw37z6);
assign Iw37z6 = (Qw37z6 & Yw37z6);
assign Yw37z6 = (~(Ao2jy6 & M018x6));
assign M018x6 = (~(Q8oiy6 & J92nv6));
assign J92nv6 = (Gx37z6 | Ppb7z6[5]);
assign Gx37z6 = (Ppb7z6[6] | Ppb7z6[7]);
assign Q8oiy6 = (!Ppb7z6[5]);
assign Qw37z6 = (~(Ffj7z6[0] & Cshov6));
assign Aw37z6 = (Ox37z6 & Wx37z6);
assign Wx37z6 = (~(Zdj7z6[0] & I2oiw6));
assign Ox37z6 = (~(Tcj7z6[0] & Rphov6));
assign Kv37z6 = (Ey37z6 & My37z6);
assign My37z6 = (Uy37z6 & Cz37z6);
assign Cz37z6 = (~(Gaj7z6[0] & Hzh7x6));
assign Uy37z6 = (~(Nbj7z6[0] & L1i7x6));
assign Ey37z6 = (Kz37z6 & Sz37z6);
assign Sz37z6 = (~(Z8j7z6[0] & P3i7x6));
assign Kz37z6 = (~(T7j7z6[0] & V6i7x6));
assign Sz3jy6 = (Ox3jy6 & Pqliw6);
assign Ox3jy6 = (S73jy6 & Omliw6);
assign Mu37z6 = (A047z6 & I047z6);
assign I047z6 = (~(Wtgjy6 & Q047z6));
assign Q047z6 = (~(Y047z6 & G147z6));
assign G147z6 = (O147z6 & W147z6);
assign W147z6 = (E247z6 & M247z6);
assign M247z6 = (U247z6 & C347z6);
assign C347z6 = (~(Lgj7z6[0] & Ao2jy6));
assign U247z6 = (~(Lgj7z6[3] & Nuniw6));
assign E247z6 = (K347z6 & S347z6);
assign S347z6 = (~(Lgj7z6[6] & Jfmiw6));
assign K347z6 = (~(Lgj7z6[9] & Cn2jy6));
assign O147z6 = (A447z6 & I447z6);
assign I447z6 = (Q447z6 & Y447z6);
assign Y447z6 = (~(Lgj7z6[12] & Cshov6));
assign Q447z6 = (~(Lgj7z6[15] & I2oiw6));
assign A447z6 = (G547z6 & O547z6);
assign O547z6 = (~(Lgj7z6[18] & Rphov6));
assign G547z6 = (~(Lgj7z6[21] & J6oiw6));
assign Y047z6 = (W547z6 & E647z6);
assign E647z6 = (M647z6 & U647z6);
assign U647z6 = (C747z6 & K747z6);
assign K747z6 = (~(Lgj7z6[24] & Uy2jy6));
assign C747z6 = (~(Lgj7z6[27] & Mbj7x6));
assign M647z6 = (S747z6 & A847z6);
assign A847z6 = (~(Lgj7z6[30] & Nfj7x6));
assign S747z6 = (~(Lgj7z6[33] & Hzh7x6));
assign W547z6 = (I847z6 & Q847z6);
assign Q847z6 = (Y847z6 & G947z6);
assign G947z6 = (~(Lgj7z6[36] & L1i7x6));
assign Y847z6 = (~(Lgj7z6[39] & Jrj7x6));
assign I847z6 = (O947z6 & W947z6);
assign W947z6 = (~(Lgj7z6[42] & P3i7x6));
assign O947z6 = (~(Lgj7z6[45] & V6i7x6));
assign Wtgjy6 = (Ea47z6 & S73jy6);
assign S73jy6 = (~(Nob7z6[5] | Nob7z6[6]));
assign Ea47z6 = (Nob7z6[4] & Pqliw6);
assign A047z6 = (~(Awcjy6 & Ma47z6));
assign Ma47z6 = (~(Ua47z6 & Cb47z6));
assign Cb47z6 = (Kb47z6 & Sb47z6);
assign Sb47z6 = (Ac47z6 & Ic47z6);
assign Ic47z6 = (Qc47z6 & Yc47z6);
assign Yc47z6 = (~(Lgj7z6[48] & Ao2jy6));
assign Qc47z6 = (~(Lgj7z6[51] & Nuniw6));
assign Ac47z6 = (Gd47z6 & Od47z6);
assign Od47z6 = (~(Lgj7z6[54] & Jfmiw6));
assign Gd47z6 = (~(Lgj7z6[57] & Cn2jy6));
assign Kb47z6 = (Wd47z6 & Ee47z6);
assign Ee47z6 = (Me47z6 & Ue47z6);
assign Ue47z6 = (~(Cshov6 & Lgj7z6[60]));
assign Me47z6 = (~(Lgj7z6[63] & I2oiw6));
assign Wd47z6 = (Cf47z6 & Kf47z6);
assign Kf47z6 = (~(Lgj7z6[66] & Rphov6));
assign Cf47z6 = (~(Lgj7z6[69] & J6oiw6));
assign Ua47z6 = (Sf47z6 & Ag47z6);
assign Ag47z6 = (Ig47z6 & Qg47z6);
assign Qg47z6 = (Yg47z6 & Gh47z6);
assign Gh47z6 = (~(Lgj7z6[72] & Uy2jy6));
assign Yg47z6 = (~(Lgj7z6[75] & Mbj7x6));
assign Ig47z6 = (Oh47z6 & Wh47z6);
assign Wh47z6 = (~(Lgj7z6[78] & Nfj7x6));
assign Oh47z6 = (~(Lgj7z6[81] & Hzh7x6));
assign Sf47z6 = (Ei47z6 & Mi47z6);
assign Mi47z6 = (Ui47z6 & Cj47z6);
assign Cj47z6 = (~(Lgj7z6[84] & L1i7x6));
assign Ui47z6 = (~(Lgj7z6[87] & Jrj7x6));
assign Ei47z6 = (Kj47z6 & Sj47z6);
assign Sj47z6 = (~(Lgj7z6[90] & P3i7x6));
assign Kj47z6 = (~(Lgj7z6[93] & V6i7x6));
assign Awcjy6 = (~(Ak47z6 | Nob7z6[4]));
assign Wt37z6 = (Ik47z6 & Qk47z6);
assign Qk47z6 = (~(Maajy6 & Yk47z6));
assign Yk47z6 = (~(Gl47z6 & Ol47z6));
assign Ol47z6 = (Wl47z6 & Em47z6);
assign Em47z6 = (Mm47z6 & Um47z6);
assign Um47z6 = (Cn47z6 & Kn47z6);
assign Kn47z6 = (~(Lgj7z6[96] & Ao2jy6));
assign Cn47z6 = (~(Lgj7z6[99] & Nuniw6));
assign Mm47z6 = (Sn47z6 & Ao47z6);
assign Ao47z6 = (~(Lgj7z6[102] & Jfmiw6));
assign Sn47z6 = (~(Lgj7z6[105] & Cn2jy6));
assign Wl47z6 = (Io47z6 & Qo47z6);
assign Qo47z6 = (Yo47z6 & Gp47z6);
assign Gp47z6 = (~(Lgj7z6[108] & Cshov6));
assign Yo47z6 = (~(Lgj7z6[111] & I2oiw6));
assign Io47z6 = (Op47z6 & Wp47z6);
assign Wp47z6 = (~(Lgj7z6[114] & Rphov6));
assign Op47z6 = (~(Lgj7z6[117] & J6oiw6));
assign Gl47z6 = (Eq47z6 & Mq47z6);
assign Mq47z6 = (Uq47z6 & Cr47z6);
assign Cr47z6 = (Kr47z6 & Sr47z6);
assign Sr47z6 = (~(Lgj7z6[120] & Uy2jy6));
assign Kr47z6 = (~(Lgj7z6[123] & Mbj7x6));
assign Uq47z6 = (As47z6 & Is47z6);
assign Is47z6 = (~(Lgj7z6[126] & Nfj7x6));
assign As47z6 = (~(Lgj7z6[129] & Hzh7x6));
assign Eq47z6 = (Qs47z6 & Ys47z6);
assign Ys47z6 = (Gt47z6 & Ot47z6);
assign Ot47z6 = (~(Lgj7z6[132] & L1i7x6));
assign Gt47z6 = (~(Lgj7z6[135] & Jrj7x6));
assign Qs47z6 = (Wt47z6 & Eu47z6);
assign Eu47z6 = (~(Lgj7z6[138] & P3i7x6));
assign Wt47z6 = (~(Lgj7z6[141] & V6i7x6));
assign Maajy6 = (~(Ak47z6 | Omliw6));
assign Ak47z6 = (~(Mu47z6 & Nob7z6[5]));
assign Mu47z6 = (Gpliw6 & Pqliw6);
assign Gpliw6 = (!Nob7z6[6]);
assign Ik47z6 = (~(A87jy6 & Uu47z6));
assign Uu47z6 = (~(Cv47z6 & Kv47z6));
assign Kv47z6 = (Sv47z6 & Aw47z6);
assign Aw47z6 = (Iw47z6 & Qw47z6);
assign Qw47z6 = (Yw47z6 & Gx47z6);
assign Gx47z6 = (~(Lgj7z6[144] & Ao2jy6));
assign Ao2jy6 = (!Rqmiw6);
assign Rqmiw6 = (~(Ox47z6 & Me3jy6));
assign Ox47z6 = (Giliw6 & Flliw6);
assign Yw47z6 = (~(Lgj7z6[147] & Nuniw6));
assign Nuniw6 = (!Daoiw6);
assign Daoiw6 = (~(Qc3jy6 & Kf3jy6));
assign Iw47z6 = (Wx47z6 & Ey47z6);
assign Ey47z6 = (~(Lgj7z6[150] & Jfmiw6));
assign Jfmiw6 = (!Zumiw6);
assign Zumiw6 = (~(My47z6 & Me3jy6));
assign My47z6 = (Nob7z6[1] & Flliw6);
assign Wx47z6 = (~(Lgj7z6[153] & Cn2jy6));
assign Cn2jy6 = (!Xdoiw6);
assign Xdoiw6 = (~(Qc3jy6 & Uy47z6));
assign Qc3jy6 = (Wjliw6 & Flliw6);
assign Sv47z6 = (Cz47z6 & Kz47z6);
assign Kz47z6 = (Sz47z6 & A057z6);
assign A057z6 = (~(Lgj7z6[156] & Cshov6));
assign Cshov6 = (!Ue5jy6);
assign Ue5jy6 = (~(I057z6 & Ee3jy6));
assign Sz47z6 = (~(Lgj7z6[159] & I2oiw6));
assign I2oiw6 = (Kf3jy6 & Ee3jy6);
assign Cz47z6 = (Q057z6 & Y057z6);
assign Y057z6 = (~(Lgj7z6[162] & Rphov6));
assign Rphov6 = (Ee3jy6 & Gh3jy6);
assign Q057z6 = (~(Lgj7z6[165] & J6oiw6));
assign J6oiw6 = (Uy47z6 & Ee3jy6);
assign Ee3jy6 = (Nob7z6[2] & Flliw6);
assign Cv47z6 = (G157z6 & O157z6);
assign O157z6 = (W157z6 & E257z6);
assign E257z6 = (M257z6 & U257z6);
assign U257z6 = (~(Lgj7z6[168] & Uy2jy6));
assign Uy2jy6 = (Cz3jy6 & Giliw6);
assign M257z6 = (~(Lgj7z6[171] & Mbj7x6));
assign Mbj7x6 = (!U7k7x6);
assign U7k7x6 = (~(C357z6 & Kf3jy6));
assign W157z6 = (K357z6 & S357z6);
assign S357z6 = (~(Lgj7z6[174] & Nfj7x6));
assign Nfj7x6 = (Cz3jy6 & Nob7z6[1]);
assign Cz3jy6 = (Me3jy6 & Nob7z6[3]);
assign Me3jy6 = (~(Nob7z6[0] | Nob7z6[2]));
assign K357z6 = (~(Lgj7z6[177] & Hzh7x6));
assign Hzh7x6 = (!Pfk7x6);
assign Pfk7x6 = (~(C357z6 & Uy47z6));
assign C357z6 = (Nob7z6[3] & Wjliw6);
assign G157z6 = (A457z6 & I457z6);
assign I457z6 = (Q457z6 & Y457z6);
assign Y457z6 = (~(Lgj7z6[180] & L1i7x6));
assign L1i7x6 = (!Qpl7x6);
assign Qpl7x6 = (~(I057z6 & Yc3jy6));
assign I057z6 = (Krliw6 & Giliw6);
assign Q457z6 = (~(Lgj7z6[183] & Jrj7x6));
assign Jrj7x6 = (Yc3jy6 & Kf3jy6);
assign Kf3jy6 = (~(Krliw6 | Nob7z6[1]));
assign A457z6 = (G557z6 & O557z6);
assign O557z6 = (~(Lgj7z6[186] & P3i7x6));
assign P3i7x6 = (Yc3jy6 & Gh3jy6);
assign Gh3jy6 = (~(Giliw6 | Nob7z6[0]));
assign G557z6 = (~(Lgj7z6[189] & V6i7x6));
assign V6i7x6 = (Yc3jy6 & Uy47z6);
assign Uy47z6 = (~(Krliw6 | Giliw6));
assign Giliw6 = (!Nob7z6[1]);
assign Krliw6 = (!Nob7z6[0]);
assign Yc3jy6 = (~(Wjliw6 | Flliw6));
assign Flliw6 = (!Nob7z6[3]);
assign Wjliw6 = (!Nob7z6[2]);
assign A87jy6 = (W557z6 & E657z6);
assign E657z6 = (Xnliw6 & Pqliw6);
assign Pqliw6 = (!Nob7z6[7]);
assign Xnliw6 = (!Nob7z6[5]);
assign W557z6 = (Nob7z6[6] & Omliw6);
assign Omliw6 = (!Nob7z6[4]);
assign BRCHSTAT[2] = (M657z6 & Aciiy6);
assign M657z6 = (~(U657z6 & C757z6));
assign C757z6 = (~(V9mnv6 & K757z6));
assign K757z6 = (Csohw6 | Rrnnv6);
assign U657z6 = (~(S757z6 | Ir0ov6));
assign BRCHSTAT[1] = (~(A857z6 & I857z6));
assign I857z6 = (~(Camnv6 & Q857z6));
assign Q857z6 = (Jamnv6 | S757z6);
assign Jamnv6 = (~(Pcmhw6 & Y857z6));
assign Y857z6 = (~(V9mnv6 & G957z6));
assign G957z6 = (Vmnnv6 | Amnnv6);
assign Amnnv6 = (Nginv6 | Rrnnv6);
assign Rrnnv6 = (U6uiy6 & Zec7z6[28]);
assign Vmnnv6 = (~(Sfohw6 & U9inv6));
assign Sfohw6 = (!Csohw6);
assign Csohw6 = (Yksiy6 & O957z6);
assign Pcmhw6 = (!Ir0ov6);
assign Ir0ov6 = (V9mnv6 & Awiiy6);
assign Awiiy6 = (W957z6 & Ea57z6);
assign Ea57z6 = (Ma57z6 & Ua57z6);
assign Camnv6 = (!Aciiy6);
assign A857z6 = (~(V9mnv6 & Cb57z6));
assign Cb57z6 = (~(Kb57z6 & Sb57z6));
assign Sb57z6 = (U9inv6 | Zec7z6[7]);
assign Kb57z6 = (Ac57z6 & A2sov6);
assign Ac57z6 = (~(Nginv6 & Painv6));
assign BRCHSTAT[0] = (S757z6 | Ic57z6);
assign Ic57z6 = (V9mnv6 & Qc57z6);
assign Qc57z6 = (~(A2sov6 & Yc57z6));
assign Yc57z6 = (~(Gd57z6 & Aciiy6));
assign Aciiy6 = (~(Od57z6 & Wd57z6));
assign Wd57z6 = (Wqfov6 | Gpsiw6);
assign Gpsiw6 = (Cmbdt6 | L2gdt6);
assign Od57z6 = (~(N6xiw6 & Drfov6));
assign Drfov6 = (!L2gdt6);
assign N6xiw6 = (!Ghkiy6);
assign Ghkiy6 = (~(Ee57z6 & Ashnv6));
assign Ashnv6 = (Yrfov6 | L2gdt6);
assign Ee57z6 = (S6cdt6 | Yrfov6);
assign Yrfov6 = (~(Wqfov6 | Ohe7z6[4]));
assign Wqfov6 = (Me57z6 | Ohe7z6[1]);
assign Me57z6 = (Ohe7z6[2] | Ohe7z6[3]);
assign Gd57z6 = (~(Flnnv6 & Htnnv6));
assign Htnnv6 = (~(Nginv6 & Zec7z6[10]));
assign Nginv6 = (Ue57z6 & Cf57z6);
assign Cf57z6 = (~(Kf57z6 | I5cdt6));
assign Kf57z6 = (~(Sf57z6 & Adohw6));
assign Ue57z6 = (U6uiy6 & K7uiy6);
assign K7uiy6 = (!Cvtiy6);
assign Flnnv6 = (U9inv6 | Xeinv6);
assign U9inv6 = (T1sov6 | I5cdt6);
assign T1sov6 = (~(Ag57z6 & Xgmhw6));
assign Xgmhw6 = (Ig57z6 & Zec7z6[15]);
assign Ig57z6 = (Zec7z6[14] & Uqsiy6);
assign Ag57z6 = (~(D6siw6 | Z3fhw6));
assign Z3fhw6 = (Cvehw6 & Zec7z6[11]);
assign A2sov6 = (!Btpiw6);
assign Btpiw6 = (S3riy6 & Painv6);
assign S3riy6 = (I5fhw6 & Zec7z6[8]);
assign S757z6 = (V9mnv6 & Qg57z6);
assign Qg57z6 = (~(Bhaov6 & Ofmhw6));
assign Ofmhw6 = (Yg57z6 & Gh57z6);
assign Gh57z6 = (Oh57z6 & Jkc7x6);
assign Jkc7x6 = (~(Agmiy6 & Zec7z6[4]));
assign Agmiy6 = (~(Cvmiy6 | Elviw6));
assign Elviw6 = (!Zec7z6[31]);
assign Cvmiy6 = (~(Wh57z6 & Eauiy6));
assign Wh57z6 = (Xqwiw6 & Fcinv6);
assign Xqwiw6 = (B0xiw6 | Obwiw6);
assign B0xiw6 = (Zec7z6[8] & Xeinv6);
assign Oh57z6 = (~(Igmiy6 | Znvnv6));
assign Znvnv6 = (Sfiiy6 & Sjtiy6);
assign Sjtiy6 = (Ei57z6 & W9tiy6);
assign Ei57z6 = (Gbfhw6 & Bainv6);
assign Igmiy6 = (Qkc7x6 & Zec7z6[8]);
assign Qkc7x6 = (Mqiiy6 & Zec7z6[11]);
assign Mqiiy6 = (I5fhw6 & Gbfhw6);
assign Gbfhw6 = (Zec7z6[10] & Qeinv6);
assign I5fhw6 = (~(Kntiy6 | D6siw6));
assign Kntiy6 = (!Sntiy6);
assign Sntiy6 = (Mi57z6 & Zec7z6[15]);
assign Mi57z6 = (Zec7z6[13] & Sbtiy6);
assign Sbtiy6 = (!Zec7z6[14]);
assign Yg57z6 = (Ui57z6 & Cj57z6);
assign Cj57z6 = (~(Kj57z6 & Sj57z6));
assign Sj57z6 = (Ak57z6 & Ik57z6);
assign Ik57z6 = (Qk57z6 & O957z6);
assign Qk57z6 = (Yk57z6 & Bainv6);
assign Yk57z6 = (Gl57z6 | Hxihw6);
assign Hxihw6 = (!U2uiy6);
assign U2uiy6 = (Xeinv6 & Rktov6);
assign Rktov6 = (!K0riw6);
assign K0riw6 = (Ol57z6 & Zec7z6[3]);
assign Ol57z6 = (!Wl57z6);
assign Gl57z6 = (Zec7z6[27] ? Utihw6 : Em57z6);
assign Utihw6 = (!Kzqiy6);
assign Em57z6 = (Mm57z6 & Um57z6);
assign Um57z6 = (Cn57z6 & Buihw6);
assign Buihw6 = (!Zec7z6[25]);
assign Mm57z6 = (Kzqiy6 & Kn57z6);
assign Kzqiy6 = (Lofhw6 & Jlohw6);
assign Jlohw6 = (!Zec7z6[26]);
assign Lofhw6 = (!Zec7z6[24]);
assign Ak57z6 = (Q8riy6 & Zec7z6[30]);
assign Q8riy6 = (Zec7z6[28] & Zec7z6[29]);
assign Kj57z6 = (Sn57z6 & Ao57z6);
assign Ao57z6 = (Io57z6 & Zec7z6[12]);
assign Io57z6 = (Zec7z6[11] & Zec7z6[31]);
assign Sn57z6 = (Qo57z6 & Zec7z6[4]);
assign Qo57z6 = (Nbfhw6 & Kdfhw6);
assign Ui57z6 = (~(Yo57z6 & Gp57z6));
assign Gp57z6 = (Kn57z6 & Cn57z6);
assign Kn57z6 = (!Zec7z6[22]);
assign Yo57z6 = (Cbuiy6 & Op57z6);
assign Op57z6 = (!Zec7z6[21]);
assign Cbuiy6 = (Wp57z6 & Eq57z6);
assign Eq57z6 = (Obwiw6 & Nbfhw6);
assign Nbfhw6 = (Zec7z6[6] & Zpehw6);
assign Zpehw6 = (!Zec7z6[5]);
assign Obwiw6 = (Zec7z6[7] & Bainv6);
assign Wp57z6 = (Zec7z6[4] & Eauiy6);
assign Eauiy6 = (Kdfhw6 & Zhmhw6);
assign Zhmhw6 = (Ydfhw6 & O957z6);
assign Ydfhw6 = (Zec7z6[11] & D6siw6);
assign Kdfhw6 = (Painv6 & Qeinv6);
assign Qeinv6 = (!Zec7z6[9]);
assign Bhaov6 = (Mq57z6 & Uq57z6);
assign Uq57z6 = (~(Cr57z6 & Kr57z6));
assign Kr57z6 = (Sr57z6 & As57z6);
assign As57z6 = (Is57z6 & Qs57z6);
assign Qs57z6 = (!Zec7z6[20]);
assign Is57z6 = (Cn57z6 & Sf57z6);
assign Sf57z6 = (!Zec7z6[28]);
assign Cn57z6 = (!Zec7z6[23]);
assign Sr57z6 = (Zec7z6[22] & Zec7z6[21]);
assign Cr57z6 = (Ys57z6 & Gt57z6);
assign Gt57z6 = (Ot57z6 & Cvtiy6);
assign Cvtiy6 = (Sywiw6 & Zec7z6[9]);
assign Sywiw6 = (~(Xeinv6 | Bainv6));
assign Ot57z6 = (U6uiy6 & Zec7z6[4]);
assign U6uiy6 = (M2uiy6 & Zec7z6[31]);
assign M2uiy6 = (Wt57z6 & Zec7z6[12]);
assign Wt57z6 = (O957z6 & Gginv6);
assign Ys57z6 = (E3fhw6 & H2riw6);
assign H2riw6 = (Painv6 & Adohw6);
assign Adohw6 = (!Zec7z6[30]);
assign Painv6 = (!Zec7z6[10]);
assign E3fhw6 = (Zec7z6[5] & Fcinv6);
assign Fcinv6 = (!Zec7z6[6]);
assign Mq57z6 = (~(Ua57z6 & Eu57z6));
assign Eu57z6 = (~(W957z6 & Ma57z6));
assign Ma57z6 = (~(Zec7z6[3] | X0cdt6));
assign W957z6 = (Qzuiw6 & Zec7z6[4]);
assign Qzuiw6 = (Zec7z6[5] & Zec7z6[6]);
assign Ua57z6 = (~(Mu57z6 & Amtov6));
assign Amtov6 = (~(Uu57z6 & W9tiy6));
assign Uu57z6 = (Cvehw6 & Zec7z6[8]);
assign Mu57z6 = (Q9fhw6 | Aktiy6);
assign Aktiy6 = (!Sfiiy6);
assign Sfiiy6 = (~(Wl57z6 | Xeinv6));
assign Xeinv6 = (!Zec7z6[7]);
assign Wl57z6 = (~(Cv57z6 & Zec7z6[2]));
assign Cv57z6 = (Zec7z6[1] & Zec7z6[0]);
assign Q9fhw6 = (~(Kv57z6 & W9tiy6));
assign W9tiy6 = (Yksiy6 & Gpuiy6);
assign Gpuiy6 = (!Icuiy6);
assign Icuiy6 = (~(Sv57z6 & Zec7z6[14]));
assign Sv57z6 = (Uqsiy6 & Eqsiy6);
assign Eqsiy6 = (!Zec7z6[15]);
assign Uqsiy6 = (!Zec7z6[13]);
assign Kv57z6 = (Cvehw6 & Bainv6);
assign Bainv6 = (!Zec7z6[8]);
assign Cvehw6 = (Zec7z6[10] & Zec7z6[9]);
assign V9mnv6 = (Aw57z6 & Iw57z6);
assign Iw57z6 = (Qw57z6 & Yw57z6);
assign Yw57z6 = (Gx57z6 & Fetov6);
assign Fetov6 = (!Pacdt6);
assign Gx57z6 = (~(Efcdt6 | Vjddt6));
assign Qw57z6 = (Ox57z6 & Wx57z6);
assign Wx57z6 = (~(Ey57z6 & My57z6));
assign My57z6 = (~(Uy57z6 & Cz57z6));
assign Cz57z6 = (~(Bfd7z6[1] & Otiiy6));
assign Uy57z6 = (Nbtov6 & D6tov6);
assign D6tov6 = (!Bfd7z6[3]);
assign Nbtov6 = (!Bfd7z6[2]);
assign Ey57z6 = (L9d7z6[3] | L9d7z6[2]);
assign Ox57z6 = (~(Myuiy6 | L9cdt6));
assign Myuiy6 = (Kz57z6 & Sz57z6);
assign Sz57z6 = (~(Fjaov6 | Pacdt6));
assign Fjaov6 = (G597z6 & A067z6);
assign A067z6 = (~(I067z6 & Q067z6));
assign Q067z6 = (~(Pmc7z6[1] & W1k6z6));
assign W1k6z6 = (Y067z6 ^ Lpc7z6[1]);
assign I067z6 = (G167z6 & O167z6);
assign O167z6 = (~(Pmc7z6[2] & W167z6));
assign G167z6 = (~(Pmc7z6[0] & O1k6z6));
assign Kz57z6 = (E267z6 & Igiiy6);
assign Igiiy6 = (~(Yiaov6 & M267z6));
assign M267z6 = (U267z6 | Bfd7z6[0]);
assign U267z6 = (Bfd7z6[2] | Bfd7z6[4]);
assign E267z6 = (~(Yiaov6 & Kbriy6));
assign Kbriy6 = (!Otiiy6);
assign Yiaov6 = (C367z6 & G597z6);
assign C367z6 = (W167z6 ? Pmc7z6[1] : K367z6);
assign W167z6 = (~(Y067z6 | Lpc7z6[1]));
assign K367z6 = (O1k6z6 | Pmc7z6[0]);
assign O1k6z6 = (Lpc7z6[1] & Y067z6);
assign Y067z6 = (!Lpc7z6[0]);
assign Aw57z6 = (S367z6 & A467z6);
assign A467z6 = (I467z6 & K3jnv6);
assign K3jnv6 = (~(Q467z6 | Y807z6));
assign Y807z6 = (Y3fet6 & Qg2nv6);
assign Q467z6 = (~(SLEEPHOLDACKn & W8h7v6));
assign SLEEPHOLDACKn = (!Gwj8v6);
assign Gwj8v6 = (D2fet6 & Qg2nv6);
assign Qg2nv6 = (!Tnzdt6);
assign I467z6 = (Y467z6 & G567z6);
assign G567z6 = (~(O567z6 & W567z6));
assign W567z6 = (L9d7z6[1] | L9d7z6[0]);
assign O567z6 = (~(E667z6 & M667z6));
assign M667z6 = (~(Bfd7z6[5] & Otiiy6));
assign E667z6 = (~(Bfd7z6[0] | Bfd7z6[1]));
assign Y467z6 = (~(U667z6 & C767z6));
assign C767z6 = (L9d7z6[5] | L9d7z6[4]);
assign U667z6 = (~(K767z6 & S767z6));
assign S767z6 = (~(Bfd7z6[3] & Otiiy6));
assign Otiiy6 = (O957z6 & Kbtiy6);
assign Kbtiy6 = (!Yksiy6);
assign Yksiy6 = (Gginv6 & D6siw6);
assign D6siw6 = (!Zec7z6[12]);
assign Gginv6 = (!Zec7z6[11]);
assign O957z6 = (A867z6 & Zec7z6[15]);
assign A867z6 = (Zec7z6[14] & Zec7z6[13]);
assign K767z6 = (~(Bfd7z6[4] | Bfd7z6[5]));
assign S367z6 = (O4piw6 & Ktfxx6);
assign Ktfxx6 = (~(Ddmhw6 | Qdcdt6));
assign Ddmhw6 = (Tk8iw6 ? Osd7z6[1] : Osd7z6[2]);
assign Tk8iw6 = (Myhiy6 & Iwhiy6);
assign Iwhiy6 = (I867z6 & Q867z6);
assign Q867z6 = (Y867z6 & G967z6);
assign G967z6 = (~(O967z6 | Fhc7z6[15]));
assign O967z6 = (Fhc7z6[8] | Fhc7z6[9]);
assign Y867z6 = (~(Fhc7z6[13] | Fhc7z6[14]));
assign I867z6 = (W967z6 & Ea67z6);
assign Ea67z6 = (~(Fhc7z6[11] | Fhc7z6[12]));
assign W967z6 = (~(Q4oiy6 | Fhc7z6[10]));
assign Q4oiy6 = (~(Ma67z6 & Ua67z6));
assign Ua67z6 = (Cb67z6 & Kb67z6);
assign Kb67z6 = (~(Fhc7z6[6] | Fhc7z6[7]));
assign Cb67z6 = (~(E3c7z6[4] | Fhc7z6[5]));
assign Ma67z6 = (Sb67z6 & Ac67z6);
assign Ac67z6 = (~(E3c7z6[2] | E3c7z6[3]));
assign Sb67z6 = (~(E3c7z6[0] | E3c7z6[1]));
assign Myhiy6 = (!Lntiw6);
assign Lntiw6 = (~(Ic67z6 & Qc67z6));
assign Qc67z6 = (Yc67z6 & Gd67z6);
assign Gd67z6 = (Od67z6 & Wd67z6);
assign Wd67z6 = (~(Fhc7z6[30] | Fhc7z6[31]));
assign Od67z6 = (~(Fhc7z6[28] | Fhc7z6[29]));
assign Yc67z6 = (Ee67z6 & Me67z6);
assign Me67z6 = (~(Fhc7z6[26] | Fhc7z6[27]));
assign Ee67z6 = (~(Fhc7z6[24] | Fhc7z6[25]));
assign Ic67z6 = (Ue67z6 & Cf67z6);
assign Cf67z6 = (Kf67z6 & Sf67z6);
assign Sf67z6 = (~(Fhc7z6[22] | Fhc7z6[23]));
assign Kf67z6 = (~(Fhc7z6[20] | Fhc7z6[21]));
assign Ue67z6 = (Ag67z6 & Ig67z6);
assign Ig67z6 = (~(Fhc7z6[18] | Fhc7z6[19]));
assign Ag67z6 = (~(Fhc7z6[16] | Fhc7z6[17]));
assign O4piw6 = (Ldo7v6 & X6xnv6);
assign X6xnv6 = (~(Kzy6z6 & I51ov6));
assign I51ov6 = (Cgc7z6[3] & O4jhw6);
assign O4jhw6 = (!Cgc7z6[0]);
assign Kzy6z6 = (P1piw6 & A4jhw6);
assign A4jhw6 = (!Cgc7z6[2]);
assign P1piw6 = (!Cgc7z6[1]);

always @(posedge FCLK or negedge PORESETn)
  if(~PORESETn)
    Sj2nz6 <= 1'b0;
  else
    Sj2nz6 <= 1'b1;

always @(posedge FCLK or negedge PORESETn)
  if(~PORESETn)
    Ik2nz6 <= 1'b0;
  else
    Ik2nz6 <= M4adt6;

always @(posedge FCLK or negedge SYSRESETn)
  if(~SYSRESETn)
    Zk2nz6 <= 1'b0;
  else
    Zk2nz6 <= 1'b1;

always @(posedge FCLK or negedge SYSRESETn)
  if(~SYSRESETn)
    Ql2nz6 <= 1'b0;
  else
    Ql2nz6 <= Y4adt6;

always @(posedge SWCLKTCK or negedge PORESETn)
  if(~PORESETn)
    Im2nz6 <= 1'b0;
  else
    Im2nz6 <= 1'b1;

always @(posedge SWCLKTCK or negedge PORESETn)
  if(~PORESETn)
    Ym2nz6 <= 1'b0;
  else
    Ym2nz6 <= L5adt6;

always @(posedge TRACECLKIN or negedge Ox9dt6)
  if(~Ox9dt6)
    Pn2nz6 <= 1'b0;
  else
    Pn2nz6 <= Ox9dt6;

always @(posedge TRACECLKIN or negedge Ox9dt6)
  if(~Ox9dt6)
    Go2nz6 <= 1'b0;
  else
    Go2nz6 <= X5adt6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yo2nz6 <= 1'b0;
  else
    Yo2nz6 <= CDBGPWRUPACK;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Eq2nz6 <= 1'b0;
  else
    Eq2nz6 <= Aabdt6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Er2nz6 <= 1'b0;
  else
    Er2nz6 <= DBGEN;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hs2nz6 <= 1'b0;
  else
    Hs2nz6 <= Cbbdt6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Et2nz6 <= 1'b0;
  else
    Et2nz6 <= DBGEN;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Su2nz6 <= 1'b0;
  else
    Su2nz6 <= Bcbdt6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Aw2nz6 <= 1'b0;
  else
    Aw2nz6 <= I8o7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ny2nz6 <= 1'b0;
  else
    Ny2nz6 <= B8o7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    A13nz6 <= 1'b0;
  else
    A13nz6 <= U7o7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N33nz6 <= 1'b0;
  else
    N33nz6 <= N7o7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    A63nz6 <= 1'b0;
  else
    A63nz6 <= G7o7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N83nz6 <= 1'b0;
  else
    N83nz6 <= Z6o7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ab3nz6 <= 1'b0;
  else
    Ab3nz6 <= DBGRESTART;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cd3nz6 <= 1'b0;
  else
    Cd3nz6 <= 1'b1;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bf3nz6 <= 1'b0;
  else
    Bf3nz6 <= S6o7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Yg3nz6 <= 1'b0;
  else
    Yg3nz6 <= WICENREQ;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Xh3nz6 <= 1'b0;
  else
    Xh3nz6 <= CDBGPWRUPACK;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Vj3nz6 <= 1'b0;
  else
    Vj3nz6 <= Mp67v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ul3nz6 <= 1'b0;
  else
    Ul3nz6 <= 1'b1;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Un3nz6 <= 1'b0;
  else
    Un3nz6 <= NIDEN;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ip3nz6 <= 1'b0;
  else
    Ip3nz6 <= I977v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vq3nz6 <= 1'b0;
  else
    Vq3nz6 <= Fy67v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ms3nz6 <= 1'b0;
  else
    Ms3nz6 <= 1'b1;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Su3nz6 <= 1'b0;
  else
    Su3nz6 <= Tho7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mw3nz6 <= 1'b0;
  else
    Mw3nz6 <= L6o7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sx3nz6 <= 1'b0;
  else
    Sx3nz6 <= Fql8v6;

always @(posedge HCLK) T04nz6 <= Qny7v6;
always @(posedge HCLK) D34nz6 <= Etl8v6;
always @(posedge FCLK) B64nz6 <= Cel8v6;
always @(posedge FCLK) P84nz6 <= Vdl8v6;
always @(posedge FCLK) Ab4nz6 <= Odl8v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pd4nz6 <= 1'b0;
  else
    Pd4nz6 <= Adl8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jf4nz6 <= 1'b0;
  else
    Jf4nz6 <= Hdl8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jh4nz6 <= 1'b0;
  else
    Jh4nz6 <= Kmp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jj4nz6 <= 1'b0;
  else
    Jj4nz6 <= Kbl8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hl4nz6 <= 1'b0;
  else
    Hl4nz6 <= G9l8v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Un4nz6 <= 1'b0;
  else
    Un4nz6 <= U81nz6[1];

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Nq4nz6 <= 1'b0;
  else
    Nq4nz6 <= J1h7v6;

always @(posedge HCLK) Gt4nz6 <= Ltl8v6;
always @(posedge HCLK) Yv4nz6 <= Tks7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    My4nz6 <= 1'b0;
  else
    My4nz6 <= Loj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L15nz6 <= 1'b0;
  else
    L15nz6 <= F2p7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    R45nz6 <= 1'b0;
  else
    R45nz6 <= Tm48v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H65nz6 <= 1'b0;
  else
    H65nz6 <= Eoj8v6;

always @(posedge HCLK) G95nz6 <= P7p7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kc5nz6 <= 1'b0;
  else
    Kc5nz6 <= Fjl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jf5nz6 <= 1'b0;
  else
    Jf5nz6 <= Eaj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mi5nz6 <= 1'b0;
  else
    Mi5nz6 <= Fly7v6;

always @(posedge HCLK) Kl5nz6 <= Yky7v6;
always @(posedge HCLK) Ho5nz6 <= X0l8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qq5nz6 <= 1'b0;
  else
    Qq5nz6 <= Efl8v6;

always @(posedge FCLK) Rs5nz6 <= H1r7v6;
always @(posedge FCLK) Ou5nz6 <= Gyp7v6;
always @(posedge FCLK) Zw5nz6 <= Sxp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Oz5nz6 <= 1'b0;
  else
    Oz5nz6 <= Cpp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    O16nz6 <= 1'b0;
  else
    O16nz6 <= Ohp7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M36nz6 <= 1'b0;
  else
    M36nz6 <= Hrl8v6;

always @(posedge HCLK) N66nz6 <= Amy7v6;
always @(posedge HCLK) X86nz6 <= C0l8v6;
always @(posedge HCLK) Vb6nz6 <= Tys7v6;
always @(posedge HCLK) Pe6nz6 <= Mys7v6;
always @(posedge HCLK) Jh6nz6 <= Fys7v6;
always @(posedge HCLK) Dk6nz6 <= Yxs7v6;
always @(posedge HCLK) Ym6nz6 <= Rxs7v6;
always @(posedge HCLK) Tp6nz6 <= Kxs7v6;
always @(posedge HCLK) Os6nz6 <= Dxs7v6;
always @(posedge HCLK) Jv6nz6 <= Wws7v6;
always @(posedge HCLK) Ey6nz6 <= Pws7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z07nz6 <= 1'b0;
  else
    Z07nz6 <= Ggl8v6;

always @(posedge HCLK) A37nz6 <= Ngl8v6;
always @(posedge HCLK) P57nz6 <= Ivl8v6;
always @(posedge HCLK) H87nz6 <= E358v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z97nz6 <= 1'b0;
  else
    Z97nz6 <= Vl68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oc7nz6 <= 1'b0;
  else
    Oc7nz6 <= Jwh8v6;

always @(posedge HCLK) Af7nz6 <= Jr88v6;
always @(posedge HCLK) Qh7nz6 <= Egs7v6;
always @(posedge HCLK) Fk7nz6 <= Fey7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cn7nz6 <= 1'b0;
  else
    Cn7nz6 <= Vkl8v6;

always @(posedge HCLK) Cq7nz6 <= Mzy7v6;
always @(posedge HCLK) Ls7nz6 <= Vzk8v6;
always @(posedge HCLK) Jv7nz6 <= Be38v6;
always @(posedge HCLK) Dy7nz6 <= Ud38v6;
always @(posedge HCLK) X08nz6 <= Nd38v6;
always @(posedge HCLK) S38nz6 <= Gd38v6;
always @(posedge HCLK) N68nz6 <= Zc38v6;
always @(posedge HCLK) I98nz6 <= Sc38v6;
always @(posedge HCLK) Dc8nz6 <= Lc38v6;
always @(posedge HCLK) Ye8nz6 <= J0l8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Th8nz6 <= 1'b0;
  else
    Th8nz6 <= P3l8v6;

always @(posedge FCLK) Uj8nz6 <= V1r7v6;
always @(posedge FCLK) Rl8nz6 <= U5q7v6;
always @(posedge FCLK) Co8nz6 <= G5q7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rq8nz6 <= 1'b0;
  else
    Rq8nz6 <= Aop7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rs8nz6 <= 1'b0;
  else
    Rs8nz6 <= Sjp7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pu8nz6 <= 1'b0;
  else
    Pu8nz6 <= Tql8v6;

always @(posedge HCLK) Qx8nz6 <= Hmy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    A09nz6 <= 1'b0;
  else
    A09nz6 <= Sfl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X29nz6 <= 1'b0;
  else
    X29nz6 <= Mly7v6;

always @(posedge HCLK) R59nz6 <= Fdk8v6;
always @(posedge HCLK) P89nz6 <= Zpi8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lb9nz6 <= 1'b0;
  else
    Lb9nz6 <= Q4a7z6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Le9nz6 <= 1'b0;
  else
    Le9nz6 <= Ycs7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oh9nz6 <= 1'b0;
  else
    Oh9nz6 <= N098v6;

always @(posedge HCLK) Ik9nz6 <= Rky7v6;
always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gn9nz6 <= 1'b0;
  else
    Gn9nz6 <= Djk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fq9nz6 <= 1'b0;
  else
    Fq9nz6 <= Ask8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ct9nz6 <= 1'b0;
  else
    Ct9nz6 <= Mrk8v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Av9nz6 <= 1'b0;
  else
    Av9nz6 <= Ad78v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Zv9nz6 <= 1'b0;
  else
    Zv9nz6 <= Gv68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Zw9nz6 <= 1'b0;
  else
    Zw9nz6 <= Nv68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Zx9nz6 <= 1'b0;
  else
    Zx9nz6 <= Uv68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Zy9nz6 <= 1'b0;
  else
    Zy9nz6 <= Bw68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Zz9nz6 <= 1'b0;
  else
    Zz9nz6 <= Iw68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Z0anz6 <= 1'b0;
  else
    Z0anz6 <= Pw68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Z1anz6 <= 1'b0;
  else
    Z1anz6 <= Ww68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Z2anz6 <= 1'b0;
  else
    Z2anz6 <= Dx68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Z3anz6 <= 1'b0;
  else
    Z3anz6 <= Kx68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Z4anz6 <= 1'b0;
  else
    Z4anz6 <= Rx68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    A6anz6 <= 1'b0;
  else
    A6anz6 <= Yx68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    B7anz6 <= 1'b0;
  else
    B7anz6 <= Fy68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    C8anz6 <= 1'b0;
  else
    C8anz6 <= My68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    D9anz6 <= 1'b0;
  else
    D9anz6 <= Ty68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Eaanz6 <= 1'b0;
  else
    Eaanz6 <= Az68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Fbanz6 <= 1'b0;
  else
    Fbanz6 <= Hz68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Gcanz6 <= 1'b0;
  else
    Gcanz6 <= Oz68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Hdanz6 <= 1'b0;
  else
    Hdanz6 <= Vz68v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Ieanz6 <= 1'b0;
  else
    Ieanz6 <= C078v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Jfanz6 <= 1'b0;
  else
    Jfanz6 <= J078v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Kganz6 <= 1'b0;
  else
    Kganz6 <= Q078v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Lhanz6 <= 1'b0;
  else
    Lhanz6 <= X078v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Mianz6 <= 1'b0;
  else
    Mianz6 <= E178v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Njanz6 <= 1'b0;
  else
    Njanz6 <= L178v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Okanz6 <= 1'b0;
  else
    Okanz6 <= S178v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Planz6 <= 1'b0;
  else
    Planz6 <= Z178v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Qmanz6 <= 1'b0;
  else
    Qmanz6 <= G278v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Rnanz6 <= 1'b0;
  else
    Rnanz6 <= N278v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Soanz6 <= 1'b0;
  else
    Soanz6 <= U278v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Tpanz6 <= 1'b0;
  else
    Tpanz6 <= B378v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Uqanz6 <= 1'b0;
  else
    Uqanz6 <= I378v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Vranz6 <= 1'b0;
  else
    Vranz6 <= P378v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Wsanz6 <= 1'b0;
  else
    Wsanz6 <= W378v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Xtanz6 <= 1'b0;
  else
    Xtanz6 <= D478v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Yuanz6 <= 1'b0;
  else
    Yuanz6 <= K478v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Zvanz6 <= 1'b0;
  else
    Zvanz6 <= R478v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Axanz6 <= 1'b0;
  else
    Axanz6 <= Y478v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Byanz6 <= 1'b0;
  else
    Byanz6 <= F578v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Czanz6 <= 1'b0;
  else
    Czanz6 <= M578v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    D0bnz6 <= 1'b0;
  else
    D0bnz6 <= T578v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    E1bnz6 <= 1'b0;
  else
    E1bnz6 <= A678v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    F2bnz6 <= 1'b0;
  else
    F2bnz6 <= H678v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    G3bnz6 <= 1'b0;
  else
    G3bnz6 <= O678v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    H4bnz6 <= 1'b0;
  else
    H4bnz6 <= V678v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    I5bnz6 <= 1'b0;
  else
    I5bnz6 <= C778v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    J6bnz6 <= 1'b0;
  else
    J6bnz6 <= J778v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    K7bnz6 <= 1'b0;
  else
    K7bnz6 <= Q778v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    L8bnz6 <= 1'b0;
  else
    L8bnz6 <= X778v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    M9bnz6 <= 1'b0;
  else
    M9bnz6 <= E878v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Nabnz6 <= 1'b0;
  else
    Nabnz6 <= L878v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Obbnz6 <= 1'b0;
  else
    Obbnz6 <= S878v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Pcbnz6 <= 1'b0;
  else
    Pcbnz6 <= Z878v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Qdbnz6 <= 1'b0;
  else
    Qdbnz6 <= G978v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Rebnz6 <= 1'b0;
  else
    Rebnz6 <= N978v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Sfbnz6 <= 1'b0;
  else
    Sfbnz6 <= U978v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Tgbnz6 <= 1'b0;
  else
    Tgbnz6 <= Ba78v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Uhbnz6 <= 1'b0;
  else
    Uhbnz6 <= Ia78v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Vibnz6 <= 1'b0;
  else
    Vibnz6 <= Pa78v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Wjbnz6 <= 1'b0;
  else
    Wjbnz6 <= Wa78v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Xkbnz6 <= 1'b0;
  else
    Xkbnz6 <= Db78v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Ylbnz6 <= 1'b0;
  else
    Ylbnz6 <= Kb78v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Zmbnz6 <= 1'b0;
  else
    Zmbnz6 <= Rb78v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Aobnz6 <= 1'b0;
  else
    Aobnz6 <= Yb78v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Bpbnz6 <= 1'b0;
  else
    Bpbnz6 <= Fc78v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Cqbnz6 <= 1'b0;
  else
    Cqbnz6 <= Mc78v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Drbnz6 <= 1'b0;
  else
    Drbnz6 <= Tc78v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Dsbnz6 <= 1'b0;
  else
    Dsbnz6 <= Frk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Etbnz6 <= 1'b0;
  else
    Etbnz6 <= E6o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fwbnz6 <= 1'b0;
  else
    Fwbnz6 <= X5o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hzbnz6 <= 1'b0;
  else
    Hzbnz6 <= Q5o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    J2cnz6 <= 1'b0;
  else
    J2cnz6 <= J5o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    L5cnz6 <= 1'b0;
  else
    L5cnz6 <= C5o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    N8cnz6 <= 1'b0;
  else
    N8cnz6 <= V4o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pbcnz6 <= 1'b0;
  else
    Pbcnz6 <= O4o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Recnz6 <= 1'b0;
  else
    Recnz6 <= H4o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Thcnz6 <= 1'b0;
  else
    Thcnz6 <= A4o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vkcnz6 <= 1'b0;
  else
    Vkcnz6 <= T3o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xncnz6 <= 1'b0;
  else
    Xncnz6 <= M3o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zqcnz6 <= 1'b0;
  else
    Zqcnz6 <= F3o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bucnz6 <= 1'b0;
  else
    Bucnz6 <= Y2o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dxcnz6 <= 1'b0;
  else
    Dxcnz6 <= R2o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    F0dnz6 <= 1'b0;
  else
    F0dnz6 <= K2o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    H3dnz6 <= 1'b0;
  else
    H3dnz6 <= D2o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    J6dnz6 <= 1'b0;
  else
    J6dnz6 <= W1o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    L9dnz6 <= 1'b0;
  else
    L9dnz6 <= P1o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ncdnz6 <= 1'b0;
  else
    Ncdnz6 <= I1o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pfdnz6 <= 1'b0;
  else
    Pfdnz6 <= B1o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ridnz6 <= 1'b0;
  else
    Ridnz6 <= U0o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tldnz6 <= 1'b0;
  else
    Tldnz6 <= N0o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vodnz6 <= 1'b0;
  else
    Vodnz6 <= G0o7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xrdnz6 <= 1'b0;
  else
    Xrdnz6 <= Zzn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zudnz6 <= 1'b0;
  else
    Zudnz6 <= Szn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bydnz6 <= 1'b0;
  else
    Bydnz6 <= Lzn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    D1enz6 <= 1'b0;
  else
    D1enz6 <= Ezn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    F4enz6 <= 1'b0;
  else
    F4enz6 <= Xyn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    H7enz6 <= 1'b0;
  else
    H7enz6 <= Qyn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jaenz6 <= 1'b0;
  else
    Jaenz6 <= Jyn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ldenz6 <= 1'b0;
  else
    Ldenz6 <= Cyn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ngenz6 <= 1'b0;
  else
    Ngenz6 <= Vxn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pjenz6 <= 1'b0;
  else
    Pjenz6 <= Oxn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rmenz6 <= 1'b0;
  else
    Rmenz6 <= Hxn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tpenz6 <= 1'b0;
  else
    Tpenz6 <= Axn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vsenz6 <= 1'b0;
  else
    Vsenz6 <= Twn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xvenz6 <= 1'b0;
  else
    Xvenz6 <= Mwn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zyenz6 <= 1'b0;
  else
    Zyenz6 <= Fwn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    B2fnz6 <= 1'b0;
  else
    B2fnz6 <= Yvn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    D5fnz6 <= 1'b0;
  else
    D5fnz6 <= Rvn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    F8fnz6 <= 1'b0;
  else
    F8fnz6 <= Kvn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hbfnz6 <= 1'b0;
  else
    Hbfnz6 <= Dvn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jefnz6 <= 1'b0;
  else
    Jefnz6 <= Wun7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lhfnz6 <= 1'b0;
  else
    Lhfnz6 <= Pun7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nkfnz6 <= 1'b0;
  else
    Nkfnz6 <= Iun7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pnfnz6 <= 1'b0;
  else
    Pnfnz6 <= Bun7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rqfnz6 <= 1'b0;
  else
    Rqfnz6 <= Utn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ttfnz6 <= 1'b0;
  else
    Ttfnz6 <= Ntn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vwfnz6 <= 1'b0;
  else
    Vwfnz6 <= Gtn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xzfnz6 <= 1'b0;
  else
    Xzfnz6 <= Zsn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z2gnz6 <= 1'b0;
  else
    Z2gnz6 <= Ssn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    B6gnz6 <= 1'b0;
  else
    B6gnz6 <= Lsn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    D9gnz6 <= 1'b0;
  else
    D9gnz6 <= Esn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fcgnz6 <= 1'b0;
  else
    Fcgnz6 <= Xrn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hfgnz6 <= 1'b0;
  else
    Hfgnz6 <= Qrn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jignz6 <= 1'b0;
  else
    Jignz6 <= Jrn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Llgnz6 <= 1'b0;
  else
    Llgnz6 <= Crn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nognz6 <= 1'b0;
  else
    Nognz6 <= Vqn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Prgnz6 <= 1'b0;
  else
    Prgnz6 <= Oqn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rugnz6 <= 1'b0;
  else
    Rugnz6 <= Hqn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Txgnz6 <= 1'b0;
  else
    Txgnz6 <= Aqn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    V0hnz6 <= 1'b0;
  else
    V0hnz6 <= Tpn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    X3hnz6 <= 1'b0;
  else
    X3hnz6 <= Mpn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z6hnz6 <= 1'b0;
  else
    Z6hnz6 <= Fpn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bahnz6 <= 1'b0;
  else
    Bahnz6 <= Yon7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cdhnz6 <= 1'b0;
  else
    Cdhnz6 <= Ron7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dghnz6 <= 1'b0;
  else
    Dghnz6 <= Yqk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bjhnz6 <= 1'b0;
  else
    Bjhnz6 <= Oxfet6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Elhnz6 <= 1'b0;
  else
    Elhnz6 <= Qtfet6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cnhnz6 <= 1'b0;
  else
    Cnhnz6 <= Gpfet6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hphnz6 <= 1'b0;
  else
    Hphnz6 <= Svj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yrhnz6 <= 1'b0;
  else
    Yrhnz6 <= R1p7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tuhnz6 <= 1'b0;
  else
    Tuhnz6 <= Gzo7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zxhnz6 <= 1'b0;
  else
    Zxhnz6 <= R4l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pzhnz6 <= 1'b0;
  else
    Pzhnz6 <= Iqj8v6;

always @(posedge HCLK) O2inz6 <= L5p7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    S5inz6 <= 1'b0;
  else
    S5inz6 <= Ykj8v6;

always @(posedge HCLK) Q8inz6 <= M1i8v6;
always @(posedge HCLK) Vainz6 <= Kon7v6;
always @(posedge HCLK) Xdinz6 <= Don7v6;
always @(posedge HCLK) Zginz6 <= Wnn7v6;
always @(posedge HCLK) Bkinz6 <= Pnn7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dninz6 <= 1'b0;
  else
    Dninz6 <= D0i8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tpinz6 <= 1'b0;
  else
    Tpinz6 <= Wzh8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Osinz6 <= 1'b0;
  else
    Osinz6 <= W5a7z6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kvinz6 <= 1'b0;
  else
    Kvinz6 <= Z2k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Myinz6 <= 1'b0;
  else
    Myinz6 <= Id48v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O1jnz6 <= 1'b0;
  else
    O1jnz6 <= Pyx7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    N3jnz6 <= 1'b0;
  else
    N3jnz6 <= Znk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    S5jnz6 <= 1'b0;
  else
    S5jnz6 <= Ibk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Q7jnz6 <= 1'b0;
  else
    Q7jnz6 <= HALTED;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    P9jnz6 <= 1'b0;
  else
    P9jnz6 <= Z2c7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Objnz6 <= 1'b0;
  else
    Objnz6 <= HALTED;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qdjnz6 <= 1'b1;
  else
    Qdjnz6 <= Ddeet6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wfjnz6 <= 1'b0;
  else
    Wfjnz6 <= X8eet6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bijnz6 <= 1'b0;
  else
    Bijnz6 <= Ujx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fkjnz6 <= 1'b0;
  else
    Fkjnz6 <= Svc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gmjnz6 <= 1'b0;
  else
    Gmjnz6 <= Zwx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qojnz6 <= 1'b0;
  else
    Qojnz6 <= Tjl8v6;

always @(posedge HCLK) Qrjnz6 <= U638v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ztjnz6 <= 1'b0;
  else
    Ztjnz6 <= Ugl8v6;

always @(posedge FCLK) Fxjnz6 <= Hiv7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lzjnz6 <= 1'b0;
  else
    Lzjnz6 <= Iyq7v6;

always @(posedge FCLK) P2knz6 <= Uxq7v6;
always @(posedge FCLK) D5knz6 <= Lbq7v6;
always @(posedge FCLK) O7knz6 <= Lqp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Daknz6 <= 1'b0;
  else
    Daknz6 <= Eqp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dcknz6 <= 1'b0;
  else
    Dcknz6 <= Ial8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Beknz6 <= 1'b0;
  else
    Beknz6 <= Rpl8v6;

always @(posedge HCLK) Chknz6 <= K5z7v6;
always @(posedge HCLK) Mjknz6 <= Bjy7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kmknz6 <= 1'b0;
  else
    Kmknz6 <= Inn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qoknz6 <= 1'b0;
  else
    Qoknz6 <= Lrfet6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vqknz6 <= 1'b0;
  else
    Vqknz6 <= Ixj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mtknz6 <= 1'b0;
  else
    Mtknz6 <= Xp38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jwknz6 <= 1'b0;
  else
    Jwknz6 <= Zyo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pzknz6 <= 1'b1;
  else
    Pzknz6 <= Qsl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J2lnz6 <= 1'b0;
  else
    J2lnz6 <= Xuj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L5lnz6 <= 1'b0;
  else
    L5lnz6 <= Mjl8v6;

always @(posedge HCLK) L8lnz6 <= W3l8v6;
always @(posedge HCLK) Ualnz6 <= Wcy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rdlnz6 <= 1'b0;
  else
    Rdlnz6 <= Msj8v6;

always @(posedge HCLK) Pglnz6 <= T8i8v6;
always @(posedge HCLK) Uilnz6 <= Pbz7v6;
always @(posedge HCLK) Dllnz6 <= Tey7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Aolnz6 <= 1'b0;
  else
    Aolnz6 <= Jll8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Arlnz6 <= 1'b0;
  else
    Arlnz6 <= Uzo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fulnz6 <= 1'b0;
  else
    Fulnz6 <= Eq38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Exlnz6 <= 1'b0;
  else
    Exlnz6 <= Mkk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Azlnz6 <= 1'b0;
  else
    Azlnz6 <= Fuw7v6;

always @(posedge HCLK) A1mnz6 <= Mey7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X3mnz6 <= 1'b0;
  else
    X3mnz6 <= Cll8v6;

always @(posedge HCLK) X6mnz6 <= Wxy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    G9mnz6 <= 1'b0;
  else
    G9mnz6 <= Zfl8v6;

always @(posedge HCLK) Qbmnz6 <= Ycz7v6;
always @(posedge HCLK) Zdmnz6 <= Rdy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wgmnz6 <= 1'b0;
  else
    Wgmnz6 <= Hkl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wjmnz6 <= 1'b0;
  else
    Wjmnz6 <= Y1p7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cnmnz6 <= 1'b0;
  else
    Cnmnz6 <= Kil8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zpmnz6 <= 1'b0;
  else
    Zpmnz6 <= Ihl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wsmnz6 <= 1'b0;
  else
    Wsmnz6 <= Dil8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xvmnz6 <= 1'b0;
  else
    Xvmnz6 <= Phl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yymnz6 <= 1'b0;
  else
    Yymnz6 <= Whl8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Z1nnz6 <= 1'b0;
  else
    Z1nnz6 <= Bnn7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    X4nnz6 <= 1'b0;
  else
    X4nnz6 <= Umn7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    T7nnz6 <= 1'b0;
  else
    T7nnz6 <= Dsx7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    N9nnz6 <= 1'b1;
  else
    N9nnz6 <= Wrx7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gbnnz6 <= 1'b0;
  else
    Gbnnz6 <= M0r7v6;

always @(posedge FCLK) Wcnnz6 <= F0r7v6;
always @(posedge FCLK) Sennz6 <= Fup7v6;
always @(posedge FCLK) Dhnnz6 <= Rtp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Sjnnz6 <= 1'b0;
  else
    Sjnnz6 <= Tcl8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Plnnz6 <= 1'b0;
  else
    Plnnz6 <= Ybl8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mnnnz6 <= 1'b0;
  else
    Mnnnz6 <= Qip7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kpnnz6 <= 1'b0;
  else
    Kpnnz6 <= Arl8v6;

always @(posedge HCLK) Lsnnz6 <= Tyk8v6;
always @(posedge HCLK) Vunnz6 <= Kky7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Txnnz6 <= 1'b0;
  else
    Txnnz6 <= Z3y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vznnz6 <= 1'b0;
  else
    Vznnz6 <= Wol8v6;

always @(posedge HCLK) W2onz6 <= O0z7v6;
always @(posedge HCLK) G5onz6 <= Giy7v6;
always @(posedge HCLK) E8onz6 <= Zp48v6;
always @(posedge HCLK) U9onz6 <= Pu88v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nbonz6 <= 1'b0;
  else
    Nbonz6 <= Nak8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ceonz6 <= 1'b0;
  else
    Ceonz6 <= Jk88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sgonz6 <= 1'b0;
  else
    Sgonz6 <= Xms7v6;

always @(posedge HCLK) Ijonz6 <= Oes7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xlonz6 <= 1'b0;
  else
    Xlonz6 <= Mlj8v6;

always @(posedge HCLK) Voonz6 <= M9p7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yronz6 <= 1'b0;
  else
    Yronz6 <= Pqj8v6;

always @(posedge HCLK) Xuonz6 <= H2i8v6;
always @(posedge HCLK) Cxonz6 <= Myk8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mzonz6 <= 1'b0;
  else
    Mzonz6 <= I4a7z6;

always @(posedge HCLK) M2pnz6 <= Q1z7v6;
always @(posedge HCLK) V4pnz6 <= Kdy7v6;
always @(posedge FCLK) S7pnz6 <= K6r7v6;
always @(posedge FCLK) P9pnz6 <= Tmq7v6;
always @(posedge FCLK) Acpnz6 <= Tnp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pepnz6 <= 1'b0;
  else
    Pepnz6 <= Mnp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pgpnz6 <= 1'b0;
  else
    Pgpnz6 <= Ukp7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nipnz6 <= 1'b0;
  else
    Nipnz6 <= Mql8v6;

always @(posedge HCLK) Olpnz6 <= Omy7v6;
always @(posedge HCLK) Ynpnz6 <= Wjy7v6;
always @(posedge FCLK) Wqpnz6 <= Hy78v6;
always @(posedge FCLK) Etpnz6 <= Gxq7v6;
always @(posedge FCLK) Svpnz6 <= Ziq7v6;
always @(posedge FCLK) Dypnz6 <= Fnp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    S0qnz6 <= 1'b0;
  else
    S0qnz6 <= Ymp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    S2qnz6 <= 1'b0;
  else
    S2qnz6 <= Wlp7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q4qnz6 <= 1'b0;
  else
    Q4qnz6 <= Bol8v6;

always @(posedge HCLK) R7qnz6 <= C8z7v6;
always @(posedge HCLK) Baqnz6 <= Lhy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zcqnz6 <= 1'b0;
  else
    Zcqnz6 <= Wdx7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xfqnz6 <= 1'b0;
  else
    Xfqnz6 <= Pdx7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Viqnz6 <= 1'b0;
  else
    Viqnz6 <= Lgk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zkqnz6 <= 1'b0;
  else
    Zkqnz6 <= Jw38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ynqnz6 <= 1'b0;
  else
    Ynqnz6 <= Rjk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cqqnz6 <= 1'b0;
  else
    Cqqnz6 <= Sgk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Atqnz6 <= 1'b0;
  else
    Atqnz6 <= Oek8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Evqnz6 <= 1'b0;
  else
    Evqnz6 <= T8x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dyqnz6 <= 1'b0;
  else
    Dyqnz6 <= Jfk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    H0rnz6 <= 1'b0;
  else
    H0rnz6 <= Jww7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    G3rnz6 <= 1'b0;
  else
    G3rnz6 <= Hek8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K5rnz6 <= 1'b0;
  else
    K5rnz6 <= Pxj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O8rnz6 <= 1'b0;
  else
    O8rnz6 <= Ypl8v6;

always @(posedge HCLK) Pbrnz6 <= Y5z7v6;
always @(posedge HCLK) Zdrnz6 <= Ijy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xgrnz6 <= 1'b0;
  else
    Xgrnz6 <= B5y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yirnz6 <= 1'b0;
  else
    Yirnz6 <= Unl8v6;

always @(posedge HCLK) Zlrnz6 <= U3z7v6;
always @(posedge HCLK) Jornz6 <= Ehy7v6;
always @(posedge FCLK) Hrrnz6 <= Aiv7v6;
always @(posedge FCLK) Ntrnz6 <= Kgv7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tvrnz6 <= 1'b0;
  else
    Tvrnz6 <= Kpl8v6;

always @(posedge HCLK) Uyrnz6 <= Nwy7v6;
always @(posedge HCLK) E1snz6 <= Uiy7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    C4snz6 <= 1'b0;
  else
    C4snz6 <= X7l8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F6snz6 <= 1'b0;
  else
    F6snz6 <= Xle8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F8snz6 <= 1'b0;
  else
    F8snz6 <= Ulv7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hasnz6 <= 1'b1;
  else
    Hasnz6 <= Bik8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fcsnz6 <= 1'b0;
  else
    Fcsnz6 <= Axbdt6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jesnz6 <= 1'b0;
  else
    Jesnz6 <= Wxj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hhsnz6 <= 1'b0;
  else
    Hhsnz6 <= Kyj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kksnz6 <= 1'b0;
  else
    Kksnz6 <= Jsl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xmsnz6 <= 1'b0;
  else
    Xmsnz6 <= Dyj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ypsnz6 <= 1'b0;
  else
    Ypsnz6 <= Ril8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Etsnz6 <= 1'b0;
  else
    Etsnz6 <= Yl48v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ewsnz6 <= 1'b0;
  else
    Ewsnz6 <= Qnj8v6;

always @(posedge HCLK) Dzsnz6 <= D8p7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H2tnz6 <= 1'b0;
  else
    H2tnz6 <= Yrj8v6;

always @(posedge HCLK) G5tnz6 <= E4i8v6;
always @(posedge HCLK) M7tnz6 <= Yyy7v6;
always @(posedge HCLK) W9tnz6 <= Niy7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Uctnz6 <= 1'b1;
  else
    Uctnz6 <= Dp78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Oetnz6 <= 1'b0;
  else
    Oetnz6 <= Rhu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mgtnz6 <= 1'b0;
  else
    Mgtnz6 <= Iwk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kitnz6 <= 1'b0;
  else
    Kitnz6 <= Nmn7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jktnz6 <= 1'b0;
  else
    Jktnz6 <= Pwk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hmtnz6 <= 1'b0;
  else
    Hmtnz6 <= Kxk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fotnz6 <= 1'b0;
  else
    Fotnz6 <= Wwk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dqtnz6 <= 1'b0;
  else
    Dqtnz6 <= Dxk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bstnz6 <= 1'b0;
  else
    Bstnz6 <= Hzs7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wttnz6 <= 1'b0;
  else
    Wttnz6 <= Jur7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Uvtnz6 <= 1'b0;
  else
    Uvtnz6 <= Evr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Hytnz6 <= 1'b0;
  else
    Hytnz6 <= Ja1nz6[2];

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    A1unz6 <= 1'b0;
  else
    A1unz6 <= Fwg7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    T3unz6 <= 1'b0;
  else
    T3unz6 <= Xur7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    G6unz6 <= 1'b0;
  else
    G6unz6 <= Ja1nz6[1];

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Z8unz6 <= 1'b0;
  else
    Z8unz6 <= Qtg7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Sbunz6 <= 1'b0;
  else
    Sbunz6 <= Mzr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qdunz6 <= 1'b0;
  else
    Qdunz6 <= Q1s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ofunz6 <= 1'b0;
  else
    Ofunz6 <= Ixr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mhunz6 <= 1'b0;
  else
    Mhunz6 <= Lvr7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kjunz6 <= 1'b0;
  else
    Kjunz6 <= Qll8v6;

always @(posedge HCLK) Kmunz6 <= I4z7v6;
always @(posedge HCLK) Tounz6 <= Afy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qrunz6 <= 1'b0;
  else
    Qrunz6 <= T0y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Stunz6 <= 1'b0;
  else
    Stunz6 <= V7k8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uwunz6 <= 1'b0;
  else
    Uwunz6 <= Gmn7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vzunz6 <= 1'b0;
  else
    Vzunz6 <= Zln7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    W2vnz6 <= 1'b0;
  else
    W2vnz6 <= Xfk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    U5vnz6 <= 1'b0;
  else
    U5vnz6 <= Alk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y7vnz6 <= 1'b0;
  else
    Y7vnz6 <= Tkk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cavnz6 <= 1'b0;
  else
    Cavnz6 <= Ovfet6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ccvnz6 <= 1'b0;
  else
    Ccvnz6 <= Zvj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tevnz6 <= 1'b0;
  else
    Tevnz6 <= Lvj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Khvnz6 <= 1'b0;
  else
    Khvnz6 <= Evj8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pkvnz6 <= 1'b0;
  else
    Pkvnz6 <= Gwj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Smvnz6 <= 1'b0;
  else
    Smvnz6 <= Gok8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rovnz6 <= 1'b0;
  else
    Rovnz6 <= Fkk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Prvnz6 <= 1'b0;
  else
    Prvnz6 <= V6l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Stvnz6 <= 1'b0;
  else
    Stvnz6 <= Mmddt6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wvvnz6 <= 1'b0;
  else
    Wvvnz6 <= Quj8v6;

always @(posedge HCLK) Yyvnz6 <= Aez7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D1wnz6 <= 1'b0;
  else
    D1wnz6 <= Xel8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N3wnz6 <= 1'b0;
  else
    N3wnz6 <= Enk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O5wnz6 <= 1'b0;
  else
    O5wnz6 <= F0y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q7wnz6 <= 1'b0;
  else
    Q7wnz6 <= Iol8v6;

always @(posedge HCLK) Rawnz6 <= S2z7v6;
always @(posedge HCLK) Bdwnz6 <= Shy7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zfwnz6 <= 1'b0;
  else
    Zfwnz6 <= Drymz6[0];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fiwnz6 <= 1'b0;
  else
    Fiwnz6 <= Us77v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lkwnz6 <= 1'b0;
  else
    Lkwnz6 <= Eml8v6;

always @(posedge HCLK) Mnwnz6 <= W038v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Eqwnz6 <= 1'b0;
  else
    Eqwnz6 <= Z2z7v6;

always @(posedge HCLK) Oswnz6 <= Zvy7v6;
always @(posedge HCLK) Yuwnz6 <= Zhy7v6;
always @(posedge HCLK) Wxwnz6 <= Ks48v6;
always @(posedge HCLK) Mzwnz6 <= Vfy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K2xnz6 <= 1'b0;
  else
    K2xnz6 <= Lml8v6;

always @(posedge HCLK) L5xnz6 <= E2z7v6;
always @(posedge FCLK) V7xnz6 <= Lkv7v6;
always @(posedge FCLK) Baxnz6 <= Viv7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hcxnz6 <= 1'b0;
  else
    Hcxnz6 <= Zml8v6;

always @(posedge HCLK) Ifxnz6 <= Kyy7v6;
always @(posedge HCLK) Shxnz6 <= Jgy7v6;
always @(posedge FCLK) Qkxnz6 <= V948v6;
always @(posedge FCLK) Wmxnz6 <= Ca48v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cpxnz6 <= 1'b0;
  else
    Cpxnz6 <= Azk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Drxnz6 <= 1'b0;
  else
    Drxnz6 <= Rzx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ftxnz6 <= 1'b0;
  else
    Ftxnz6 <= Sml8v6;

always @(posedge HCLK) Gwxnz6 <= A0z7v6;
always @(posedge HCLK) Qyxnz6 <= Cgy7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    O1ynz6 <= 1'b0;
  else
    O1ynz6 <= Ql78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    L3ynz6 <= 1'b0;
  else
    L3ynz6 <= Mj78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    J5ynz6 <= 1'b0;
  else
    J5ynz6 <= Tj78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    E7ynz6 <= 1'b0;
  else
    E7ynz6 <= Sln7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Y8ynz6 <= 1'b0;
  else
    Y8ynz6 <= W3e7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ebynz6 <= 1'b0;
  else
    Ebynz6 <= Thg7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kdynz6 <= 1'b0;
  else
    Kdynz6 <= Lln7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gfynz6 <= 1'b0;
  else
    Gfynz6 <= Eln7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Chynz6 <= 1'b0;
  else
    Chynz6 <= Xkn7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yiynz6 <= 1'b1;
  else
    Yiynz6 <= Ijr7v6;

always @(posedge FCLK) Xkynz6 <= Bcr7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rmynz6 <= 1'b0;
  else
    Rmynz6 <= Ehr7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hoynz6 <= 1'b1;
  else
    Hoynz6 <= Ubr7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gqynz6 <= 1'b0;
  else
    Gqynz6 <= Qkn7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gsynz6 <= 1'b0;
  else
    Gsynz6 <= Jkn7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Guynz6 <= 1'b0;
  else
    Guynz6 <= Ckn7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gwynz6 <= 1'b0;
  else
    Gwynz6 <= Vjn7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gyynz6 <= 1'b1;
  else
    Gyynz6 <= Ojn7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    G0znz6 <= 1'b0;
  else
    G0znz6 <= Xvq7v6;

always @(posedge FCLK) Y2znz6 <= Qvq7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    J5znz6 <= 1'b0;
  else
    J5znz6 <= Jvq7v6;

always @(posedge FCLK) B8znz6 <= N5q7v6;
always @(posedge FCLK) Maznz6 <= Zxp7v6;
always @(posedge FCLK) Xcznz6 <= Ytp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ifznz6 <= 1'b0;
  else
    Ifznz6 <= Brq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Aiznz6 <= 1'b0;
  else
    Aiznz6 <= Uqq7v6;

always @(posedge FCLK) Skznz6 <= Ktp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dnznz6 <= 1'b1;
  else
    Dnznz6 <= Nqq7v6;

always @(posedge HCLK) Kpznz6 <= Qgy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Isznz6 <= 1'b0;
  else
    Isznz6 <= Gnl8v6;

always @(posedge HCLK) Jvznz6 <= E9z7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Txznz6 <= 1'b0;
  else
    Txznz6 <= Kex7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    R00oz6 <= 1'b0;
  else
    R00oz6 <= Qfk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    P30oz6 <= 1'b0;
  else
    P30oz6 <= Olk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T50oz6 <= 1'b0;
  else
    T50oz6 <= Pik8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T70oz6 <= 1'b0;
  else
    T70oz6 <= D4l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ba0oz6 <= 1'b0;
  else
    Ba0oz6 <= Ej38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ec0oz6 <= 1'b0;
  else
    Ec0oz6 <= S1l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ge0oz6 <= 1'b0;
  else
    Ge0oz6 <= Gk38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jg0oz6 <= 1'b0;
  else
    Jg0oz6 <= Wpk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ki0oz6 <= 1'b0;
  else
    Ki0oz6 <= H3adt6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ek0oz6 <= 1'b0;
  else
    Ek0oz6 <= H3adt6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Em0oz6 <= 1'b0;
  else
    Em0oz6 <= T5b7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Io0oz6 <= 1'b0;
  else
    Io0oz6 <= Wha7z6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Sq0oz6 <= 1'b0;
  else
    Sq0oz6 <= U7a7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qs0oz6 <= 1'b0;
  else
    Qs0oz6 <= Xm87v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wu0oz6 <= 1'b0;
  else
    Wu0oz6 <= Fj87v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xw0oz6 <= 1'b0;
  else
    Xw0oz6 <= Ih87v6;

always @(posedge HCLK) Yy0oz6 <= Dau7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    V01oz6 <= 1'b0;
  else
    V01oz6 <= N3s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Q21oz6 <= 1'b0;
  else
    Q21oz6 <= C1s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    O41oz6 <= 1'b0;
  else
    O41oz6 <= Yyr7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M61oz6 <= 1'b0;
  else
    M61oz6 <= L1l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O81oz6 <= 1'b0;
  else
    O81oz6 <= Zj38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ra1oz6 <= 1'b0;
  else
    Ra1oz6 <= E1l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Md1oz6 <= 1'b0;
  else
    Md1oz6 <= J1k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Eg1oz6 <= 1'b1;
  else
    Eg1oz6 <= H9i8v6;

always @(posedge FCLK) Ji1oz6 <= Ja48v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pk1oz6 <= 1'b0;
  else
    Pk1oz6 <= Otc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ln1oz6 <= 1'b0;
  else
    Ln1oz6 <= P648v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qp1oz6 <= 1'b0;
  else
    Qp1oz6 <= P0b7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Or1oz6 <= 1'b0;
  else
    Or1oz6 <= Mya7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zt1oz6 <= 1'b0;
  else
    Zt1oz6 <= Xco7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wv1oz6 <= 1'b0;
  else
    Wv1oz6 <= Ox67v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jx1oz6 <= 1'b0;
  else
    Jx1oz6 <= Uia7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Oz1oz6 <= 1'b0;
  else
    Oz1oz6 <= W387v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    H12oz6 <= 1'b0;
  else
    H12oz6 <= Nfu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    H32oz6 <= 1'b0;
  else
    H32oz6 <= Gfu7v6;

always @(posedge HCLK) H52oz6 <= O6t7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    E72oz6 <= 1'b0;
  else
    E72oz6 <= U3s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Z82oz6 <= 1'b0;
  else
    Z82oz6 <= J1s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xa2oz6 <= 1'b0;
  else
    Xa2oz6 <= Fzr7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vc2oz6 <= 1'b0;
  else
    Vc2oz6 <= Jmk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Df2oz6 <= 1'b0;
  else
    Df2oz6 <= Fzj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Eh2oz6 <= 1'b0;
  else
    Eh2oz6 <= Yyj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gj2oz6 <= 1'b0;
  else
    Gj2oz6 <= Ryj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lm2oz6 <= 1'b0;
  else
    Lm2oz6 <= Mti8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ip2oz6 <= 1'b0;
  else
    Ip2oz6 <= Saj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fs2oz6 <= 1'b0;
  else
    Fs2oz6 <= Laj8v6;

always @(posedge HCLK) Cv2oz6 <= Fc08v6;
always @(posedge HCLK) Sx2oz6 <= Rb08v6;
always @(posedge HCLK) J03oz6 <= O608v6;
always @(posedge HCLK) A33oz6 <= W308v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q53oz6 <= 1'b0;
  else
    Q53oz6 <= Qmk8v6;

always @(posedge HCLK) Z73oz6 <= Uaz7v6;
always @(posedge HCLK) Ja3oz6 <= Hfy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hd3oz6 <= 1'b0;
  else
    Hd3oz6 <= Kfa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tg3oz6 <= 1'b0;
  else
    Tg3oz6 <= Lxh8v6;

always @(posedge HCLK) Sj3oz6 <= Exh8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lm3oz6 <= 1'b0;
  else
    Lm3oz6 <= Nnl8v6;

always @(posedge HCLK) Mp3oz6 <= W4z7v6;
always @(posedge HCLK) Wr3oz6 <= Xgy7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Uu3oz6 <= 1'b0;
  else
    Uu3oz6 <= W288v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ww3oz6 <= 1'b0;
  else
    Ww3oz6 <= Vhw7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wy3oz6 <= 1'b0;
  else
    Wy3oz6 <= W8zmz6[0];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    A14oz6 <= 1'b0;
  else
    A14oz6 <= Vzymz6[0];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    J34oz6 <= 1'b0;
  else
    J34oz6 <= Vzymz6[1];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    S54oz6 <= 1'b0;
  else
    S54oz6 <= Vzymz6[2];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    B84oz6 <= 1'b0;
  else
    B84oz6 <= Vzymz6[3];

always @(posedge HCLK) Ka4oz6 <= Ocu7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hc4oz6 <= 1'b0;
  else
    Hc4oz6 <= S2s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ce4oz6 <= 1'b0;
  else
    Ce4oz6 <= H0s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ag4oz6 <= 1'b0;
  else
    Ag4oz6 <= Dyr7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yh4oz6 <= 1'b0;
  else
    Yh4oz6 <= Lvc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ak4oz6 <= 1'b0;
  else
    Ak4oz6 <= Sj38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dm4oz6 <= 1'b0;
  else
    Dm4oz6 <= V0k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vo4oz6 <= 1'b0;
  else
    Vo4oz6 <= Yil8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ds4oz6 <= 1'b0;
  else
    Ds4oz6 <= Vtj8v6;

always @(posedge HCLK) Gv4oz6 <= Fao7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ky4oz6 <= 1'b0;
  else
    Ky4oz6 <= Htj8v6;

always @(posedge HCLK) O15oz6 <= Ke48v6;
always @(posedge HCLK) R45oz6 <= Uos7v6;
always @(posedge HCLK) V75oz6 <= Mrs7v6;
always @(posedge HCLK) Za5oz6 <= Ei48v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ce5oz6 <= 1'b0;
  else
    Ce5oz6 <= Juj8v6;

always @(posedge HCLK) Fh5oz6 <= P8o7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jk5oz6 <= 1'b0;
  else
    Jk5oz6 <= Cuj8v6;

always @(posedge HCLK) Nn5oz6 <= De48v6;
always @(posedge HCLK) Qq5oz6 <= Nos7v6;
always @(posedge HCLK) Ut5oz6 <= Frs7v6;
always @(posedge HCLK) Yw5oz6 <= Xh48v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B06oz6 <= 1'b0;
  else
    B06oz6 <= Atj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    E36oz6 <= 1'b0;
  else
    E36oz6 <= Xnj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D66oz6 <= 1'b0;
  else
    D66oz6 <= Fti8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    A96oz6 <= 1'b0;
  else
    A96oz6 <= Hjn7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Db6oz6 <= 1'b0;
  else
    Db6oz6 <= Iyx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hd6oz6 <= 1'b0;
  else
    Hd6oz6 <= N2l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ig6oz6 <= 1'b0;
  else
    Ig6oz6 <= U2l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jj6oz6 <= 1'b0;
  else
    Jj6oz6 <= Iws7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mm6oz6 <= 1'b0;
  else
    Mm6oz6 <= Z1l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pp6oz6 <= 1'b0;
  else
    Pp6oz6 <= Quc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rr6oz6 <= 1'b0;
  else
    Rr6oz6 <= O7k8v6;

always @(posedge HCLK) Yt6oz6 <= Y408v6;
always @(posedge HCLK) Ow6oz6 <= Gz28v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fz6oz6 <= 1'b0;
  else
    Fz6oz6 <= V0z7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O17oz6 <= 1'b0;
  else
    O17oz6 <= Rsi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O47oz6 <= 1'b0;
  else
    O47oz6 <= Abo7v6;

always @(posedge HCLK) O77oz6 <= Lvy7v6;
always @(posedge HCLK) Ka7oz6 <= Gqi8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gd7oz6 <= 1'b0;
  else
    Gd7oz6 <= O0k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hf7oz6 <= 1'b0;
  else
    Hf7oz6 <= Csl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Li7oz6 <= 1'b0;
  else
    Li7oz6 <= Mao7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kl7oz6 <= 1'b0;
  else
    Kl7oz6 <= Lbi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    No7oz6 <= 1'b0;
  else
    No7oz6 <= U3d7z6[1];

always @(posedge HCLK) Pr7oz6 <= N6p7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tu7oz6 <= 1'b0;
  else
    Tu7oz6 <= Jgj8v6;

always @(posedge HCLK) Rx7oz6 <= Vap7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U08oz6 <= 1'b0;
  else
    U08oz6 <= Gpj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T38oz6 <= 1'b0;
  else
    T38oz6 <= Evc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V58oz6 <= 1'b0;
  else
    V58oz6 <= Xuc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X78oz6 <= 1'b0;
  else
    X78oz6 <= Lj38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Aa8oz6 <= 1'b0;
  else
    Aa8oz6 <= Q1k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sc8oz6 <= 1'b0;
  else
    Sc8oz6 <= J7l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sf8oz6 <= 1'b0;
  else
    Sf8oz6 <= J8k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ui8oz6 <= 1'b1;
  else
    Ui8oz6 <= C8k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xk8oz6 <= 1'b0;
  else
    Xk8oz6 <= Rzb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ko8oz6 <= 1'b0;
  else
    Ko8oz6 <= Ssnet6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hr8oz6 <= 1'b0;
  else
    Hr8oz6 <= Nt88v6;

always @(posedge HCLK) Vt8oz6 <= Wis7v6;
always @(posedge HCLK) Jw8oz6 <= Zi48v6;
always @(posedge HCLK) Mz8oz6 <= Gj48v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P29oz6 <= 1'b0;
  else
    P29oz6 <= Wqj8v6;

always @(posedge HCLK) O59oz6 <= X4p7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    S89oz6 <= 1'b0;
  else
    S89oz6 <= Tlj8v6;

always @(posedge HCLK) Qb9oz6 <= Y0i8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vd9oz6 <= 1'b0;
  else
    Vd9oz6 <= C1k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ng9oz6 <= 1'b0;
  else
    Ng9oz6 <= X1k8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qj9oz6 <= 1'b0;
  else
    Qj9oz6 <= Ppk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ql9oz6 <= 1'b0;
  else
    Ql9oz6 <= Nw97v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Nn9oz6 <= 1'b0;
  else
    Nn9oz6 <= Yk87v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Up9oz6 <= 1'b0;
  else
    Up9oz6 <= Zz97v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zr9oz6 <= 1'b0;
  else
    Zr9oz6 <= T1zmz6[7];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gu9oz6 <= 1'b1;
  else
    Gu9oz6 <= Rxk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gw9oz6 <= 1'b0;
  else
    Gw9oz6 <= Bwk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gy9oz6 <= 1'b0;
  else
    Gy9oz6 <= Uvk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    G0aoz6 <= 1'b0;
  else
    G0aoz6 <= Zuk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    G2aoz6 <= 1'b0;
  else
    G2aoz6 <= L2s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    B4aoz6 <= 1'b0;
  else
    B4aoz6 <= A0s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Z5aoz6 <= 1'b0;
  else
    Z5aoz6 <= Wxr7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X7aoz6 <= 1'b0;
  else
    X7aoz6 <= H0k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z9aoz6 <= 1'b0;
  else
    Z9aoz6 <= M0y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bcaoz6 <= 1'b0;
  else
    Bcaoz6 <= Cuc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xeaoz6 <= 1'b0;
  else
    Xeaoz6 <= D748v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Chaoz6 <= 1'b0;
  else
    Chaoz6 <= Uy38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bkaoz6 <= 1'b0;
  else
    Bkaoz6 <= Ny38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Anaoz6 <= 1'b0;
  else
    Anaoz6 <= Msc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wpaoz6 <= 1'b0;
  else
    Wpaoz6 <= Aek8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bsaoz6 <= 1'b0;
  else
    Bsaoz6 <= Cww7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Avaoz6 <= 1'b0;
  else
    Avaoz6 <= Vvw7v6;

always @(posedge HCLK) Zxaoz6 <= B4s7v6;
always @(posedge HCLK) R0boz6 <= Qfs7v6;
always @(posedge HCLK) G3boz6 <= Bps7v6;
always @(posedge HCLK) K6boz6 <= Ips7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O9boz6 <= 1'b0;
  else
    O9boz6 <= Jnj8v6;

always @(posedge HCLK) Ncboz6 <= K8p7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rfboz6 <= 1'b0;
  else
    Rfboz6 <= Rrj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qiboz6 <= 1'b0;
  else
    Qiboz6 <= K6j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Plboz6 <= 1'b0;
  else
    Plboz6 <= U798v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Foboz6 <= 1'b1;
  else
    Foboz6 <= I898v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zqboz6 <= 1'b0;
  else
    Zqboz6 <= Ysi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qtboz6 <= 1'b0;
  else
    Qtboz6 <= Bxj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jwboz6 <= 1'b0;
  else
    Jwboz6 <= Rv88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wyboz6 <= 1'b0;
  else
    Wyboz6 <= Sb48v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y1coz6 <= 1'b0;
  else
    Y1coz6 <= Ytw7v6;

always @(posedge HCLK) Y3coz6 <= Aio7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Q6coz6 <= 1'b0;
  else
    Q6coz6 <= Buf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    L8coz6 <= 1'b0;
  else
    L8coz6 <= F9h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Eacoz6 <= 1'b0;
  else
    Eacoz6 <= Y8h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Xbcoz6 <= 1'b0;
  else
    Xbcoz6 <= R8h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Qdcoz6 <= 1'b0;
  else
    Qdcoz6 <= K8h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Jfcoz6 <= 1'b0;
  else
    Jfcoz6 <= D8h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Chcoz6 <= 1'b0;
  else
    Chcoz6 <= W7h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Vicoz6 <= 1'b0;
  else
    Vicoz6 <= P7h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Okcoz6 <= 1'b0;
  else
    Okcoz6 <= I7h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Hmcoz6 <= 1'b0;
  else
    Hmcoz6 <= B7h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Aocoz6 <= 1'b0;
  else
    Aocoz6 <= Fpf8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cqcoz6 <= 1'b0;
  else
    Cqcoz6 <= Eqh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Xrcoz6 <= 1'b0;
  else
    Xrcoz6 <= Jqg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Aucoz6 <= 1'b0;
  else
    Aucoz6 <= Ajn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Pvcoz6 <= 1'b0;
  else
    Pvcoz6 <= Rfh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Fxcoz6 <= 1'b0;
  else
    Fxcoz6 <= Kfh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Vycoz6 <= 1'b0;
  else
    Vycoz6 <= Dfh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    J0doz6 <= 1'b0;
  else
    J0doz6 <= Jv47v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    X1doz6 <= 1'b0;
  else
    X1doz6 <= Weh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    T3doz6 <= 1'b0;
  else
    T3doz6 <= Peh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    P5doz6 <= 1'b0;
  else
    P5doz6 <= Ieh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    L7doz6 <= 1'b0;
  else
    L7doz6 <= Beh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    H9doz6 <= 1'b0;
  else
    H9doz6 <= Udh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Dbdoz6 <= 1'b0;
  else
    Dbdoz6 <= Ndh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Zcdoz6 <= 1'b0;
  else
    Zcdoz6 <= Ech8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Vedoz6 <= 1'b0;
  else
    Vedoz6 <= Sch8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Rgdoz6 <= 1'b0;
  else
    Rgdoz6 <= Zch8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Nidoz6 <= 1'b0;
  else
    Nidoz6 <= Gdh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Jkdoz6 <= 1'b0;
  else
    Jkdoz6 <= Lch8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Fmdoz6 <= 1'b0;
  else
    Fmdoz6 <= Xbh8v6;

always @(posedge SWCLKTCK or negedge nTRST)
  if(~nTRST)
    Bodoz6 <= 1'b1;
  else
    Bodoz6 <= Z3ymz6[2];

always @(posedge SWCLKTCK or negedge nTRST)
  if(~nTRST)
    Updoz6 <= 1'b1;
  else
    Updoz6 <= Z3ymz6[0];

always @(posedge SWCLKTCK or negedge nTRST)
  if(~nTRST)
    Nrdoz6 <= 1'b1;
  else
    Nrdoz6 <= Z3ymz6[3];

always @(posedge SWCLKTCK or negedge nTRST)
  if(~nTRST)
    Gtdoz6 <= 1'b1;
  else
    Gtdoz6 <= Z3ymz6[1];

always @(posedge C3a7z6 or negedge Sz9dt6)
  if(~Sz9dt6)
    Zudoz6 <= 1'b0;
  else
    Zudoz6 <= D567v6;

always @(posedge SWCLKTCK or negedge nTRST)
  if(~nTRST)
    Nwdoz6 <= 1'b0;
  else
    Nwdoz6 <= Vah8v6;

always @(posedge SWCLKTCK or negedge nTRST)
  if(~nTRST)
    Fydoz6 <= 1'b0;
  else
    Fydoz6 <= Cbh8v6;

always @(posedge SWCLKTCK or negedge nTRST)
  if(~nTRST)
    Xzdoz6 <= 1'b0;
  else
    Xzdoz6 <= Qbh8v6;

always @(posedge SWCLKTCK or negedge nTRST)
  if(~nTRST)
    P1eoz6 <= 1'b0;
  else
    P1eoz6 <= Jbh8v6;

always @(posedge SWCLKTCK or negedge nTRST)
  if(~nTRST)
    H3eoz6 <= 1'b0;
  else
    H3eoz6 <= Oah8v6;

always @(posedge SWCLKTCK or negedge nTRST)
  if(~nTRST)
    Y4eoz6 <= 1'b1;
  else
    Y4eoz6 <= Hah8v6;

always @(posedge SWCLKTCK or negedge nTRST)
  if(~nTRST)
    P6eoz6 <= 1'b1;
  else
    P6eoz6 <= Aah8v6;

always @(posedge SWCLKTCK or negedge nTRST)
  if(~nTRST)
    G8eoz6 <= 1'b1;
  else
    G8eoz6 <= T9h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    X9eoz6 <= 1'b0;
  else
    X9eoz6 <= Pmg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Nbeoz6 <= 1'b0;
  else
    Nbeoz6 <= Img8v6;

always @(posedge SWCLKTCK) Edeoz6 <= Ymh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Veeoz6 <= 1'b0;
  else
    Veeoz6 <= Itg8v6;

always @(posedge FCLK) Ngeoz6 <= Fag8v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Djeoz6 <= 1'b0;
  else
    Djeoz6 <= H4g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ykeoz6 <= 1'b0;
  else
    Ykeoz6 <= C4h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Rmeoz6 <= 1'b0;
  else
    Rmeoz6 <= V3h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Koeoz6 <= 1'b0;
  else
    Koeoz6 <= O3h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Dqeoz6 <= 1'b0;
  else
    Dqeoz6 <= H3h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Wreoz6 <= 1'b0;
  else
    Wreoz6 <= A3h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Pteoz6 <= 1'b0;
  else
    Pteoz6 <= T2h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Hveoz6 <= 1'b0;
  else
    Hveoz6 <= M2h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Zweoz6 <= 1'b0;
  else
    Zweoz6 <= F2h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ryeoz6 <= 1'b0;
  else
    Ryeoz6 <= Rof8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    I0foz6 <= 1'b0;
  else
    I0foz6 <= Tin7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    M2foz6 <= 1'b0;
  else
    M2foz6 <= Min7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Q4foz6 <= 1'b0;
  else
    Q4foz6 <= Fin7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    U6foz6 <= 1'b0;
  else
    U6foz6 <= Yhn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Y8foz6 <= 1'b0;
  else
    Y8foz6 <= Rhn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Cbfoz6 <= 1'b0;
  else
    Cbfoz6 <= Khn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Gdfoz6 <= 1'b0;
  else
    Gdfoz6 <= Dhn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Lffoz6 <= 1'b0;
  else
    Lffoz6 <= Wgn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Qhfoz6 <= 1'b0;
  else
    Qhfoz6 <= Pgn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Vjfoz6 <= 1'b0;
  else
    Vjfoz6 <= Ign7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Amfoz6 <= 1'b0;
  else
    Amfoz6 <= Bgn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Fofoz6 <= 1'b0;
  else
    Fofoz6 <= Ufn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Kqfoz6 <= 1'b0;
  else
    Kqfoz6 <= Nfn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Psfoz6 <= 1'b0;
  else
    Psfoz6 <= Gfn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Uufoz6 <= 1'b0;
  else
    Uufoz6 <= Zen7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Zwfoz6 <= 1'b0;
  else
    Zwfoz6 <= Sen7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ezfoz6 <= 1'b0;
  else
    Ezfoz6 <= Len7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    J1goz6 <= 1'b0;
  else
    J1goz6 <= Een7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    V2goz6 <= 1'b0;
  else
    V2goz6 <= Esf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    K4goz6 <= 1'b0;
  else
    K4goz6 <= Oa67v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    A6goz6 <= 1'b0;
  else
    A6goz6 <= Xdn7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    X7goz6 <= 1'b0;
  else
    X7goz6 <= Qdn7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    V9goz6 <= 1'b0;
  else
    V9goz6 <= Jdn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Nbgoz6 <= 1'b0;
  else
    Nbgoz6 <= Up47v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Jdgoz6 <= 1'b0;
  else
    Jdgoz6 <= Un67v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Gfgoz6 <= 1'b0;
  else
    Gfgoz6 <= Cdn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Sggoz6 <= 1'b0;
  else
    Sggoz6 <= Vcn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ligoz6 <= 1'b0;
  else
    Ligoz6 <= Ocn7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ckgoz6 <= 1'b0;
  else
    Ckgoz6 <= Xrf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Rlgoz6 <= 1'b0;
  else
    Rlgoz6 <= G967v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jngoz6 <= 1'b0;
  else
    Jngoz6 <= Hcn7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ipgoz6 <= 1'b0;
  else
    Ipgoz6 <= Acn7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Irgoz6 <= 1'b0;
  else
    Irgoz6 <= Xph8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ctgoz6 <= 1'b0;
  else
    Ctgoz6 <= Cqg8v6;

always @(posedge SWCLKTCK) Evgoz6 <= Plh8v6;
always @(posedge SWCLKTCK) Wwgoz6 <= Wlh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Oygoz6 <= 1'b0;
  else
    Oygoz6 <= Fog8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    P0hoz6 <= 1'b0;
  else
    P0hoz6 <= Bvl8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    A2hoz6 <= 1'b0;
  else
    A2hoz6 <= Tuh8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    L3hoz6 <= 1'b0;
  else
    L3hoz6 <= Tbn7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Z5hoz6 <= 1'b0;
  else
    Z5hoz6 <= Dth8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    P8hoz6 <= 1'b0;
  else
    P8hoz6 <= Wsh8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Abhoz6 <= 1'b0;
  else
    Abhoz6 <= Vvh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Uchoz6 <= 1'b0;
  else
    Uchoz6 <= Voh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Jehoz6 <= 1'b0;
  else
    Jehoz6 <= Btg8v6;

always @(posedge SWCLKTCK) Wfhoz6 <= Hvh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ohhoz6 <= 1'b0;
  else
    Ohhoz6 <= Avh8v6;

always @(posedge SWCLKTCK) Cjhoz6 <= Tgh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ukhoz6 <= 1'b0;
  else
    Ukhoz6 <= Kug8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Imhoz6 <= 1'b0;
  else
    Imhoz6 <= Kng8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Dohoz6 <= 1'b0;
  else
    Dohoz6 <= O667v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Sphoz6 <= 1'b0;
  else
    Sphoz6 <= R1adt6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wqhoz6 <= 1'b0;
  else
    Wqhoz6 <= A9bdt6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Urhoz6 <= 1'b0;
  else
    Urhoz6 <= R1adt6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Sthoz6 <= 1'b0;
  else
    Sthoz6 <= Gr67v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Rvhoz6 <= 1'b0;
  else
    Rvhoz6 <= Gul8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Kxhoz6 <= 1'b0;
  else
    Kxhoz6 <= Mbn7v6;

always @(posedge FCLK) Pzhoz6 <= Ztl8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F2ioz6 <= 1'b0;
  else
    F2ioz6 <= Fbn7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    X4ioz6 <= 1'b0;
  else
    X4ioz6 <= I9f8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    W7ioz6 <= 1'b0;
  else
    W7ioz6 <= Bkx7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Faioz6 <= 1'b0;
  else
    Faioz6 <= Yan7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mcioz6 <= 1'b0;
  else
    Mcioz6 <= Y5k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Veioz6 <= 1'b0;
  else
    Veioz6 <= K5k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xhioz6 <= 1'b0;
  else
    Xhioz6 <= D5k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xkioz6 <= 1'b0;
  else
    Xkioz6 <= Pkx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xnioz6 <= 1'b0;
  else
    Xnioz6 <= Bhl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Arioz6 <= 1'b0;
  else
    Arioz6 <= B4k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Utioz6 <= 1'b0;
  else
    Utioz6 <= I4k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Twioz6 <= 1'b0;
  else
    Twioz6 <= N3k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pzioz6 <= 1'b0;
  else
    Pzioz6 <= G3k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L2joz6 <= 1'b0;
  else
    L2joz6 <= Uok8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N5joz6 <= 1'b0;
  else
    N5joz6 <= R5k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F8joz6 <= 1'b0;
  else
    F8joz6 <= Jvi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fbjoz6 <= 1'b0;
  else
    Fbjoz6 <= Ran7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jdjoz6 <= 1'b0;
  else
    Jdjoz6 <= Yrc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cgjoz6 <= 1'b0;
  else
    Cgjoz6 <= Snk8v6;

always @(posedge HCLK) Eijoz6 <= Z538v6;
always @(posedge HCLK) Wkjoz6 <= B038v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nnjoz6 <= 1'b0;
  else
    Nnjoz6 <= Tdk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wpjoz6 <= 1'b0;
  else
    Wpjoz6 <= Kan7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yrjoz6 <= 1'b0;
  else
    Yrjoz6 <= E2k8v6;

always @(posedge HCLK) Yujoz6 <= Xny7v6;
always @(posedge HCLK) Fxjoz6 <= Tdz7v6;
always @(posedge HCLK) Lzjoz6 <= B738v6;
always @(posedge HCLK) R1koz6 <= Mdz7v6;
always @(posedge HCLK) X3koz6 <= Fdz7v6;
always @(posedge HCLK) D6koz6 <= Rcz7v6;
always @(posedge HCLK) J8koz6 <= Kcz7v6;
always @(posedge HCLK) Pakoz6 <= Dcz7v6;
always @(posedge HCLK) Vckoz6 <= Wbz7v6;
always @(posedge HCLK) Bfkoz6 <= Ibz7v6;
always @(posedge HCLK) Hhkoz6 <= Bbz7v6;
always @(posedge HCLK) Ojkoz6 <= Naz7v6;
always @(posedge HCLK) Vlkoz6 <= Gaz7v6;
always @(posedge HCLK) Cokoz6 <= Z9z7v6;
always @(posedge HCLK) Jqkoz6 <= S9z7v6;
always @(posedge HCLK) Qskoz6 <= L9z7v6;
always @(posedge HCLK) Xukoz6 <= X8z7v6;
always @(posedge HCLK) Exkoz6 <= Q8z7v6;
always @(posedge HCLK) Lzkoz6 <= J8z7v6;
always @(posedge HCLK) S1loz6 <= V7z7v6;
always @(posedge HCLK) Z3loz6 <= O7z7v6;
always @(posedge HCLK) G6loz6 <= H7z7v6;
always @(posedge HCLK) N8loz6 <= A7z7v6;
always @(posedge HCLK) Ualoz6 <= T6z7v6;
always @(posedge HCLK) Bdloz6 <= M6z7v6;
always @(posedge HCLK) Ifloz6 <= F6z7v6;
always @(posedge HCLK) Phloz6 <= Gpy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wjloz6 <= 1'b0;
  else
    Wjloz6 <= W738v6;

always @(posedge HCLK) Gmloz6 <= Pjy7v6;
always @(posedge HCLK) Eploz6 <= Hls7v6;
always @(posedge HCLK) Srloz6 <= Ff48v6;
always @(posedge HCLK) Vuloz6 <= Mf48v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yxloz6 <= 1'b0;
  else
    Yxloz6 <= Zoj8v6;

always @(posedge HCLK) X0moz6 <= U6p7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B4moz6 <= 1'b0;
  else
    B4moz6 <= Cgj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z6moz6 <= 1'b0;
  else
    Z6moz6 <= Tti8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W9moz6 <= 1'b0;
  else
    W9moz6 <= A8j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tcmoz6 <= 1'b0;
  else
    Tcmoz6 <= Kqk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ufmoz6 <= 1'b0;
  else
    Ufmoz6 <= Hjf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dimoz6 <= 1'b0;
  else
    Dimoz6 <= Dan7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kkmoz6 <= 1'b0;
  else
    Kkmoz6 <= W9n7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mmmoz6 <= 1'b0;
  else
    Mmmoz6 <= V0d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gpmoz6 <= 1'b0;
  else
    Gpmoz6 <= P9n7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Krmoz6 <= 1'b0;
  else
    Krmoz6 <= I9n7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ptmoz6 <= 1'b1;
  else
    Ptmoz6 <= Vcf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tvmoz6 <= 1'b0;
  else
    Tvmoz6 <= Ocf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wxmoz6 <= 1'b0;
  else
    Wxmoz6 <= L9k8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    J0noz6 <= 1'b0;
  else
    J0noz6 <= B9n7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    W2noz6 <= 1'b1;
  else
    W2noz6 <= U8n7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    G5noz6 <= 1'b0;
  else
    G5noz6 <= Hpg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Y6noz6 <= 1'b0;
  else
    Y6noz6 <= Wmg8v6;

always @(posedge SWCLKTCK) N8noz6 <= Tnh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Eanoz6 <= 1'b0;
  else
    Eanoz6 <= Dug8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wbnoz6 <= 1'b0;
  else
    Wbnoz6 <= Yth8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Menoz6 <= 1'b0;
  else
    Menoz6 <= N8n7v6;

always @(posedge HCLK) Dhnoz6 <= Hnx7v6;
always @(posedge HCLK) Vjnoz6 <= Sgs7v6;
always @(posedge HCLK) Kmnoz6 <= Zus7v6;
always @(posedge HCLK) Opnoz6 <= Gvs7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ssnoz6 <= 1'b0;
  else
    Ssnoz6 <= Vfj8v6;

always @(posedge HCLK) Qvnoz6 <= Jbp7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tynoz6 <= 1'b0;
  else
    Tynoz6 <= Soj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    S1ooz6 <= 1'b0;
  else
    S1ooz6 <= Pdi8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    S3ooz6 <= 1'b0;
  else
    S3ooz6 <= Trk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R5ooz6 <= 1'b0;
  else
    R5ooz6 <= Vrl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O8ooz6 <= 1'b0;
  else
    O8ooz6 <= Wcj8v6;

always @(posedge HCLK) Kbooz6 <= Xwh8v6;
always @(posedge HCLK) Deooz6 <= Xfs7v6;
always @(posedge HCLK) Sgooz6 <= Xbp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kjooz6 <= 1'b0;
  else
    Kjooz6 <= Puf8v6;

always @(posedge SWCLKTCK) Flooz6 <= Ahh8v6;
always @(posedge SWCLKTCK) Xmooz6 <= Hhh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Poooz6 <= 1'b0;
  else
    Poooz6 <= Yug8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Dqooz6 <= 1'b0;
  else
    Dqooz6 <= Rng8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Yrooz6 <= 1'b0;
  else
    Yrooz6 <= Bmg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ltooz6 <= 1'b0;
  else
    Ltooz6 <= Jph8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Yuooz6 <= 1'b0;
  else
    Yuooz6 <= Zkg8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Twooz6 <= 1'b0;
  else
    Twooz6 <= Zsf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Nyooz6 <= 1'b0;
  else
    Nyooz6 <= Ssf8v6;

always @(posedge SWCLKTCK) E0poz6 <= Mgh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    V1poz6 <= 1'b0;
  else
    V1poz6 <= Dng8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    O3poz6 <= 1'b0;
  else
    O3poz6 <= Uzg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    C5poz6 <= 1'b0;
  else
    C5poz6 <= Hwg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    U6poz6 <= 1'b0;
  else
    U6poz6 <= Iuf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    M8poz6 <= 1'b0;
  else
    M8poz6 <= A4g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Eapoz6 <= 1'b0;
  else
    Eapoz6 <= Utf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Wbpoz6 <= 1'b0;
  else
    Wbpoz6 <= S6g8v6;

always @(posedge SWCLKTCK) Ndpoz6 <= Fnh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Efpoz6 <= 1'b0;
  else
    Efpoz6 <= Ptg8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wgpoz6 <= 1'b0;
  else
    Wgpoz6 <= Kth8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mjpoz6 <= 1'b0;
  else
    Mjpoz6 <= G8n7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zlpoz6 <= 1'b0;
  else
    Zlpoz6 <= E9k8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Nopoz6 <= 1'b0;
  else
    Nopoz6 <= Blzet6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Drpoz6 <= 1'b0;
  else
    Drpoz6 <= T21ft6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ntpoz6 <= 1'b0;
  else
    Ntpoz6 <= Hgzet6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fwpoz6 <= 1'b0;
  else
    Fwpoz6 <= Hgzet6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yypoz6 <= 1'b0;
  else
    Yypoz6 <= F51ft6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    L1qoz6 <= 1'b0;
  else
    L1qoz6 <= Z7n7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    A4qoz6 <= 1'b0;
  else
    A4qoz6 <= S7n7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    S6qoz6 <= 1'b0;
  else
    S6qoz6 <= L7n7v6;

always @(posedge HCLK) J9qoz6 <= Irx7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bcqoz6 <= 1'b0;
  else
    Bcqoz6 <= R9g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Vdqoz6 <= 1'b0;
  else
    Vdqoz6 <= K9g8v6;

always @(posedge SWCLKTCK) Mfqoz6 <= Ooh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Dhqoz6 <= 1'b0;
  else
    Dhqoz6 <= E7n7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fjqoz6 <= 1'b0;
  else
    Fjqoz6 <= Sdg8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zlqoz6 <= 1'b0;
  else
    Zlqoz6 <= X6n7v6;

always @(posedge FCLK) Qoqoz6 <= Mag8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Grqoz6 <= 1'b0;
  else
    Grqoz6 <= Q6n7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ytqoz6 <= 1'b0;
  else
    Ytqoz6 <= V4g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Tvqoz6 <= 1'b0;
  else
    Tvqoz6 <= O4g8v6;

always @(posedge SWCLKTCK) Lxqoz6 <= Dmh8v6;
always @(posedge SWCLKTCK) Dzqoz6 <= Kmh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    U0roz6 <= 1'b0;
  else
    U0roz6 <= Yfh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    K2roz6 <= 1'b0;
  else
    K2roz6 <= Gzg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Y3roz6 <= 1'b0;
  else
    Y3roz6 <= Nzg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    M5roz6 <= 1'b0;
  else
    M5roz6 <= Zyg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    A7roz6 <= 1'b0;
  else
    A7roz6 <= B0h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    O8roz6 <= 1'b0;
  else
    O8roz6 <= Jxg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Earoz6 <= 1'b0;
  else
    Earoz6 <= Cxg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ubroz6 <= 1'b1;
  else
    Ubroz6 <= Nlg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Pdroz6 <= 1'b0;
  else
    Pdroz6 <= J6n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Bfroz6 <= 1'b0;
  else
    Bfroz6 <= C6n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ogroz6 <= 1'b1;
  else
    Ogroz6 <= Owg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Hiroz6 <= 1'b0;
  else
    Hiroz6 <= V5n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ujroz6 <= 1'b0;
  else
    Ujroz6 <= O5n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Wlroz6 <= 1'b0;
  else
    Wlroz6 <= H5n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ynroz6 <= 1'b0;
  else
    Ynroz6 <= A5n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Aqroz6 <= 1'b0;
  else
    Aqroz6 <= T4n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Csroz6 <= 1'b0;
  else
    Csroz6 <= M4n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Furoz6 <= 1'b0;
  else
    Furoz6 <= F4n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Iwroz6 <= 1'b0;
  else
    Iwroz6 <= Y3n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Lyroz6 <= 1'b0;
  else
    Lyroz6 <= R3n7v6;

always @(posedge FCLK) O0soz6 <= Neg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    E3soz6 <= 1'b0;
  else
    E3soz6 <= K3n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    W5soz6 <= 1'b0;
  else
    W5soz6 <= D3n7v6;

always @(posedge FCLK) Z7soz6 <= Geg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pasoz6 <= 1'b0;
  else
    Pasoz6 <= W2n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Hdsoz6 <= 1'b0;
  else
    Hdsoz6 <= P2n7v6;

always @(posedge FCLK) Kfsoz6 <= Zdg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Aisoz6 <= 1'b0;
  else
    Aisoz6 <= I2n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Sksoz6 <= 1'b0;
  else
    Sksoz6 <= B2n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Vmsoz6 <= 1'b0;
  else
    Vmsoz6 <= U1n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Xosoz6 <= 1'b0;
  else
    Xosoz6 <= N1n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Pqsoz6 <= 1'b0;
  else
    Pqsoz6 <= G1n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Hssoz6 <= 1'b0;
  else
    Hssoz6 <= Z0n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ttsoz6 <= 1'b0;
  else
    Ttsoz6 <= Awg8v6;

always @(posedge SWCLKTCK) Ivsoz6 <= Hoh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Zwsoz6 <= 1'b0;
  else
    Zwsoz6 <= S0n7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Bzsoz6 <= 1'b0;
  else
    Bzsoz6 <= Vpg8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    E1toz6 <= 1'b0;
  else
    E1toz6 <= Uul8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Z2toz6 <= 1'b0;
  else
    Z2toz6 <= Qph8v6;

always @(posedge SWCLKTCK) C5toz6 <= Qih8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    U6toz6 <= 1'b0;
  else
    U6toz6 <= L0n7v6;

always @(posedge FCLK) X8toz6 <= Wfg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Nbtoz6 <= 1'b0;
  else
    Nbtoz6 <= E0n7v6;

always @(posedge SWCLKTCK) Fetoz6 <= Xih8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Xftoz6 <= 1'b0;
  else
    Xftoz6 <= Xzm7v6;

always @(posedge FCLK) Aitoz6 <= Dgg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qktoz6 <= 1'b0;
  else
    Qktoz6 <= Qzm7v6;

always @(posedge SWCLKTCK) Odazz6 <= Ejh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Gfazz6 <= 1'b0;
  else
    Gfazz6 <= Jzm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Jhazz6 <= 1'b0;
  else
    Jhazz6 <= Qqg8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ljazz6 <= 1'b0;
  else
    Ljazz6 <= Lqh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Flazz6 <= 1'b0;
  else
    Flazz6 <= Mpf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Gnazz6 <= 1'b0;
  else
    Gnazz6 <= U6h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Zoazz6 <= 1'b0;
  else
    Zoazz6 <= Czm7v6;

always @(posedge FCLK) Erazz6 <= Kgg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Utazz6 <= 1'b0;
  else
    Utazz6 <= Vym7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Mwazz6 <= 1'b0;
  else
    Mwazz6 <= N6h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Fyazz6 <= 1'b0;
  else
    Fyazz6 <= Oym7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    K0bzz6 <= 1'b0;
  else
    K0bzz6 <= Tpf8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    L2bzz6 <= 1'b0;
  else
    L2bzz6 <= Sqh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    F4bzz6 <= 1'b0;
  else
    F4bzz6 <= Xqg8v6;

always @(posedge SWCLKTCK) H6bzz6 <= Ljh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Z7bzz6 <= 1'b0;
  else
    Z7bzz6 <= Hym7v6;

always @(posedge FCLK) Cabzz6 <= Rgg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Scbzz6 <= 1'b0;
  else
    Scbzz6 <= Aym7v6;

always @(posedge SWCLKTCK) Kfbzz6 <= Sjh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Chbzz6 <= 1'b0;
  else
    Chbzz6 <= Txm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Fjbzz6 <= 1'b0;
  else
    Fjbzz6 <= Erg8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hlbzz6 <= 1'b0;
  else
    Hlbzz6 <= Zqh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Bnbzz6 <= 1'b0;
  else
    Bnbzz6 <= Aqf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Cpbzz6 <= 1'b0;
  else
    Cpbzz6 <= G6h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Vqbzz6 <= 1'b0;
  else
    Vqbzz6 <= Mxm7v6;

always @(posedge FCLK) Atbzz6 <= Ygg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qvbzz6 <= 1'b0;
  else
    Qvbzz6 <= Fxm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Iybzz6 <= 1'b0;
  else
    Iybzz6 <= Z5h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    B0czz6 <= 1'b0;
  else
    B0czz6 <= Ywm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    G2czz6 <= 1'b0;
  else
    G2czz6 <= Hqf8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    H4czz6 <= 1'b0;
  else
    H4czz6 <= Grh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    B6czz6 <= 1'b0;
  else
    B6czz6 <= Lrg8v6;

always @(posedge SWCLKTCK) D8czz6 <= Zjh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    V9czz6 <= 1'b0;
  else
    V9czz6 <= Rwm7v6;

always @(posedge FCLK) Ybczz6 <= Fhg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Oeczz6 <= 1'b0;
  else
    Oeczz6 <= Kwm7v6;

always @(posedge SWCLKTCK) Ghczz6 <= Gkh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Yiczz6 <= 1'b0;
  else
    Yiczz6 <= Dwm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Blczz6 <= 1'b0;
  else
    Blczz6 <= Srg8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dnczz6 <= 1'b0;
  else
    Dnczz6 <= Nrh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Xoczz6 <= 1'b0;
  else
    Xoczz6 <= Oqf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Yqczz6 <= 1'b0;
  else
    Yqczz6 <= S5h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Rsczz6 <= 1'b0;
  else
    Rsczz6 <= Wvm7v6;

always @(posedge FCLK) Wuczz6 <= Mhg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mxczz6 <= 1'b0;
  else
    Mxczz6 <= Pvm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    E0dzz6 <= 1'b0;
  else
    E0dzz6 <= L5h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    X1dzz6 <= 1'b0;
  else
    X1dzz6 <= Ivm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    C4dzz6 <= 1'b0;
  else
    C4dzz6 <= Vqf8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    D6dzz6 <= 1'b0;
  else
    D6dzz6 <= Urh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    X7dzz6 <= 1'b0;
  else
    X7dzz6 <= Zrg8v6;

always @(posedge SWCLKTCK) Z9dzz6 <= Nkh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Rbdzz6 <= 1'b0;
  else
    Rbdzz6 <= Bvm7v6;

always @(posedge FCLK) Uddzz6 <= Thg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kgdzz6 <= 1'b0;
  else
    Kgdzz6 <= Uum7v6;

always @(posedge SWCLKTCK) Cjdzz6 <= Ukh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ukdzz6 <= 1'b0;
  else
    Ukdzz6 <= Num7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Xmdzz6 <= 1'b0;
  else
    Xmdzz6 <= Gsg8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zodzz6 <= 1'b0;
  else
    Zodzz6 <= Bsh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Tqdzz6 <= 1'b0;
  else
    Tqdzz6 <= Crf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Usdzz6 <= 1'b0;
  else
    Usdzz6 <= E5h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Nudzz6 <= 1'b0;
  else
    Nudzz6 <= Gum7v6;

always @(posedge FCLK) Swdzz6 <= Aig8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Izdzz6 <= 1'b0;
  else
    Izdzz6 <= Ztm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    A2ezz6 <= 1'b0;
  else
    A2ezz6 <= X4h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    T3ezz6 <= 1'b0;
  else
    T3ezz6 <= Stm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Y5ezz6 <= 1'b0;
  else
    Y5ezz6 <= Jrf8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Z7ezz6 <= 1'b0;
  else
    Z7ezz6 <= Ish8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    T9ezz6 <= 1'b0;
  else
    T9ezz6 <= Nsg8v6;

always @(posedge SWCLKTCK) Vbezz6 <= Blh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ndezz6 <= 1'b0;
  else
    Ndezz6 <= Ltm7v6;

always @(posedge FCLK) Qfezz6 <= Hig8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Giezz6 <= 1'b0;
  else
    Giezz6 <= Etm7v6;

always @(posedge SWCLKTCK) Ykezz6 <= Ilh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Qmezz6 <= 1'b0;
  else
    Qmezz6 <= Xsm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Toezz6 <= 1'b0;
  else
    Toezz6 <= Usg8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vqezz6 <= 1'b0;
  else
    Vqezz6 <= Psh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Psezz6 <= 1'b0;
  else
    Psezz6 <= Qrf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Quezz6 <= 1'b0;
  else
    Quezz6 <= Q4h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Jwezz6 <= 1'b0;
  else
    Jwezz6 <= Qsm7v6;

always @(posedge FCLK) Oyezz6 <= Oig8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    E1fzz6 <= 1'b0;
  else
    E1fzz6 <= Jsm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    W3fzz6 <= 1'b0;
  else
    W3fzz6 <= J4h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    P5fzz6 <= 1'b0;
  else
    P5fzz6 <= Csm7v6;

always @(posedge FCLK) U7fzz6 <= Vig8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kafzz6 <= 1'b0;
  else
    Kafzz6 <= Vrm7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cdfzz6 <= 1'b0;
  else
    Cdfzz6 <= Kh88v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yefzz6 <= 1'b1;
  else
    Yefzz6 <= B9f8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vhfzz6 <= 1'b0;
  else
    Vhfzz6 <= Nmf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pkfzz6 <= 1'b0;
  else
    Pkfzz6 <= G5a7z6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cnfzz6 <= 1'b0;
  else
    Cnfzz6 <= Bt0ft6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ppfzz6 <= 1'b0;
  else
    Ppfzz6 <= Orm7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dsfzz6 <= 1'b0;
  else
    Dsfzz6 <= Xczet6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wufzz6 <= 1'b0;
  else
    Wufzz6 <= U71ft6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jxfzz6 <= 1'b0;
  else
    Jxfzz6 <= Hrm7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xzfzz6 <= 1'b0;
  else
    Xzfzz6 <= Pvl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P2gzz6 <= 1'b0;
  else
    P2gzz6 <= Arm7v6;

always @(posedge HCLK) P5gzz6 <= Y9g8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D8gzz6 <= 1'b0;
  else
    D8gzz6 <= Cm68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dbgzz6 <= 1'b0;
  else
    Dbgzz6 <= Jm68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Degzz6 <= 1'b0;
  else
    Degzz6 <= Qm68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dhgzz6 <= 1'b0;
  else
    Dhgzz6 <= Xm68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dkgzz6 <= 1'b0;
  else
    Dkgzz6 <= Bu88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cngzz6 <= 1'b0;
  else
    Cngzz6 <= S4yet6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wpgzz6 <= 1'b0;
  else
    Wpgzz6 <= M5l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Msgzz6 <= 1'b0;
  else
    Msgzz6 <= L3oet6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jvgzz6 <= 1'b0;
  else
    Jvgzz6 <= Hn48v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bygzz6 <= 1'b0;
  else
    Bygzz6 <= Y4l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D1hzz6 <= 1'b0;
  else
    D1hzz6 <= Mm48v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D4hzz6 <= 1'b0;
  else
    D4hzz6 <= Fm48v6;

always @(posedge HCLK) D7hzz6 <= Jh48v6;
always @(posedge HCLK) Gahzz6 <= Qh48v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jdhzz6 <= 1'b0;
  else
    Jdhzz6 <= Bqj8v6;

always @(posedge HCLK) Ighzz6 <= S5p7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mjhzz6 <= 1'b0;
  else
    Mjhzz6 <= Ijj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kmhzz6 <= 1'b0;
  else
    Kmhzz6 <= Rdj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tohzz6 <= 1'b0;
  else
    Tohzz6 <= Kdj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Prhzz6 <= 1'b0;
  else
    Prhzz6 <= Gt88v6;

always @(posedge HCLK) Duhzz6 <= Ols7v6;
always @(posedge HCLK) Rwhzz6 <= Uqx7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jzhzz6 <= 1'b0;
  else
    Jzhzz6 <= P8g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    D1izz6 <= 1'b0;
  else
    D1izz6 <= I8g8v6;

always @(posedge SWCLKTCK) U2izz6 <= Aoh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    L4izz6 <= 1'b0;
  else
    L4izz6 <= Tqm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    N6izz6 <= 1'b0;
  else
    N6izz6 <= Opg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Q8izz6 <= 1'b0;
  else
    Q8izz6 <= Lkg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Haizz6 <= 1'b0;
  else
    Haizz6 <= Skg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ybizz6 <= 1'b0;
  else
    Ybizz6 <= Cph8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ldizz6 <= 1'b0;
  else
    Ldizz6 <= Y1h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Dfizz6 <= 1'b0;
  else
    Dfizz6 <= Mqm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Hhizz6 <= 1'b0;
  else
    Hhizz6 <= R1h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ziizz6 <= 1'b0;
  else
    Ziizz6 <= Fqm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Dlizz6 <= 1'b0;
  else
    Dlizz6 <= K1h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Vmizz6 <= 1'b0;
  else
    Vmizz6 <= Ypm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Zoizz6 <= 1'b0;
  else
    Zoizz6 <= D1h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Rqizz6 <= 1'b0;
  else
    Rqizz6 <= Rpm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Vsizz6 <= 1'b0;
  else
    Vsizz6 <= W0h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Nuizz6 <= 1'b0;
  else
    Nuizz6 <= Kpm7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ewizz6 <= 1'b0;
  else
    Ewizz6 <= Fuh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Uyizz6 <= 1'b0;
  else
    Uyizz6 <= P0h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    M0jzz6 <= 1'b0;
  else
    M0jzz6 <= Dpm7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    D2jzz6 <= 1'b1;
  else
    D2jzz6 <= Ekg8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    X4jzz6 <= 1'b0;
  else
    X4jzz6 <= Wom7v6;

always @(posedge HCLK) N7jzz6 <= Ens7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fajzz6 <= 1'b0;
  else
    Fajzz6 <= Ldg8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zcjzz6 <= 1'b0;
  else
    Zcjzz6 <= Pom7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mfjzz6 <= 1'b0;
  else
    Mfjzz6 <= Cwh8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bijzz6 <= 1'b0;
  else
    Bijzz6 <= Ppzet6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rkjzz6 <= 1'b0;
  else
    Rkjzz6 <= Ov0ft6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bnjzz6 <= 1'b0;
  else
    Bnjzz6 <= Iom7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xpjzz6 <= 1'b0;
  else
    Xpjzz6 <= F5l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Osjzz6 <= 1'b0;
  else
    Osjzz6 <= Pnf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fvjzz6 <= 1'b0;
  else
    Fvjzz6 <= Inf8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rxjzz6 <= 1'b0;
  else
    Rxjzz6 <= Bom7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    H0kzz6 <= 1'b0;
  else
    H0kzz6 <= Unm7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Y2kzz6 <= 1'b0;
  else
    Y2kzz6 <= Muh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    O5kzz6 <= 1'b0;
  else
    O5kzz6 <= M9h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    G7kzz6 <= 1'b0;
  else
    G7kzz6 <= Nnm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    I9kzz6 <= 1'b0;
  else
    I9kzz6 <= Gnm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Kbkzz6 <= 1'b0;
  else
    Kbkzz6 <= Zmm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ndkzz6 <= 1'b0;
  else
    Ndkzz6 <= Smm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Qfkzz6 <= 1'b0;
  else
    Qfkzz6 <= Lmm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Thkzz6 <= 1'b0;
  else
    Thkzz6 <= Emm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Wjkzz6 <= 1'b0;
  else
    Wjkzz6 <= Xlm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Plkzz6 <= 1'b0;
  else
    Plkzz6 <= Qlm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Knkzz6 <= 1'b0;
  else
    Knkzz6 <= Jlm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Fpkzz6 <= 1'b0;
  else
    Fpkzz6 <= Clm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Xqkzz6 <= 1'b0;
  else
    Xqkzz6 <= Nul8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Zskzz6 <= 1'b0;
  else
    Zskzz6 <= Ovh8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Qukzz6 <= 1'b0;
  else
    Qukzz6 <= Vkm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Gwkzz6 <= 1'b0;
  else
    Gwkzz6 <= Okm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Wxkzz6 <= 1'b0;
  else
    Wxkzz6 <= Hkm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Mzkzz6 <= 1'b0;
  else
    Mzkzz6 <= Akm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    C1lzz6 <= 1'b0;
  else
    C1lzz6 <= Tjm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    S2lzz6 <= 1'b0;
  else
    S2lzz6 <= Mjm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    I4lzz6 <= 1'b0;
  else
    I4lzz6 <= Fjm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Y5lzz6 <= 1'b0;
  else
    Y5lzz6 <= Yim7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    S7lzz6 <= 1'b0;
  else
    S7lzz6 <= Rim7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    M9lzz6 <= 1'b0;
  else
    M9lzz6 <= Rth8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cclzz6 <= 1'b0;
  else
    Cclzz6 <= B1g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Xdlzz6 <= 1'b0;
  else
    Xdlzz6 <= U0g8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pflzz6 <= 1'b0;
  else
    Pflzz6 <= Dvf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Khlzz6 <= 1'b0;
  else
    Khlzz6 <= Wuf8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cjlzz6 <= 1'b0;
  else
    Cjlzz6 <= Twf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Xklzz6 <= 1'b0;
  else
    Xklzz6 <= Mwf8v6;

always @(posedge SWCLKTCK) Pmlzz6 <= Cih8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Holzz6 <= 1'b0;
  else
    Holzz6 <= Kim7v6;

always @(posedge FCLK) Kqlzz6 <= Ifg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Atlzz6 <= 1'b0;
  else
    Atlzz6 <= Dim7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Svlzz6 <= 1'b0;
  else
    Svlzz6 <= Ut88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gylzz6 <= 1'b0;
  else
    Gylzz6 <= Bnf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    S0mzz6 <= 1'b0;
  else
    S0mzz6 <= Dmyet6;

always @(posedge HCLK) L3mzz6 <= Whm7v6;
always @(posedge HCLK) B6mzz6 <= Phm7v6;
always @(posedge HCLK) R8mzz6 <= Ihm7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hbmzz6 <= 1'b0;
  else
    Hbmzz6 <= Dhyet6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wdmzz6 <= 1'b0;
  else
    Wdmzz6 <= Umf8v6;

always @(posedge HCLK) Igmzz6 <= K9o7v6;
always @(posedge HCLK) Mjmzz6 <= Gos7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qmmzz6 <= 1'b0;
  else
    Qmmzz6 <= H6l8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lpmzz6 <= 1'b0;
  else
    Lpmzz6 <= T5l8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ksmzz6 <= 1'b0;
  else
    Ksmzz6 <= A6l8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jvmzz6 <= 1'b0;
  else
    Jvmzz6 <= Hes7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Iymzz6 <= 1'b0;
  else
    Iymzz6 <= C7l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K1nzz6 <= 1'b0;
  else
    K1nzz6 <= Gak8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    B4nzz6 <= 1'b0;
  else
    B4nzz6 <= Bhm7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    V6nzz6 <= 1'b0;
  else
    V6nzz6 <= Wnf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    P9nzz6 <= 1'b0;
  else
    P9nzz6 <= Dof8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jcnzz6 <= 1'b0;
  else
    Jcnzz6 <= Stl8v6;

always @(posedge HCLK) Dfnzz6 <= Brx7v6;
always @(posedge HCLK) Vhnzz6 <= Lpx7v6;
always @(posedge HCLK) Nknzz6 <= Ves7v6;
always @(posedge HCLK) Cnnzz6 <= Dlx7v6;
always @(posedge HCLK) Upnzz6 <= Rqs7v6;
always @(posedge HCLK) Ysnzz6 <= Yqs7v6;
always @(posedge HCLK) Cwnzz6 <= Jfs7v6;
always @(posedge HCLK) Rynzz6 <= I4s7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    J1ozz6 <= 1'b0;
  else
    J1ozz6 <= Rvf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    E3ozz6 <= 1'b0;
  else
    E3ozz6 <= Kvf8v6;

always @(posedge SWCLKTCK) W4ozz6 <= Ohh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    O6ozz6 <= 1'b0;
  else
    O6ozz6 <= Ugm7v6;

always @(posedge FCLK) R8ozz6 <= Ueg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hbozz6 <= 1'b0;
  else
    Hbozz6 <= Ngm7v6;

always @(posedge SWCLKTCK) Zdozz6 <= Vhh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Rfozz6 <= 1'b0;
  else
    Rfozz6 <= Ggm7v6;

always @(posedge HCLK) Uhozz6 <= Imv7v6;
always @(posedge HCLK) Mkozz6 <= Cfs7v6;
always @(posedge HCLK) Bnozz6 <= Dqs7v6;
always @(posedge HCLK) Fqozz6 <= Kqs7v6;
always @(posedge FCLK) Jtozz6 <= Bfg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zvozz6 <= 1'b0;
  else
    Zvozz6 <= Zfm7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ryozz6 <= 1'b0;
  else
    Ryozz6 <= Fwf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    M0pzz6 <= 1'b0;
  else
    M0pzz6 <= Yvf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    E2pzz6 <= 1'b0;
  else
    E2pzz6 <= Mvg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    S3pzz6 <= 1'b0;
  else
    S3pzz6 <= Yng8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    L5pzz6 <= 1'b0;
  else
    L5pzz6 <= Fvg8v6;

always @(posedge HCLK) Z6pzz6 <= Pps7v6;
always @(posedge HCLK) Dapzz6 <= Wps7v6;
always @(posedge HCLK) Hdpzz6 <= Vls7v6;
always @(posedge HCLK) Vfpzz6 <= Nqx7v6;
always @(posedge HCLK) Nipzz6 <= Hg48v6;
always @(posedge HCLK) Qlpzz6 <= Og48v6;
always @(posedge HCLK) Topzz6 <= Cms7v6;
always @(posedge HCLK) Hrpzz6 <= Gqx7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ztpzz6 <= 1'b0;
  else
    Ztpzz6 <= N7g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Tvpzz6 <= 1'b0;
  else
    Tvpzz6 <= G7g8v6;

always @(posedge SWCLKTCK) Kxpzz6 <= Mnh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Bzpzz6 <= 1'b0;
  else
    Bzpzz6 <= Sfm7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    D1qzz6 <= 1'b0;
  else
    D1qzz6 <= Jjg8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    A4qzz6 <= 1'b0;
  else
    A4qzz6 <= Qjg8v6;

always @(posedge FCLK) X6qzz6 <= Tag8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    M9qzz6 <= 1'b0;
  else
    M9qzz6 <= Lfm7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dcqzz6 <= 1'b0;
  else
    Dcqzz6 <= J5g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Xdqzz6 <= 1'b0;
  else
    Xdqzz6 <= C5g8v6;

always @(posedge FCLK) Ofqzz6 <= Abg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Diqzz6 <= 1'b0;
  else
    Diqzz6 <= Efm7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ukqzz6 <= 1'b0;
  else
    Ukqzz6 <= X5g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Omqzz6 <= 1'b0;
  else
    Omqzz6 <= Q5g8v6;

always @(posedge SWCLKTCK) Foqzz6 <= Rmh8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Wpqzz6 <= 1'b0;
  else
    Wpqzz6 <= Xem7v6;

always @(posedge HCLK) Yrqzz6 <= Onx7v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Quqzz6 <= 1'b0;
  else
    Quqzz6 <= I0h8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Gwqzz6 <= 1'b0;
  else
    Gwqzz6 <= Apg8v6;

always @(posedge FCLK) Hyqzz6 <= Hbg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    W0rzz6 <= 1'b0;
  else
    W0rzz6 <= Qem7v6;

always @(posedge FCLK) N3rzz6 <= Obg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    C6rzz6 <= 1'b0;
  else
    C6rzz6 <= Jem7v6;

always @(posedge FCLK) T8rzz6 <= Vbg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ibrzz6 <= 1'b0;
  else
    Ibrzz6 <= Cem7v6;

always @(posedge FCLK) Zdrzz6 <= Ccg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ogrzz6 <= 1'b0;
  else
    Ogrzz6 <= Vdm7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fjrzz6 <= 1'b0;
  else
    Fjrzz6 <= Dh88v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Blrzz6 <= 1'b0;
  else
    Blrzz6 <= Pg88v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xmrzz6 <= 1'b0;
  else
    Xmrzz6 <= Wg88v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Torzz6 <= 1'b0;
  else
    Torzz6 <= Ig88v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pqrzz6 <= 1'b0;
  else
    Pqrzz6 <= Bg88v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lsrzz6 <= 1'b0;
  else
    Lsrzz6 <= Uf88v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hurzz6 <= 1'b0;
  else
    Hurzz6 <= B8g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Bwrzz6 <= 1'b0;
  else
    Bwrzz6 <= U7g8v6;

always @(posedge FCLK) Sxrzz6 <= Jcg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    H0szz6 <= 1'b0;
  else
    H0szz6 <= Odm7v6;

always @(posedge FCLK) Y2szz6 <= Qcg8v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    N5szz6 <= 1'b0;
  else
    N5szz6 <= D9g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    H7szz6 <= 1'b0;
  else
    H7szz6 <= W8g8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Y8szz6 <= 1'b0;
  else
    Y8szz6 <= Hdm7v6;

always @(posedge FCLK) Pbszz6 <= Xcg8v6;
always @(posedge FCLK) Eeszz6 <= Edg8v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tgszz6 <= 1'b0;
  else
    Tgszz6 <= Cjg8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ijszz6 <= 1'b0;
  else
    Ijszz6 <= Bizet6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vlszz6 <= 1'b0;
  else
    Vlszz6 <= K01ft6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Coszz6 <= 1'b0;
  else
    Coszz6 <= Mezet6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Vqszz6 <= 1'b0;
  else
    Vqszz6 <= Wtg8v6;

always @(posedge HCLK) Nsszz6 <= Vg48v6;
always @(posedge HCLK) Qvszz6 <= Ch48v6;
always @(posedge HCLK) Tyszz6 <= Jms7v6;
always @(posedge HCLK) H1tzz6 <= Zpx7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Z3tzz6 <= 1'b0;
  else
    Z3tzz6 <= Z6g8v6;

always @(posedge HCLK) T5tzz6 <= Qms7v6;
always @(posedge HCLK) H8tzz6 <= Spx7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zatzz6 <= 1'b0;
  else
    Zatzz6 <= L6g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Tctzz6 <= 1'b0;
  else
    Tctzz6 <= E6g8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ketzz6 <= 1'b1;
  else
    Ketzz6 <= Xjg8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dhtzz6 <= 1'b0;
  else
    Dhtzz6 <= Adm7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Sjtzz6 <= 1'b0;
  else
    Sjtzz6 <= Kp78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Oltzz6 <= 1'b0;
  else
    Oltzz6 <= Rp78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kntzz6 <= 1'b0;
  else
    Kntzz6 <= Fq78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gptzz6 <= 1'b0;
  else
    Gptzz6 <= Mq78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Crtzz6 <= 1'b0;
  else
    Crtzz6 <= Ar78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ystzz6 <= 1'b0;
  else
    Ystzz6 <= Js78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vutzz6 <= 1'b0;
  else
    Vutzz6 <= Qs78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Swtzz6 <= 1'b0;
  else
    Swtzz6 <= Xs78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pytzz6 <= 1'b0;
  else
    Pytzz6 <= Et78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    M0uzz6 <= 1'b0;
  else
    M0uzz6 <= Lt78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    J2uzz6 <= 1'b0;
  else
    J2uzz6 <= Yp78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F4uzz6 <= 1'b0;
  else
    F4uzz6 <= Tq78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    B6uzz6 <= 1'b0;
  else
    B6uzz6 <= Hr78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Y7uzz6 <= 1'b0;
  else
    Y7uzz6 <= Or78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    V9uzz6 <= 1'b0;
  else
    V9uzz6 <= St78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Sbuzz6 <= 1'b0;
  else
    Sbuzz6 <= Dqk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pduzz6 <= 1'b0;
  else
    Pduzz6 <= Sdo7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ofuzz6 <= 1'b0;
  else
    Ofuzz6 <= D16ft6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jhuzz6 <= 1'b1;
  else
    Jhuzz6 <= Z9k8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Hjuzz6 <= 1'b0;
  else
    Hjuzz6 <= Tvg8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vkuzz6 <= 1'b0;
  else
    Vkuzz6 <= Hxf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Qmuzz6 <= 1'b0;
  else
    Qmuzz6 <= Axf8v6;

always @(posedge SWCLKTCK) Iouzz6 <= Jih8v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Aquzz6 <= 1'b0;
  else
    Aquzz6 <= Tcm7v6;

always @(posedge HCLK) Dsuzz6 <= Wkx7v6;
always @(posedge FCLK) Vuuzz6 <= Pfg8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lxuzz6 <= 1'b0;
  else
    Lxuzz6 <= Mcm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    D0vzz6 <= 1'b0;
  else
    D0vzz6 <= Ulg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    R1vzz6 <= 1'b0;
  else
    R1vzz6 <= Fcm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    L3vzz6 <= 1'b0;
  else
    L3vzz6 <= Ybm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    F5vzz6 <= 1'b0;
  else
    F5vzz6 <= Rbm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    V6vzz6 <= 1'b0;
  else
    V6vzz6 <= Kbm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    S8vzz6 <= 1'b1;
  else
    S8vzz6 <= Dbm7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Iavzz6 <= 1'b1;
  else
    Iavzz6 <= Wam7v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ybvzz6 <= 1'b0;
  else
    Ybvzz6 <= Lsf8v6;

always @(posedge HCLK) Odvzz6 <= Tf48v6;
always @(posedge HCLK) Rgvzz6 <= Ag48v6;
always @(posedge HCLK) Ujvzz6 <= Epx7v6;
always @(posedge HCLK) Mmvzz6 <= Djs7v6;
always @(posedge HCLK) Bpvzz6 <= Nj48v6;
always @(posedge HCLK) Fsvzz6 <= Uj48v6;
always @(posedge HCLK) Jvvzz6 <= Xox7v6;
always @(posedge HCLK) Byvzz6 <= Kjs7v6;
always @(posedge HCLK) Q0wzz6 <= Bk48v6;
always @(posedge HCLK) U3wzz6 <= Ik48v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y6wzz6 <= 1'b0;
  else
    Y6wzz6 <= Krj8v6;

always @(posedge HCLK) X9wzz6 <= J4p7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bdwzz6 <= 1'b0;
  else
    Bdwzz6 <= Cnj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Agwzz6 <= 1'b0;
  else
    Agwzz6 <= Vmj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Eiwzz6 <= 1'b0;
  else
    Eiwzz6 <= Omj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ikwzz6 <= 1'b0;
  else
    Ikwzz6 <= Ebi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jnwzz6 <= 1'b0;
  else
    Jnwzz6 <= Zbi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mqwzz6 <= 1'b0;
  else
    Mqwzz6 <= U3d7z6[3];

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Otwzz6 <= 1'b0;
  else
    Otwzz6 <= Nci8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rwwzz6 <= 1'b0;
  else
    Rwwzz6 <= U3d7z6[5];

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tzwzz6 <= 1'b0;
  else
    Tzwzz6 <= Uci8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W2xzz6 <= 1'b0;
  else
    W2xzz6 <= U3d7z6[0];

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y5xzz6 <= 1'b0;
  else
    Y5xzz6 <= Sbi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B9xzz6 <= 1'b0;
  else
    B9xzz6 <= Gci8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ecxzz6 <= 1'b0;
  else
    Ecxzz6 <= U3d7z6[4];

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gfxzz6 <= 1'b0;
  else
    Gfxzz6 <= U3d7z6[2];

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Iixzz6 <= 1'b0;
  else
    Iixzz6 <= Drj8v6;

always @(posedge HCLK) Hlxzz6 <= Q4p7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Loxzz6 <= 1'b0;
  else
    Loxzz6 <= Amj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Krxzz6 <= 1'b0;
  else
    Krxzz6 <= Qai8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ktxzz6 <= 1'b0;
  else
    Ktxzz6 <= Pam7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lwxzz6 <= 1'b0;
  else
    Lwxzz6 <= Jai8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lyxzz6 <= 1'b0;
  else
    Lyxzz6 <= Xsddt6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M0yzz6 <= 1'b0;
  else
    M0yzz6 <= V9i8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N2yzz6 <= 1'b0;
  else
    N2yzz6 <= O9i8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O4yzz6 <= 1'b0;
  else
    O4yzz6 <= Cp38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q6yzz6 <= 1'b0;
  else
    Q6yzz6 <= Flj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q8yzz6 <= 1'b0;
  else
    Q8yzz6 <= Hmj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vayzz6 <= 1'b0;
  else
    Vayzz6 <= A0k8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ycyzz6 <= 1'b0;
  else
    Ycyzz6 <= D4adt6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Weyzz6 <= 1'b0;
  else
    Weyzz6 <= Iam7v6;

always @(posedge HCLK) Ygyzz6 <= Y8p7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ckyzz6 <= 1'b0;
  else
    Ckyzz6 <= G2l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fnyzz6 <= 1'b0;
  else
    Fnyzz6 <= Uij8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ipyzz6 <= 1'b0;
  else
    Ipyzz6 <= Pjj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nryzz6 <= 1'b0;
  else
    Nryzz6 <= Cai8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ptyzz6 <= 1'b0;
  else
    Ptyzz6 <= Ubj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xvyzz6 <= 1'b0;
  else
    Xvyzz6 <= Dv88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uyyzz6 <= 1'b0;
  else
    Uyyzz6 <= Kv88v6;

always @(posedge HCLK) R1zzz6 <= R8p7v6;
always @(posedge HCLK) V4zzz6 <= Qox7v6;
always @(posedge HCLK) N7zzz6 <= Rjs7v6;
always @(posedge HCLK) Cazzz6 <= Pk48v6;
always @(posedge HCLK) Gdzzz6 <= Wk48v6;
always @(posedge HCLK) Kgzzz6 <= Jox7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cjzzz6 <= 1'b0;
  else
    Cjzzz6 <= F3g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Xkzzz6 <= 1'b0;
  else
    Xkzzz6 <= Y2g8v6;

always @(posedge HCLK) Pmzzz6 <= Yjs7v6;
always @(posedge HCLK) Epzzz6 <= Dl48v6;
always @(posedge HCLK) Iszzz6 <= Kl48v6;
always @(posedge HCLK) Mvzzz6 <= Cox7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Eyzzz6 <= 1'b0;
  else
    Eyzzz6 <= R2g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Zzzzz6 <= 1'b0;
  else
    Zzzzz6 <= K2g8v6;

always @(posedge HCLK) R10007 <= Fks7v6;
always @(posedge HCLK) G40007 <= W7p7v6;
always @(posedge HCLK) K70007 <= R9o7v6;
always @(posedge HCLK) Oa0007 <= Rl48v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sd0007 <= 1'b0;
  else
    Sd0007 <= Fsj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rg0007 <= 1'b0;
  else
    Rg0007 <= Bjj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cj0007 <= 1'b0;
  else
    Cj0007 <= Dkj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nl0007 <= 1'b0;
  else
    Nl0007 <= Kkj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yn0007 <= 1'b0;
  else
    Yn0007 <= Rkj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jq0007 <= 1'b0;
  else
    Jq0007 <= Wjj8v6;

always @(posedge HCLK) Os0007 <= K408v6;
always @(posedge HCLK) Ev0007 <= F508v6;
always @(posedge HCLK) Ux0007 <= M508v6;
always @(posedge HCLK) K01007 <= A608v6;
always @(posedge HCLK) A31007 <= I038v6;
always @(posedge HCLK) R51007 <= V608v6;
always @(posedge HCLK) I81007 <= D138v6;
always @(posedge HCLK) Ab1007 <= C708v6;
always @(posedge HCLK) Rd1007 <= K138v6;
always @(posedge HCLK) Jg1007 <= J708v6;
always @(posedge HCLK) Aj1007 <= R138v6;
always @(posedge HCLK) Sl1007 <= X708v6;
always @(posedge HCLK) Jo1007 <= F238v6;
always @(posedge HCLK) Br1007 <= E808v6;
always @(posedge HCLK) St1007 <= M238v6;
always @(posedge HCLK) Kw1007 <= S808v6;
always @(posedge HCLK) Bz1007 <= A338v6;
always @(posedge HCLK) T12007 <= Z808v6;
always @(posedge HCLK) K42007 <= H338v6;
always @(posedge HCLK) C72007 <= G908v6;
always @(posedge HCLK) T92007 <= O338v6;
always @(posedge HCLK) Lc2007 <= N908v6;
always @(posedge HCLK) Cf2007 <= V338v6;
always @(posedge HCLK) Uh2007 <= U908v6;
always @(posedge HCLK) Lk2007 <= C438v6;
always @(posedge HCLK) Dn2007 <= Ba08v6;
always @(posedge HCLK) Up2007 <= J438v6;
always @(posedge HCLK) Ms2007 <= Ia08v6;
always @(posedge HCLK) Dv2007 <= Q438v6;
always @(posedge HCLK) Vx2007 <= H608v6;
always @(posedge HCLK) M03007 <= P038v6;
always @(posedge HCLK) E33007 <= L808v6;
always @(posedge HCLK) V53007 <= T238v6;
always @(posedge HCLK) N83007 <= Pa08v6;
always @(posedge HCLK) Eb3007 <= X438v6;
always @(posedge HCLK) Wd3007 <= R408v6;
always @(posedge HCLK) Mg3007 <= D408v6;
always @(posedge HCLK) Cj3007 <= N638v6;
always @(posedge HCLK) Tl3007 <= T508v6;
always @(posedge HCLK) Jo3007 <= Wa08v6;
always @(posedge HCLK) Ar3007 <= E538v6;
always @(posedge HCLK) St3007 <= Q708v6;
always @(posedge HCLK) Jw3007 <= Y138v6;
always @(posedge HCLK) Bz3007 <= Kb08v6;
always @(posedge HCLK) S14007 <= S538v6;
always @(posedge HCLK) K44007 <= Db08v6;
always @(posedge HCLK) B74007 <= L538v6;
always @(posedge HCLK) T94007 <= Zuz7v6;
always @(posedge HCLK) Jc4007 <= Luz7v6;
always @(posedge HCLK) Af4007 <= Euz7v6;
always @(posedge HCLK) Rh4007 <= Xtz7v6;
always @(posedge HCLK) Ik4007 <= Qtz7v6;
always @(posedge HCLK) Zm4007 <= Jtz7v6;
always @(posedge HCLK) Qp4007 <= Ctz7v6;
always @(posedge HCLK) Hs4007 <= Vsz7v6;
always @(posedge HCLK) Yu4007 <= Osz7v6;
always @(posedge HCLK) Px4007 <= Hsz7v6;
always @(posedge HCLK) G05007 <= Asz7v6;
always @(posedge HCLK) X25007 <= Trz7v6;
always @(posedge HCLK) O55007 <= Mrz7v6;
always @(posedge HCLK) F85007 <= Frz7v6;
always @(posedge HCLK) Wa5007 <= Yqz7v6;
always @(posedge HCLK) Nd5007 <= Rqz7v6;
always @(posedge HCLK) Eg5007 <= Kqz7v6;
always @(posedge HCLK) Vi5007 <= Dqz7v6;
always @(posedge HCLK) Ml5007 <= Wpz7v6;
always @(posedge HCLK) Do5007 <= Ppz7v6;
always @(posedge HCLK) Uq5007 <= Ipz7v6;
always @(posedge HCLK) Lt5007 <= Bpz7v6;
always @(posedge HCLK) Cw5007 <= Uoz7v6;
always @(posedge HCLK) Sy5007 <= Noz7v6;
always @(posedge HCLK) I16007 <= Goz7v6;
always @(posedge HCLK) Y36007 <= Znz7v6;
always @(posedge HCLK) O66007 <= Snz7v6;
always @(posedge HCLK) E96007 <= Lnz7v6;
always @(posedge HCLK) Ub6007 <= Enz7v6;
always @(posedge HCLK) Ke6007 <= Xmz7v6;
always @(posedge HCLK) Ah6007 <= Qmz7v6;
always @(posedge HCLK) Qj6007 <= Lt08v6;
always @(posedge HCLK) Gm6007 <= Xs08v6;
always @(posedge HCLK) Xo6007 <= Qs08v6;
always @(posedge HCLK) Or6007 <= Js08v6;
always @(posedge HCLK) Fu6007 <= Cs08v6;
always @(posedge HCLK) Ww6007 <= Vr08v6;
always @(posedge HCLK) Nz6007 <= Or08v6;
always @(posedge HCLK) E27007 <= Hr08v6;
always @(posedge HCLK) V47007 <= Ar08v6;
always @(posedge HCLK) M77007 <= Tq08v6;
always @(posedge HCLK) Da7007 <= Mq08v6;
always @(posedge HCLK) Uc7007 <= Fq08v6;
always @(posedge HCLK) Lf7007 <= Yp08v6;
always @(posedge HCLK) Ci7007 <= Rp08v6;
always @(posedge HCLK) Tk7007 <= Kp08v6;
always @(posedge HCLK) Kn7007 <= Dp08v6;
always @(posedge HCLK) Bq7007 <= Wo08v6;
always @(posedge HCLK) Ss7007 <= Po08v6;
always @(posedge HCLK) Jv7007 <= Io08v6;
always @(posedge HCLK) Ay7007 <= Bo08v6;
always @(posedge HCLK) R08007 <= Un08v6;
always @(posedge HCLK) I38007 <= Nn08v6;
always @(posedge HCLK) Z58007 <= Gn08v6;
always @(posedge HCLK) P88007 <= Zm08v6;
always @(posedge HCLK) Fb8007 <= Sm08v6;
always @(posedge HCLK) Vd8007 <= Lm08v6;
always @(posedge HCLK) Lg8007 <= Em08v6;
always @(posedge HCLK) Bj8007 <= Xl08v6;
always @(posedge HCLK) Rl8007 <= Ql08v6;
always @(posedge HCLK) Ho8007 <= Jl08v6;
always @(posedge HCLK) Xq8007 <= Cl08v6;
always @(posedge HCLK) Nt8007 <= Ra18v6;
always @(posedge HCLK) Dw8007 <= Da18v6;
always @(posedge HCLK) Uy8007 <= W918v6;
always @(posedge HCLK) L19007 <= P918v6;
always @(posedge HCLK) C49007 <= I918v6;
always @(posedge HCLK) T69007 <= B918v6;
always @(posedge HCLK) K99007 <= U818v6;
always @(posedge HCLK) Bc9007 <= N818v6;
always @(posedge HCLK) Se9007 <= G818v6;
always @(posedge HCLK) Jh9007 <= Z718v6;
always @(posedge HCLK) Ak9007 <= S718v6;
always @(posedge HCLK) Rm9007 <= L718v6;
always @(posedge HCLK) Ip9007 <= E718v6;
always @(posedge HCLK) Zr9007 <= X618v6;
always @(posedge HCLK) Qu9007 <= Q618v6;
always @(posedge HCLK) Hx9007 <= J618v6;
always @(posedge HCLK) Yz9007 <= C618v6;
always @(posedge HCLK) P2a007 <= V518v6;
always @(posedge HCLK) G5a007 <= O518v6;
always @(posedge HCLK) X7a007 <= H518v6;
always @(posedge HCLK) Oaa007 <= A518v6;
always @(posedge HCLK) Fda007 <= T418v6;
always @(posedge HCLK) Wfa007 <= M418v6;
always @(posedge HCLK) Mia007 <= F418v6;
always @(posedge HCLK) Cla007 <= Y318v6;
always @(posedge HCLK) Sna007 <= R318v6;
always @(posedge HCLK) Iqa007 <= K318v6;
always @(posedge HCLK) Ysa007 <= D318v6;
always @(posedge HCLK) Ova007 <= W218v6;
always @(posedge HCLK) Eya007 <= P218v6;
always @(posedge HCLK) U0b007 <= I218v6;
always @(posedge HCLK) K3b007 <= Hj18v6;
always @(posedge HCLK) A6b007 <= Ti18v6;
always @(posedge HCLK) R8b007 <= Mi18v6;
always @(posedge HCLK) Ibb007 <= Fi18v6;
always @(posedge HCLK) Zdb007 <= Yh18v6;
always @(posedge HCLK) Qgb007 <= Rh18v6;
always @(posedge HCLK) Hjb007 <= Kh18v6;
always @(posedge HCLK) Ylb007 <= Dh18v6;
always @(posedge HCLK) Pob007 <= Wg18v6;
always @(posedge HCLK) Grb007 <= Pg18v6;
always @(posedge HCLK) Xtb007 <= Ig18v6;
always @(posedge HCLK) Owb007 <= Bg18v6;
always @(posedge HCLK) Fzb007 <= Uf18v6;
always @(posedge HCLK) W1c007 <= Nf18v6;
always @(posedge HCLK) N4c007 <= Gf18v6;
always @(posedge HCLK) E7c007 <= Ze18v6;
always @(posedge HCLK) V9c007 <= Se18v6;
always @(posedge HCLK) Mcc007 <= Le18v6;
always @(posedge HCLK) Dfc007 <= Ee18v6;
always @(posedge HCLK) Uhc007 <= Xd18v6;
always @(posedge HCLK) Lkc007 <= Qd18v6;
always @(posedge HCLK) Cnc007 <= Jd18v6;
always @(posedge HCLK) Tpc007 <= Cd18v6;
always @(posedge HCLK) Jsc007 <= Vc18v6;
always @(posedge HCLK) Zuc007 <= Oc18v6;
always @(posedge HCLK) Pxc007 <= Hc18v6;
always @(posedge HCLK) F0d007 <= Ac18v6;
always @(posedge HCLK) V2d007 <= Tb18v6;
always @(posedge HCLK) L5d007 <= Mb18v6;
always @(posedge HCLK) B8d007 <= Fb18v6;
always @(posedge HCLK) Rad007 <= Ya18v6;
always @(posedge HCLK) Hdd007 <= Xr18v6;
always @(posedge HCLK) Xfd007 <= Jr18v6;
always @(posedge HCLK) Oid007 <= Cr18v6;
always @(posedge HCLK) Fld007 <= Vq18v6;
always @(posedge HCLK) Wnd007 <= Oq18v6;
always @(posedge HCLK) Nqd007 <= Hq18v6;
always @(posedge HCLK) Etd007 <= Aq18v6;
always @(posedge HCLK) Vvd007 <= Tp18v6;
always @(posedge HCLK) Myd007 <= Mp18v6;
always @(posedge HCLK) D1e007 <= Fp18v6;
always @(posedge HCLK) U3e007 <= Yo18v6;
always @(posedge HCLK) L6e007 <= Ro18v6;
always @(posedge HCLK) C9e007 <= Ko18v6;
always @(posedge HCLK) Tbe007 <= Do18v6;
always @(posedge HCLK) Kee007 <= Wn18v6;
always @(posedge HCLK) Bhe007 <= Pn18v6;
always @(posedge HCLK) Sje007 <= In18v6;
always @(posedge HCLK) Jme007 <= Bn18v6;
always @(posedge HCLK) Ape007 <= Um18v6;
always @(posedge HCLK) Rre007 <= Nm18v6;
always @(posedge HCLK) Iue007 <= Gm18v6;
always @(posedge HCLK) Zwe007 <= Zl18v6;
always @(posedge HCLK) Qze007 <= Sl18v6;
always @(posedge HCLK) G2f007 <= Ll18v6;
always @(posedge HCLK) W4f007 <= El18v6;
always @(posedge HCLK) M7f007 <= Xk18v6;
always @(posedge HCLK) Caf007 <= Qk18v6;
always @(posedge HCLK) Scf007 <= Jk18v6;
always @(posedge HCLK) Iff007 <= Ck18v6;
always @(posedge HCLK) Yhf007 <= Vj18v6;
always @(posedge HCLK) Okf007 <= Oj18v6;
always @(posedge HCLK) Enf007 <= N028v6;
always @(posedge HCLK) Vpf007 <= Zz18v6;
always @(posedge HCLK) Nsf007 <= Sz18v6;
always @(posedge HCLK) Fvf007 <= Lz18v6;
always @(posedge HCLK) Xxf007 <= Ez18v6;
always @(posedge HCLK) P0g007 <= Xy18v6;
always @(posedge HCLK) H3g007 <= Qy18v6;
always @(posedge HCLK) Z5g007 <= Jy18v6;
always @(posedge HCLK) R8g007 <= Cy18v6;
always @(posedge HCLK) Jbg007 <= Vx18v6;
always @(posedge HCLK) Beg007 <= Ox18v6;
always @(posedge HCLK) Tgg007 <= Hx18v6;
always @(posedge HCLK) Ljg007 <= Ax18v6;
always @(posedge HCLK) Dmg007 <= Tw18v6;
always @(posedge HCLK) Vog007 <= Mw18v6;
always @(posedge HCLK) Nrg007 <= Fw18v6;
always @(posedge HCLK) Fug007 <= Yv18v6;
always @(posedge HCLK) Xwg007 <= Rv18v6;
always @(posedge HCLK) Pzg007 <= Kv18v6;
always @(posedge HCLK) H2h007 <= Dv18v6;
always @(posedge HCLK) Z4h007 <= Wu18v6;
always @(posedge HCLK) R7h007 <= Pu18v6;
always @(posedge HCLK) Jah007 <= Iu18v6;
always @(posedge HCLK) Adh007 <= Bu18v6;
always @(posedge HCLK) Rfh007 <= Ut18v6;
always @(posedge HCLK) Iih007 <= Nt18v6;
always @(posedge HCLK) Zkh007 <= Gt18v6;
always @(posedge HCLK) Qnh007 <= Zs18v6;
always @(posedge HCLK) Hqh007 <= Ss18v6;
always @(posedge HCLK) Ysh007 <= Ls18v6;
always @(posedge HCLK) Pvh007 <= Es18v6;
always @(posedge HCLK) Gyh007 <= D928v6;
always @(posedge HCLK) X0i007 <= P828v6;
always @(posedge HCLK) P3i007 <= I828v6;
always @(posedge HCLK) H6i007 <= B828v6;
always @(posedge HCLK) Z8i007 <= U728v6;
always @(posedge HCLK) Rbi007 <= N728v6;
always @(posedge HCLK) Jei007 <= G728v6;
always @(posedge HCLK) Bhi007 <= Z628v6;
always @(posedge HCLK) Tji007 <= S628v6;
always @(posedge HCLK) Lmi007 <= L628v6;
always @(posedge HCLK) Dpi007 <= E628v6;
always @(posedge HCLK) Vri007 <= X528v6;
always @(posedge HCLK) Nui007 <= Q528v6;
always @(posedge HCLK) Fxi007 <= J528v6;
always @(posedge HCLK) Xzi007 <= C528v6;
always @(posedge HCLK) P2j007 <= V428v6;
always @(posedge HCLK) H5j007 <= O428v6;
always @(posedge HCLK) Z7j007 <= H428v6;
always @(posedge HCLK) Raj007 <= A428v6;
always @(posedge HCLK) Jdj007 <= T328v6;
always @(posedge HCLK) Bgj007 <= M328v6;
always @(posedge HCLK) Tij007 <= F328v6;
always @(posedge HCLK) Llj007 <= Y228v6;
always @(posedge HCLK) Coj007 <= R228v6;
always @(posedge HCLK) Tqj007 <= K228v6;
always @(posedge HCLK) Ktj007 <= D228v6;
always @(posedge HCLK) Bwj007 <= W128v6;
always @(posedge HCLK) Syj007 <= P128v6;
always @(posedge HCLK) J1k007 <= I128v6;
always @(posedge HCLK) A4k007 <= B128v6;
always @(posedge HCLK) R6k007 <= U028v6;
always @(posedge HCLK) I9k007 <= Th28v6;
always @(posedge HCLK) Zbk007 <= Fh28v6;
always @(posedge HCLK) Rek007 <= Yg28v6;
always @(posedge HCLK) Jhk007 <= Rg28v6;
always @(posedge HCLK) Bkk007 <= Kg28v6;
always @(posedge HCLK) Tmk007 <= Dg28v6;
always @(posedge HCLK) Lpk007 <= Wf28v6;
always @(posedge HCLK) Dsk007 <= Pf28v6;
always @(posedge HCLK) Vuk007 <= If28v6;
always @(posedge HCLK) Nxk007 <= Bf28v6;
always @(posedge HCLK) F0l007 <= Ue28v6;
always @(posedge HCLK) X2l007 <= Ne28v6;
always @(posedge HCLK) P5l007 <= Ge28v6;
always @(posedge HCLK) H8l007 <= Zd28v6;
always @(posedge HCLK) Zal007 <= Sd28v6;
always @(posedge HCLK) Rdl007 <= Ld28v6;
always @(posedge HCLK) Jgl007 <= Ed28v6;
always @(posedge HCLK) Bjl007 <= Xc28v6;
always @(posedge HCLK) Tll007 <= Qc28v6;
always @(posedge HCLK) Lol007 <= Jc28v6;
always @(posedge HCLK) Drl007 <= Cc28v6;
always @(posedge HCLK) Vtl007 <= Vb28v6;
always @(posedge HCLK) Nwl007 <= Ob28v6;
always @(posedge HCLK) Ezl007 <= Hb28v6;
always @(posedge HCLK) V1m007 <= Ab28v6;
always @(posedge HCLK) M4m007 <= Ta28v6;
always @(posedge HCLK) D7m007 <= Ma28v6;
always @(posedge HCLK) U9m007 <= Fa28v6;
always @(posedge HCLK) Lcm007 <= Y928v6;
always @(posedge HCLK) Cfm007 <= R928v6;
always @(posedge HCLK) Thm007 <= K928v6;
always @(posedge HCLK) Kkm007 <= Vp28v6;
always @(posedge HCLK) Bnm007 <= Hp28v6;
always @(posedge HCLK) Tpm007 <= Ap28v6;
always @(posedge HCLK) Lsm007 <= To28v6;
always @(posedge HCLK) Dvm007 <= Mo28v6;
always @(posedge HCLK) Vxm007 <= Fo28v6;
always @(posedge HCLK) N0n007 <= Yn28v6;
always @(posedge HCLK) F3n007 <= Rn28v6;
always @(posedge HCLK) X5n007 <= Kn28v6;
always @(posedge HCLK) P8n007 <= Dn28v6;
always @(posedge HCLK) Hbn007 <= Wm28v6;
always @(posedge HCLK) Zdn007 <= Pm28v6;
always @(posedge HCLK) Rgn007 <= Im28v6;
always @(posedge HCLK) Jjn007 <= Bm28v6;
always @(posedge HCLK) Bmn007 <= Ul28v6;
always @(posedge HCLK) Ton007 <= Nl28v6;
always @(posedge HCLK) Lrn007 <= Gl28v6;
always @(posedge HCLK) Dun007 <= Zk28v6;
always @(posedge HCLK) Vwn007 <= Sk28v6;
always @(posedge HCLK) Nzn007 <= Lk28v6;
always @(posedge HCLK) F2o007 <= Ek28v6;
always @(posedge HCLK) X4o007 <= Xj28v6;
always @(posedge HCLK) P7o007 <= Qj28v6;
always @(posedge HCLK) Gao007 <= Jj28v6;
always @(posedge HCLK) Xco007 <= Cj28v6;
always @(posedge HCLK) Ofo007 <= Vi28v6;
always @(posedge HCLK) Fio007 <= Oi28v6;
always @(posedge HCLK) Wko007 <= Hi28v6;
always @(posedge HCLK) Nno007 <= Ai28v6;
always @(posedge HCLK) Eqo007 <= Ly28v6;
always @(posedge HCLK) Vso007 <= Xx28v6;
always @(posedge HCLK) Nvo007 <= Qx28v6;
always @(posedge HCLK) Fyo007 <= Jx28v6;
always @(posedge HCLK) X0p007 <= Cx28v6;
always @(posedge HCLK) P3p007 <= Vw28v6;
always @(posedge HCLK) H6p007 <= Ow28v6;
always @(posedge HCLK) Z8p007 <= Hw28v6;
always @(posedge HCLK) Rbp007 <= Aw28v6;
always @(posedge HCLK) Jep007 <= Tv28v6;
always @(posedge HCLK) Bhp007 <= Mv28v6;
always @(posedge HCLK) Tjp007 <= Fv28v6;
always @(posedge HCLK) Lmp007 <= Yu28v6;
always @(posedge HCLK) Dpp007 <= Ru28v6;
always @(posedge HCLK) Vrp007 <= Ku28v6;
always @(posedge HCLK) Nup007 <= Du28v6;
always @(posedge HCLK) Fxp007 <= Wt28v6;
always @(posedge HCLK) Xzp007 <= Pt28v6;
always @(posedge HCLK) P2q007 <= It28v6;
always @(posedge HCLK) H5q007 <= Bt28v6;
always @(posedge HCLK) Z7q007 <= Us28v6;
always @(posedge HCLK) Raq007 <= Ns28v6;
always @(posedge HCLK) Jdq007 <= Gs28v6;
always @(posedge HCLK) Agq007 <= Zr28v6;
always @(posedge HCLK) Riq007 <= Sr28v6;
always @(posedge HCLK) Ilq007 <= Lr28v6;
always @(posedge HCLK) Znq007 <= Er28v6;
always @(posedge HCLK) Qqq007 <= Xq28v6;
always @(posedge HCLK) Htq007 <= Qq28v6;
always @(posedge HCLK) Yvq007 <= Jq28v6;
always @(posedge HCLK) Pyq007 <= Cq28v6;
always @(posedge HCLK) G1r007 <= P308v6;
always @(posedge HCLK) W3r007 <= B308v6;
always @(posedge HCLK) N6r007 <= U208v6;
always @(posedge HCLK) E9r007 <= N208v6;
always @(posedge HCLK) Vbr007 <= G208v6;
always @(posedge HCLK) Mer007 <= Z108v6;
always @(posedge HCLK) Dhr007 <= S108v6;
always @(posedge HCLK) Ujr007 <= L108v6;
always @(posedge HCLK) Lmr007 <= E108v6;
always @(posedge HCLK) Cpr007 <= X008v6;
always @(posedge HCLK) Trr007 <= Q008v6;
always @(posedge HCLK) Kur007 <= J008v6;
always @(posedge HCLK) Bxr007 <= C008v6;
always @(posedge HCLK) Szr007 <= Vzz7v6;
always @(posedge HCLK) J2s007 <= Ozz7v6;
always @(posedge HCLK) A5s007 <= Hzz7v6;
always @(posedge HCLK) R7s007 <= Azz7v6;
always @(posedge HCLK) Ias007 <= Tyz7v6;
always @(posedge HCLK) Zcs007 <= Myz7v6;
always @(posedge HCLK) Qfs007 <= Fyz7v6;
always @(posedge HCLK) His007 <= Yxz7v6;
always @(posedge HCLK) Yks007 <= Rxz7v6;
always @(posedge HCLK) Pns007 <= Kxz7v6;
always @(posedge HCLK) Fqs007 <= Dxz7v6;
always @(posedge HCLK) Vss007 <= Wwz7v6;
always @(posedge HCLK) Lvs007 <= Pwz7v6;
always @(posedge HCLK) Bys007 <= Iwz7v6;
always @(posedge HCLK) R0t007 <= Bwz7v6;
always @(posedge HCLK) H3t007 <= Uvz7v6;
always @(posedge HCLK) X5t007 <= Nvz7v6;
always @(posedge HCLK) N8t007 <= Gvz7v6;
always @(posedge HCLK) Dbt007 <= Vk08v6;
always @(posedge HCLK) Tdt007 <= Hk08v6;
always @(posedge HCLK) Kgt007 <= Ak08v6;
always @(posedge HCLK) Bjt007 <= Tj08v6;
always @(posedge HCLK) Slt007 <= Mj08v6;
always @(posedge HCLK) Jot007 <= Fj08v6;
always @(posedge HCLK) Art007 <= Yi08v6;
always @(posedge HCLK) Rtt007 <= Ri08v6;
always @(posedge HCLK) Iwt007 <= Ki08v6;
always @(posedge HCLK) Zyt007 <= Di08v6;
always @(posedge HCLK) Q1u007 <= Wh08v6;
always @(posedge HCLK) H4u007 <= Ph08v6;
always @(posedge HCLK) Y6u007 <= Ih08v6;
always @(posedge HCLK) P9u007 <= Bh08v6;
always @(posedge HCLK) Gcu007 <= Ug08v6;
always @(posedge HCLK) Xeu007 <= Ng08v6;
always @(posedge HCLK) Ohu007 <= Gg08v6;
always @(posedge HCLK) Fku007 <= Zf08v6;
always @(posedge HCLK) Wmu007 <= Sf08v6;
always @(posedge HCLK) Npu007 <= Lf08v6;
always @(posedge HCLK) Esu007 <= Ef08v6;
always @(posedge HCLK) Vuu007 <= Xe08v6;
always @(posedge HCLK) Mxu007 <= Qe08v6;
always @(posedge HCLK) C0v007 <= Je08v6;
always @(posedge HCLK) S2v007 <= Ce08v6;
always @(posedge HCLK) I5v007 <= Vd08v6;
always @(posedge HCLK) Y7v007 <= Od08v6;
always @(posedge HCLK) Oav007 <= Hd08v6;
always @(posedge HCLK) Edv007 <= Ad08v6;
always @(posedge HCLK) Ufv007 <= Tc08v6;
always @(posedge HCLK) Kiv007 <= Mc08v6;
always @(posedge HCLK) Alv007 <= B218v6;
always @(posedge HCLK) Qnv007 <= N118v6;
always @(posedge HCLK) Hqv007 <= G118v6;
always @(posedge HCLK) Ysv007 <= Z018v6;
always @(posedge HCLK) Pvv007 <= S018v6;
always @(posedge HCLK) Gyv007 <= L018v6;
always @(posedge HCLK) X0w007 <= E018v6;
always @(posedge HCLK) O3w007 <= Xz08v6;
always @(posedge HCLK) F6w007 <= Qz08v6;
always @(posedge HCLK) W8w007 <= Jz08v6;
always @(posedge HCLK) Nbw007 <= Cz08v6;
always @(posedge HCLK) Eew007 <= Vy08v6;
always @(posedge HCLK) Vgw007 <= Oy08v6;
always @(posedge HCLK) Mjw007 <= Hy08v6;
always @(posedge HCLK) Dmw007 <= Ay08v6;
always @(posedge HCLK) Uow007 <= Tx08v6;
always @(posedge HCLK) Lrw007 <= Mx08v6;
always @(posedge HCLK) Cuw007 <= Fx08v6;
always @(posedge HCLK) Tww007 <= Yw08v6;
always @(posedge HCLK) Kzw007 <= Rw08v6;
always @(posedge HCLK) B2x007 <= Kw08v6;
always @(posedge HCLK) S4x007 <= Dw08v6;
always @(posedge HCLK) J7x007 <= Wv08v6;
always @(posedge HCLK) Z9x007 <= Pv08v6;
always @(posedge HCLK) Pcx007 <= Iv08v6;
always @(posedge HCLK) Ffx007 <= Bv08v6;
always @(posedge HCLK) Vhx007 <= Uu08v6;
always @(posedge HCLK) Lkx007 <= Nu08v6;
always @(posedge HCLK) Bnx007 <= Gu08v6;
always @(posedge HCLK) Rpx007 <= Zt08v6;
always @(posedge HCLK) Hsx007 <= St08v6;
always @(posedge HCLK) Xux007 <= Jmz7v6;
always @(posedge HCLK) Nxx007 <= Cmz7v6;
always @(posedge HCLK) E0y007 <= Vlz7v6;
always @(posedge HCLK) V2y007 <= Olz7v6;
always @(posedge HCLK) M5y007 <= Hlz7v6;
always @(posedge HCLK) D8y007 <= Alz7v6;
always @(posedge HCLK) Uay007 <= Tkz7v6;
always @(posedge HCLK) Ldy007 <= Mkz7v6;
always @(posedge HCLK) Cgy007 <= Fkz7v6;
always @(posedge HCLK) Tiy007 <= Yjz7v6;
always @(posedge HCLK) Kly007 <= Rjz7v6;
always @(posedge HCLK) Boy007 <= Kjz7v6;
always @(posedge HCLK) Sqy007 <= Djz7v6;
always @(posedge HCLK) Jty007 <= Wiz7v6;
always @(posedge HCLK) Awy007 <= Piz7v6;
always @(posedge HCLK) Ryy007 <= Iiz7v6;
always @(posedge HCLK) I1z007 <= Biz7v6;
always @(posedge HCLK) Z3z007 <= Uhz7v6;
always @(posedge HCLK) Q6z007 <= Nhz7v6;
always @(posedge HCLK) H9z007 <= Ghz7v6;
always @(posedge HCLK) Ybz007 <= Zgz7v6;
always @(posedge HCLK) Pez007 <= Sgz7v6;
always @(posedge HCLK) Ghz007 <= Lgz7v6;
always @(posedge HCLK) Wjz007 <= Egz7v6;
always @(posedge HCLK) Mmz007 <= Xfz7v6;
always @(posedge HCLK) Cpz007 <= Qfz7v6;
always @(posedge HCLK) Srz007 <= Jfz7v6;
always @(posedge HCLK) Iuz007 <= Cfz7v6;
always @(posedge HCLK) Ywz007 <= Vez7v6;
always @(posedge HCLK) Ozz007 <= Oez7v6;
always @(posedge HCLK) E20107 <= Hez7v6;
always @(posedge HCLK) U40107 <= O3p7v6;
always @(posedge HCLK) Y70107 <= Vnx7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qa0107 <= 1'b0;
  else
    Qa0107 <= D2g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Lc0107 <= 1'b0;
  else
    Lc0107 <= W1g8v6;

always @(posedge HCLK) De0107 <= Mks7v6;
always @(posedge HCLK) Sg0107 <= W8o7v6;
always @(posedge HCLK) Wj0107 <= Y9o7v6;
always @(posedge HCLK) An0107 <= Iis7v6;
always @(posedge HCLK) Pp0107 <= Rlx7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hs0107 <= 1'b0;
  else
    Hs0107 <= Vxf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Cu0107 <= 1'b0;
  else
    Cu0107 <= Oxf8v6;

always @(posedge HCLK) Uv0107 <= Trs7v6;
always @(posedge HCLK) Yy0107 <= Ass7v6;
always @(posedge HCLK) C21107 <= Bis7v6;
always @(posedge HCLK) R41107 <= Ylx7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    J71107 <= 1'b0;
  else
    J71107 <= Jyf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    E91107 <= 1'b0;
  else
    E91107 <= Cyf8v6;

always @(posedge HCLK) Wa1107 <= Hss7v6;
always @(posedge HCLK) Ae1107 <= Oss7v6;
always @(posedge HCLK) Eh1107 <= Uhs7v6;
always @(posedge HCLK) Tj1107 <= Fmx7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lm1107 <= 1'b0;
  else
    Lm1107 <= Xyf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Go1107 <= 1'b0;
  else
    Go1107 <= Qyf8v6;

always @(posedge HCLK) Yp1107 <= Vss7v6;
always @(posedge HCLK) Ct1107 <= Cts7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gw1107 <= 1'b0;
  else
    Gw1107 <= Nij8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ez1107 <= 1'b0;
  else
    Ez1107 <= Gij8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L12107 <= 1'b0;
  else
    L12107 <= Tzj8v6;

always @(posedge HCLK) S32107 <= Hap7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V62107 <= 1'b0;
  else
    V62107 <= Upj8v6;

always @(posedge HCLK) U92107 <= Z5p7v6;
always @(posedge HCLK) Yc2107 <= Nhs7v6;
always @(posedge HCLK) Nf2107 <= Mmx7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fi2107 <= 1'b0;
  else
    Fi2107 <= Lzf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ak2107 <= 1'b0;
  else
    Ak2107 <= Ezf8v6;

always @(posedge HCLK) Sl2107 <= Jts7v6;
always @(posedge HCLK) Wo2107 <= Qts7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    As2107 <= 1'b0;
  else
    As2107 <= Zhj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yu2107 <= 1'b0;
  else
    Yu2107 <= Ktw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xx2107 <= 1'b0;
  else
    Xx2107 <= Urw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W03107 <= 1'b0;
  else
    W03107 <= Bsw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V33107 <= 1'b0;
  else
    V33107 <= Isw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U63107 <= 1'b0;
  else
    U63107 <= Psw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T93107 <= 1'b0;
  else
    T93107 <= Wsw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sc3107 <= 1'b0;
  else
    Sc3107 <= Dtw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rf3107 <= 1'b0;
  else
    Rf3107 <= Vo38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sh3107 <= 1'b0;
  else
    Sh3107 <= Uwj8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sj3107 <= 1'b0;
  else
    Sj3107 <= Fwu7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yl3107 <= 1'b0;
  else
    Yl3107 <= Qgj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fo3107 <= 1'b0;
  else
    Fo3107 <= Fej8v6;

always @(posedge HCLK) Oq3107 <= Oap7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rt3107 <= 1'b0;
  else
    Rt3107 <= Npj8v6;

always @(posedge HCLK) Qw3107 <= P6i8v6;
always @(posedge HCLK) Wy3107 <= L4i8v6;
always @(posedge HCLK) C14107 <= O2i8v6;
always @(posedge HCLK) H34107 <= W6i8v6;
always @(posedge HCLK) N54107 <= S4i8v6;
always @(posedge HCLK) T74107 <= V2i8v6;
always @(posedge HCLK) Z94107 <= D7i8v6;
always @(posedge HCLK) Fc4107 <= Z4i8v6;
always @(posedge HCLK) Le4107 <= C3i8v6;
always @(posedge HCLK) Rg4107 <= G5i8v6;
always @(posedge HCLK) Xi4107 <= U5i8v6;
always @(posedge HCLK) Dl4107 <= Q3i8v6;
always @(posedge HCLK) Jn4107 <= B6i8v6;
always @(posedge HCLK) Pp4107 <= X3i8v6;
always @(posedge HCLK) Vr4107 <= I6i8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bu4107 <= 1'b0;
  else
    Bu4107 <= Y6j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ax4107 <= 1'b0;
  else
    Ax4107 <= O8j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xz4107 <= 1'b0;
  else
    Xz4107 <= H8j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U25107 <= 1'b0;
  else
    U25107 <= Zaj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L55107 <= 1'b0;
  else
    L55107 <= Wu88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    I85107 <= 1'b0;
  else
    I85107 <= R6j8v6;

always @(posedge HCLK) Ka5107 <= Qwh8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yc5107 <= 1'b0;
  else
    Yc5107 <= Vui8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wf5107 <= 1'b0;
  else
    Wf5107 <= Lwi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ui5107 <= 1'b0;
  else
    Ui5107 <= Ewi8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kl5107 <= 1'b0;
  else
    Kl5107 <= Ksx7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    En5107 <= 1'b0;
  else
    En5107 <= Rsx7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yo5107 <= 1'b1;
  else
    Yo5107 <= Xvx7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Oq5107 <= 1'b0;
  else
    Oq5107 <= Ewx7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Is5107 <= 1'b1;
  else
    Is5107 <= Ttx7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yt5107 <= 1'b1;
  else
    Yt5107 <= Oux7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ov5107 <= 1'b0;
  else
    Ov5107 <= Jel8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bx5107 <= 1'b1;
  else
    Bx5107 <= Qvx7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ry5107 <= 1'b1;
  else
    Ry5107 <= Jvx7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    I06107 <= 1'b1;
  else
    I06107 <= Cvx7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Z16107 <= 1'b1;
  else
    Z16107 <= Vux7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    P36107 <= 1'b1;
  else
    P36107 <= Hux7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F56107 <= 1'b1;
  else
    F56107 <= Aux7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    V66107 <= 1'b1;
  else
    V66107 <= Mtx7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    L86107 <= 1'b1;
  else
    L86107 <= Ftx7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ba6107 <= 1'b1;
  else
    Ba6107 <= Prx7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rb6107 <= 1'b0;
  else
    Rb6107 <= Gf88v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gd6107 <= 1'b0;
  else
    Gd6107 <= Ze88v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ve6107 <= 1'b0;
  else
    Ve6107 <= Se88v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kg6107 <= 1'b0;
  else
    Kg6107 <= Le88v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yh6107 <= 1'b0;
  else
    Yh6107 <= Ee88v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lj6107 <= 1'b0;
  else
    Lj6107 <= Nu78v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fl6107 <= 1'b0;
  else
    Fl6107 <= U3k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zn6107 <= 1'b0;
  else
    Zn6107 <= Uc48v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Br6107 <= 1'b0;
  else
    Br6107 <= Bd48v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Du6107 <= 1'b0;
  else
    Du6107 <= Zwi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bx6107 <= 1'b0;
  else
    Bx6107 <= Swi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vz6107 <= 1'b0;
  else
    Vz6107 <= Gxi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U27107 <= 1'b0;
  else
    U27107 <= D6j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T57107 <= 1'b0;
  else
    T57107 <= Pcy7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V87107 <= 1'b0;
  else
    V87107 <= D838v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xb7107 <= 1'b0;
  else
    Xb7107 <= F7j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    We7107 <= 1'b0;
  else
    We7107 <= Mej8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dh7107 <= 1'b0;
  else
    Dh7107 <= Hfj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kj7107 <= 1'b0;
  else
    Kj7107 <= Ofj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rl7107 <= 1'b0;
  else
    Rl7107 <= Ehj8v6;

always @(posedge HCLK) Yn7107 <= J3i8v6;
always @(posedge HCLK) Eq7107 <= N5i8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ks7107 <= 1'b0;
  else
    Ks7107 <= Wdi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lu7107 <= 1'b0;
  else
    Lu7107 <= Shj8v6;

always @(posedge HCLK) Qw7107 <= Pzh8v6;
always @(posedge HCLK) Qz7107 <= Izh8v6;
always @(posedge HCLK) Q28107 <= Bzh8v6;
always @(posedge HCLK) Q58107 <= Uyh8v6;
always @(posedge HCLK) Q88107 <= Nyh8v6;
always @(posedge HCLK) Gttf07 <= Gyh8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gwtf07 <= 1'b0;
  else
    Gwtf07 <= Cvi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Eztf07 <= 1'b0;
  else
    Eztf07 <= M7j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    G2uf07 <= 1'b0;
  else
    G2uf07 <= W5j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    G5uf07 <= 1'b0;
  else
    G5uf07 <= J9j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J8uf07 <= 1'b0;
  else
    J8uf07 <= Q9j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mbuf07 <= 1'b0;
  else
    Mbuf07 <= X9j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Peuf07 <= 1'b0;
  else
    Peuf07 <= Ogi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ahuf07 <= 1'b0;
  else
    Ahuf07 <= Mfi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xjuf07 <= 1'b0;
  else
    Xjuf07 <= Ffi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Umuf07 <= 1'b0;
  else
    Umuf07 <= Tfi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fpuf07 <= 1'b0;
  else
    Fpuf07 <= Xhi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Csuf07 <= 1'b0;
  else
    Csuf07 <= Kei8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zuuf07 <= 1'b0;
  else
    Zuuf07 <= Hgi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kxuf07 <= 1'b0;
  else
    Kxuf07 <= Vgi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H0vf07 <= 1'b0;
  else
    H0vf07 <= Yei8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    E3vf07 <= 1'b0;
  else
    E3vf07 <= Hui8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B6vf07 <= 1'b0;
  else
    B6vf07 <= Xgj8v6;

always @(posedge HCLK) I8vf07 <= G6p7v6;
always @(posedge HCLK) Mbvf07 <= Ghs7v6;
always @(posedge HCLK) Bevf07 <= Tmx7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tgvf07 <= 1'b0;
  else
    Tgvf07 <= Zzf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Oivf07 <= 1'b0;
  else
    Oivf07 <= Szf8v6;

always @(posedge HCLK) Gkvf07 <= Xts7v6;
always @(posedge HCLK) Knvf07 <= Eus7v6;
always @(posedge HCLK) Oqvf07 <= Zgs7v6;
always @(posedge HCLK) Dtvf07 <= Anx7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vvvf07 <= 1'b0;
  else
    Vvvf07 <= N0g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Qxvf07 <= 1'b0;
  else
    Qxvf07 <= G0g8v6;

always @(posedge HCLK) Izvf07 <= Lus7v6;
always @(posedge HCLK) M2wf07 <= Sus7v6;
always @(posedge HCLK) Q5wf07 <= Lgs7v6;
always @(posedge HCLK) F8wf07 <= Klx7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xawf07 <= 1'b0;
  else
    Xawf07 <= P1g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Scwf07 <= 1'b0;
  else
    Scwf07 <= I1g8v6;

always @(posedge HCLK) Kewf07 <= I7p7v6;
always @(posedge HCLK) Ohwf07 <= Nvs7v6;
always @(posedge HCLK) Skwf07 <= D9o7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wnwf07 <= 1'b0;
  else
    Wnwf07 <= B898v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lqwf07 <= 1'b0;
  else
    Lqwf07 <= Spnet6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ltwf07 <= 1'b0;
  else
    Ltwf07 <= Gbj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jwwf07 <= 1'b0;
  else
    Jwwf07 <= Nbj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hzwf07 <= 1'b0;
  else
    Hzwf07 <= Tzc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D2xf07 <= 1'b0;
  else
    D2xf07 <= Qvi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D5xf07 <= 1'b0;
  else
    D5xf07 <= Xvi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    A8xf07 <= 1'b0;
  else
    A8xf07 <= O6l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uaxf07 <= 1'b0;
  else
    Uaxf07 <= Fds7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Udxf07 <= 1'b0;
  else
    Udxf07 <= Zxh8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ngxf07 <= 1'b0;
  else
    Ngxf07 <= Ydj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wixf07 <= 1'b0;
  else
    Wixf07 <= Icj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xkxf07 <= 1'b0;
  else
    Xkxf07 <= Bcj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Unxf07 <= 1'b0;
  else
    Unxf07 <= Lhj8v6;

always @(posedge HCLK) Bqxf07 <= K7i8v6;
always @(posedge HCLK) Hsxf07 <= R7i8v6;
always @(posedge HCLK) Nuxf07 <= Y7i8v6;
always @(posedge HCLK) Twxf07 <= F8i8v6;
always @(posedge HCLK) Zyxf07 <= M8i8v6;
always @(posedge HCLK) F1yf07 <= K0i8v6;
always @(posedge HCLK) K3yf07 <= A2i8v6;
always @(posedge HCLK) P5yf07 <= T1i8v6;
always @(posedge HCLK) U7yf07 <= Aap7v6;
always @(posedge HCLK) Xayf07 <= Wto7v6;
always @(posedge HCLK) Ndyf07 <= Zs88v6;
always @(posedge HCLK) Dgyf07 <= Ss88v6;
always @(posedge HCLK) Tiyf07 <= Ls88v6;
always @(posedge HCLK) Jlyf07 <= Es88v6;
always @(posedge HCLK) Znyf07 <= Xr88v6;
always @(posedge HCLK) Pqyf07 <= Qr88v6;
always @(posedge HCLK) Ftyf07 <= Ck88v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tvyf07 <= 1'b0;
  else
    Tvyf07 <= Tsj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xyyf07 <= 1'b0;
  else
    Xyyf07 <= Otj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B2zf07 <= 1'b0;
  else
    B2zf07 <= Qp38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    E5zf07 <= 1'b0;
  else
    E5zf07 <= K4l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    I8zf07 <= 1'b0;
  else
    I8zf07 <= A7k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nazf07 <= 1'b0;
  else
    Nazf07 <= H7k8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sczf07 <= 1'b0;
  else
    Sczf07 <= Bam7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tfzf07 <= 1'b0;
  else
    Tfzf07 <= Icy7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Thzf07 <= 1'b0;
  else
    Thzf07 <= Uhk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vjzf07 <= 1'b0;
  else
    Vjzf07 <= Kof8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lmzf07 <= 1'b0;
  else
    Lmzf07 <= S9k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fozf07 <= 1'b1;
  else
    Fozf07 <= Hcf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zqzf07 <= 1'b0;
  else
    Zqzf07 <= Acf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ptzf07 <= 1'b0;
  else
    Ptzf07 <= U8f8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Owzf07 <= 1'b0;
  else
    Owzf07 <= Nf88v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Byzf07 <= 1'b0;
  else
    Byzf07 <= Cs78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yzzf07 <= 1'b0;
  else
    Yzzf07 <= Gu78v6;

always @(posedge HCLK) M10g07 <= U9m7v6;
always @(posedge HCLK) C30g07 <= N9m7v6;
always @(posedge HCLK) S40g07 <= G9m7v6;
always @(posedge HCLK) H60g07 <= Z8m7v6;
always @(posedge HCLK) W70g07 <= S8m7v6;
always @(posedge HCLK) L90g07 <= L8m7v6;
always @(posedge HCLK) Ab0g07 <= E8m7v6;
always @(posedge HCLK) Pc0g07 <= X7m7v6;
always @(posedge HCLK) Ee0g07 <= Q7m7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tf0g07 <= 1'b0;
  else
    Tf0g07 <= J7m7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zg0g07 <= 1'b0;
  else
    Zg0g07 <= C7m7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fi0g07 <= 1'b0;
  else
    Fi0g07 <= V6m7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lj0g07 <= 1'b0;
  else
    Lj0g07 <= O6m7v6;

always @(posedge HCLK) Rk0g07 <= H6m7v6;
always @(posedge HCLK) Om0g07 <= A6m7v6;
always @(posedge HCLK) Lo0g07 <= T5m7v6;
always @(posedge HCLK) Iq0g07 <= M5m7v6;
always @(posedge HCLK) Fs0g07 <= F5m7v6;
always @(posedge HCLK) Cu0g07 <= Y4m7v6;
always @(posedge HCLK) Zv0g07 <= R4m7v6;
always @(posedge HCLK) Wx0g07 <= K4m7v6;
always @(posedge HCLK) Uz0g07 <= D4m7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    S11g07 <= 1'b0;
  else
    S11g07 <= T3g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    N31g07 <= 1'b0;
  else
    N31g07 <= M3g8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    F51g07 <= 1'b0;
  else
    F51g07 <= Yof8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    G71g07 <= 1'b0;
  else
    G71g07 <= Syg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    V81g07 <= 1'b0;
  else
    V81g07 <= Lyg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Ka1g07 <= 1'b0;
  else
    Ka1g07 <= Eyg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Zb1g07 <= 1'b0;
  else
    Zb1g07 <= Xxg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Od1g07 <= 1'b0;
  else
    Od1g07 <= Qxg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Df1g07 <= 1'b0;
  else
    Df1g07 <= Vwg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Pg1g07 <= 1'b0;
  else
    Pg1g07 <= Tog8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Qi1g07 <= 1'b0;
  else
    Qi1g07 <= Mog8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Rk1g07 <= 1'b1;
  else
    Rk1g07 <= Fgh8v6;

always @(posedge HCLK) Mm1g07 <= Als7v6;
always @(posedge HCLK) Ap1g07 <= Re48v6;
always @(posedge HCLK) Ds1g07 <= Ye48v6;
always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Gv1g07 <= 1'b0;
  else
    Gv1g07 <= Vw47v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Uw1g07 <= 1'b0;
  else
    Uw1g07 <= Glg8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Iy1g07 <= 1'b0;
  else
    Iy1g07 <= X767v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Xz1g07 <= 1'b0;
  else
    Xz1g07 <= Rug8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L12g07 <= 1'b0;
  else
    L12g07 <= N798v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    C42g07 <= 1'b0;
  else
    C42g07 <= Obo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T62g07 <= 1'b0;
  else
    T62g07 <= G798v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M92g07 <= 1'b0;
  else
    M92g07 <= Z698v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fc2g07 <= 1'b0;
  else
    Fc2g07 <= S698v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ye2g07 <= 1'b0;
  else
    Ye2g07 <= L698v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rh2g07 <= 1'b0;
  else
    Rh2g07 <= E698v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lk2g07 <= 1'b0;
  else
    Lk2g07 <= X598v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fn2g07 <= 1'b0;
  else
    Fn2g07 <= Q598v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zp2g07 <= 1'b0;
  else
    Zp2g07 <= J598v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ts2g07 <= 1'b0;
  else
    Ts2g07 <= C598v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nv2g07 <= 1'b0;
  else
    Nv2g07 <= V498v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hy2g07 <= 1'b0;
  else
    Hy2g07 <= O498v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B13g07 <= 1'b0;
  else
    B13g07 <= H498v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V33g07 <= 1'b0;
  else
    V33g07 <= A498v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P63g07 <= 1'b0;
  else
    P63g07 <= T398v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J93g07 <= 1'b0;
  else
    J93g07 <= M398v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dc3g07 <= 1'b0;
  else
    Dc3g07 <= F398v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xe3g07 <= 1'b0;
  else
    Xe3g07 <= Y298v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rh3g07 <= 1'b0;
  else
    Rh3g07 <= R298v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lk3g07 <= 1'b0;
  else
    Lk3g07 <= K298v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fn3g07 <= 1'b0;
  else
    Fn3g07 <= D298v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zp3g07 <= 1'b0;
  else
    Zp3g07 <= W198v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ts3g07 <= 1'b0;
  else
    Ts3g07 <= P198v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nv3g07 <= 1'b0;
  else
    Nv3g07 <= I198v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hy3g07 <= 1'b0;
  else
    Hy3g07 <= B198v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B14g07 <= 1'b0;
  else
    B14g07 <= U098v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V34g07 <= 1'b0;
  else
    V34g07 <= G098v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    O64g07 <= 1'b0;
  else
    O64g07 <= A9i8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    S84g07 <= 1'b0;
  else
    S84g07 <= Nwj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ra4g07 <= 1'b0;
  else
    Ra4g07 <= Bdi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tc4g07 <= 1'b0;
  else
    Tc4g07 <= Tej8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Af4g07 <= 1'b0;
  else
    Af4g07 <= Aa38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yh4g07 <= 1'b0;
  else
    Yh4g07 <= Qi38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xk4g07 <= 1'b0;
  else
    Xk4g07 <= Ha38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vn4g07 <= 1'b0;
  else
    Vn4g07 <= Oa38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tq4g07 <= 1'b0;
  else
    Tq4g07 <= Va38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rt4g07 <= 1'b0;
  else
    Rt4g07 <= Jb38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pw4g07 <= 1'b0;
  else
    Pw4g07 <= Qb38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oz4g07 <= 1'b0;
  else
    Oz4g07 <= Xb38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N25g07 <= 1'b0;
  else
    N25g07 <= Ec38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M55g07 <= 1'b0;
  else
    M55g07 <= Bl38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L85g07 <= 1'b0;
  else
    L85g07 <= Pl38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kb5g07 <= 1'b0;
  else
    Kb5g07 <= T938v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ie5g07 <= 1'b0;
  else
    Ie5g07 <= Wl38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gh5g07 <= 1'b0;
  else
    Gh5g07 <= Dm38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bk5g07 <= 1'b0;
  else
    Bk5g07 <= Km38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ym5g07 <= 1'b0;
  else
    Ym5g07 <= Il38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xp5g07 <= 1'b0;
  else
    Xp5g07 <= Xi38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ws5g07 <= 1'b0;
  else
    Ws5g07 <= Ji38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vv5g07 <= 1'b0;
  else
    Vv5g07 <= Ci38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uy5g07 <= 1'b0;
  else
    Uy5g07 <= Vh38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T16g07 <= 1'b0;
  else
    T16g07 <= Qhi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W46g07 <= 1'b0;
  else
    W46g07 <= Iik8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z76g07 <= 1'b0;
  else
    Z76g07 <= Oui8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xa6g07 <= 1'b0;
  else
    Xa6g07 <= Dei8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ae6g07 <= 1'b0;
  else
    Ae6g07 <= Cb38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yg6g07 <= 1'b0;
  else
    Yg6g07 <= M938v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wj6g07 <= 1'b0;
  else
    Wj6g07 <= K838v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xm6g07 <= 1'b0;
  else
    Xm6g07 <= R838v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yp6g07 <= 1'b0;
  else
    Yp6g07 <= F938v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zs6g07 <= 1'b0;
  else
    Zs6g07 <= Afj8v6;

always @(posedge HCLK) Gv6g07 <= B7p7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ky6g07 <= 1'b1;
  else
    Ky6g07 <= W3m7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    T07g07 <= 1'b0;
  else
    T07g07 <= Rjzet6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    H37g07 <= 1'b0;
  else
    H37g07 <= Ay0ft6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P57g07 <= 1'b0;
  else
    P57g07 <= Pd48v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R87g07 <= 1'b0;
  else
    R87g07 <= Gc48v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tb7g07 <= 1'b0;
  else
    Tb7g07 <= Nc48v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ve7g07 <= 1'b0;
  else
    Ve7g07 <= Wd48v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xh7g07 <= 1'b0;
  else
    Xh7g07 <= Yhf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ak7g07 <= 1'b0;
  else
    Ak7g07 <= Fif8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dm7g07 <= 1'b0;
  else
    Dm7g07 <= Mif8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Go7g07 <= 1'b0;
  else
    Go7g07 <= Tif8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jq7g07 <= 1'b0;
  else
    Jq7g07 <= Ckf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ss7g07 <= 1'b0;
  else
    Ss7g07 <= Xkf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bv7g07 <= 1'b0;
  else
    Bv7g07 <= Llf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lx7g07 <= 1'b0;
  else
    Lx7g07 <= Slf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vz7g07 <= 1'b0;
  else
    Vz7g07 <= Gmf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    V18g07 <= 1'b0;
  else
    V18g07 <= Zlf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    E48g07 <= 1'b0;
  else
    E48g07 <= Elf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    N68g07 <= 1'b0;
  else
    N68g07 <= Qkf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    W88g07 <= 1'b0;
  else
    W88g07 <= Jkf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fb8g07 <= 1'b0;
  else
    Fb8g07 <= P3m7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kd8g07 <= 1'b0;
  else
    Kd8g07 <= I3m7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pf8g07 <= 1'b0;
  else
    Pf8g07 <= B3m7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uh8g07 <= 1'b0;
  else
    Uh8g07 <= U2m7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zj8g07 <= 1'b0;
  else
    Zj8g07 <= N2m7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Em8g07 <= 1'b0;
  else
    Em8g07 <= G2m7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jo8g07 <= 1'b0;
  else
    Jo8g07 <= Z1m7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oq8g07 <= 1'b0;
  else
    Oq8g07 <= S1m7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ts8g07 <= 1'b0;
  else
    Ts8g07 <= L1m7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yu8g07 <= 1'b0;
  else
    Yu8g07 <= E1m7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dx8g07 <= 1'b0;
  else
    Dx8g07 <= X0m7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Iz8g07 <= 1'b0;
  else
    Iz8g07 <= Q0m7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N19g07 <= 1'b0;
  else
    N19g07 <= J0m7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    S39g07 <= 1'b0;
  else
    S39g07 <= C0m7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W59g07 <= 1'b0;
  else
    W59g07 <= Vzl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    A89g07 <= 1'b0;
  else
    A89g07 <= Ozl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ea9g07 <= 1'b0;
  else
    Ea9g07 <= Hzl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ic9g07 <= 1'b0;
  else
    Ic9g07 <= Azl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Me9g07 <= 1'b0;
  else
    Me9g07 <= Tyl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qg9g07 <= 1'b0;
  else
    Qg9g07 <= Myl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ui9g07 <= 1'b0;
  else
    Ui9g07 <= Fyl7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yk9g07 <= 1'b0;
  else
    Yk9g07 <= Vjf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hn9g07 <= 1'b0;
  else
    Hn9g07 <= Ojf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qp9g07 <= 1'b0;
  else
    Qp9g07 <= Yxl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sr9g07 <= 1'b0;
  else
    Sr9g07 <= Rxl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ut9g07 <= 1'b0;
  else
    Ut9g07 <= Kxl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wv9g07 <= 1'b0;
  else
    Wv9g07 <= Dxl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zx9g07 <= 1'b0;
  else
    Zx9g07 <= Wwl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    C0ag07 <= 1'b0;
  else
    C0ag07 <= Pwl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F2ag07 <= 1'b0;
  else
    F2ag07 <= Iwl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H4ag07 <= 1'b0;
  else
    H4ag07 <= Bwl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J6ag07 <= 1'b0;
  else
    J6ag07 <= Uvl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L8ag07 <= 1'b0;
  else
    L8ag07 <= B4d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Paag07 <= 1'b0;
  else
    Paag07 <= X8d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tcag07 <= 1'b0;
  else
    Tcag07 <= Tdd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xeag07 <= 1'b0;
  else
    Xeag07 <= Znd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bhag07 <= 1'b0;
  else
    Bhag07 <= Vsd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gjag07 <= 1'b0;
  else
    Gjag07 <= Rxd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Llag07 <= 1'b0;
  else
    Llag07 <= J7e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qnag07 <= 1'b0;
  else
    Qnag07 <= Fce8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vpag07 <= 1'b0;
  else
    Vpag07 <= U1f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Asag07 <= 1'b0;
  else
    Asag07 <= Q6f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fuag07 <= 1'b0;
  else
    Fuag07 <= Nff8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kwag07 <= 1'b0;
  else
    Kwag07 <= X1d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nyag07 <= 1'b0;
  else
    Nyag07 <= T6d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q0bg07 <= 1'b0;
  else
    Q0bg07 <= Pbd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T2bg07 <= 1'b0;
  else
    T2bg07 <= Vld8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W4bg07 <= 1'b0;
  else
    W4bg07 <= Rqd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z6bg07 <= 1'b0;
  else
    Z6bg07 <= Nvd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    C9bg07 <= 1'b0;
  else
    C9bg07 <= F5e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fbbg07 <= 1'b0;
  else
    Fbbg07 <= Bae8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Idbg07 <= 1'b0;
  else
    Idbg07 <= Qze8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lfbg07 <= 1'b0;
  else
    Lfbg07 <= M4f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Phbg07 <= 1'b0;
  else
    Phbg07 <= Rhf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tjbg07 <= 1'b0;
  else
    Tjbg07 <= I4d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ylbg07 <= 1'b0;
  else
    Ylbg07 <= E9d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dobg07 <= 1'b0;
  else
    Dobg07 <= Aed8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Iqbg07 <= 1'b0;
  else
    Iqbg07 <= God8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nsbg07 <= 1'b0;
  else
    Nsbg07 <= Ctd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Subg07 <= 1'b0;
  else
    Subg07 <= Yxd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xwbg07 <= 1'b0;
  else
    Xwbg07 <= Q7e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Czbg07 <= 1'b0;
  else
    Czbg07 <= Mce8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H1cg07 <= 1'b0;
  else
    H1cg07 <= B2f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M3cg07 <= 1'b0;
  else
    M3cg07 <= X6f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R5cg07 <= 1'b0;
  else
    R5cg07 <= Gff8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W7cg07 <= 1'b0;
  else
    W7cg07 <= E2d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Aacg07 <= 1'b0;
  else
    Aacg07 <= A7d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Eccg07 <= 1'b0;
  else
    Eccg07 <= Wbd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Iecg07 <= 1'b0;
  else
    Iecg07 <= Cmd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mgcg07 <= 1'b0;
  else
    Mgcg07 <= Yqd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qicg07 <= 1'b0;
  else
    Qicg07 <= Uvd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ukcg07 <= 1'b0;
  else
    Ukcg07 <= M5e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ymcg07 <= 1'b0;
  else
    Ymcg07 <= Iae8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cpcg07 <= 1'b0;
  else
    Cpcg07 <= Xze8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Grcg07 <= 1'b0;
  else
    Grcg07 <= T4f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ktcg07 <= 1'b0;
  else
    Ktcg07 <= Khf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ovcg07 <= 1'b0;
  else
    Ovcg07 <= Nvl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nxcg07 <= 1'b0;
  else
    Nxcg07 <= Gvl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mzcg07 <= 1'b0;
  else
    Mzcg07 <= Rh88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P1dg07 <= 1'b0;
  else
    P1dg07 <= Pxc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    S3dg07 <= 1'b0;
  else
    S3dg07 <= Fzc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V5dg07 <= 1'b0;
  else
    V5dg07 <= A0d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y7dg07 <= 1'b0;
  else
    Y7dg07 <= J1d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Badg07 <= 1'b0;
  else
    Badg07 <= F6d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ecdg07 <= 1'b0;
  else
    Ecdg07 <= Bbd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hedg07 <= 1'b0;
  else
    Hedg07 <= Pid8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kgdg07 <= 1'b0;
  else
    Kgdg07 <= Kjd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nidg07 <= 1'b0;
  else
    Nidg07 <= Fkd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qkdg07 <= 1'b0;
  else
    Qkdg07 <= Tkd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tmdg07 <= 1'b0;
  else
    Tmdg07 <= Hld8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wodg07 <= 1'b0;
  else
    Wodg07 <= Dqd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zqdg07 <= 1'b0;
  else
    Zqdg07 <= Zud8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ctdg07 <= 1'b0;
  else
    Ctdg07 <= Fje8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fvdg07 <= 1'b0;
  else
    Fvdg07 <= Ywe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ixdg07 <= 1'b0;
  else
    Ixdg07 <= Mxe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lzdg07 <= 1'b0;
  else
    Lzdg07 <= Aye8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O1eg07 <= 1'b0;
  else
    O1eg07 <= Oye8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R3eg07 <= 1'b0;
  else
    R3eg07 <= Cze8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U5eg07 <= 1'b0;
  else
    U5eg07 <= Y3f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X7eg07 <= 1'b0;
  else
    X7eg07 <= Jdf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Aaeg07 <= 1'b0;
  else
    Aaeg07 <= N2e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dceg07 <= 1'b0;
  else
    Dceg07 <= B3e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Geeg07 <= 1'b0;
  else
    Geeg07 <= P3e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jgeg07 <= 1'b0;
  else
    Jgeg07 <= D4e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mieg07 <= 1'b0;
  else
    Mieg07 <= R4e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pkeg07 <= 1'b0;
  else
    Pkeg07 <= N9e8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Smeg07 <= 1'b0;
  else
    Smeg07 <= Yjk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qpeg07 <= 1'b0;
  else
    Qpeg07 <= Zul7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rseg07 <= 1'b0;
  else
    Rseg07 <= Sul7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vueg07 <= 1'b0;
  else
    Vueg07 <= Lul7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xweg07 <= 1'b0;
  else
    Xweg07 <= Lef8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Czeg07 <= 1'b0;
  else
    Czeg07 <= S7f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H1fg07 <= 1'b0;
  else
    H1fg07 <= W2f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M3fg07 <= 1'b0;
  else
    M3fg07 <= Hde8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R5fg07 <= 1'b0;
  else
    R5fg07 <= L8e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W7fg07 <= 1'b0;
  else
    W7fg07 <= Tyd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bafg07 <= 1'b0;
  else
    Bafg07 <= Xtd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gcfg07 <= 1'b0;
  else
    Gcfg07 <= Bpd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lefg07 <= 1'b0;
  else
    Lefg07 <= Ved8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qgfg07 <= 1'b0;
  else
    Qgfg07 <= Z9d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vifg07 <= 1'b0;
  else
    Vifg07 <= D5d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Alfg07 <= 1'b0;
  else
    Alfg07 <= Pgf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Enfg07 <= 1'b0;
  else
    Enfg07 <= O5f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ipfg07 <= 1'b0;
  else
    Ipfg07 <= S0f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mrfg07 <= 1'b0;
  else
    Mrfg07 <= Dbe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qtfg07 <= 1'b0;
  else
    Qtfg07 <= H6e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uvfg07 <= 1'b0;
  else
    Uvfg07 <= Pwd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yxfg07 <= 1'b0;
  else
    Yxfg07 <= Trd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    C0gg07 <= 1'b0;
  else
    C0gg07 <= Xmd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    G2gg07 <= 1'b0;
  else
    G2gg07 <= Rcd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K4gg07 <= 1'b0;
  else
    K4gg07 <= V7d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O6gg07 <= 1'b0;
  else
    O6gg07 <= Z2d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    S8gg07 <= 1'b0;
  else
    S8gg07 <= Eul7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pagg07 <= 1'b0;
  else
    Pagg07 <= Xtl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qcgg07 <= 1'b0;
  else
    Qcgg07 <= C4w7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oegg07 <= 1'b0;
  else
    Oegg07 <= Ajf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tggg07 <= 1'b1;
  else
    Tggg07 <= Qtl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bjgg07 <= 1'b0;
  else
    Bjgg07 <= F6k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Klgg07 <= 1'b0;
  else
    Klgg07 <= Bbk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ongg07 <= 1'b1;
  else
    Ongg07 <= Uak8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cqgg07 <= 1'b0;
  else
    Cqgg07 <= Jtl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jsgg07 <= 1'b0;
  else
    Jsgg07 <= Ctl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qugg07 <= 1'b0;
  else
    Qugg07 <= Vsl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xwgg07 <= 1'b0;
  else
    Xwgg07 <= Osl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ezgg07 <= 1'b0;
  else
    Ezgg07 <= C9j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B2hg07 <= 1'b0;
  else
    B2hg07 <= V8j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y4hg07 <= 1'b0;
  else
    Y4hg07 <= Hsl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F7hg07 <= 1'b0;
  else
    F7hg07 <= Asl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M9hg07 <= 1'b0;
  else
    M9hg07 <= Trl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pbhg07 <= 1'b0;
  else
    Pbhg07 <= Mrl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sdhg07 <= 1'b0;
  else
    Sdhg07 <= Frl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vfhg07 <= 1'b0;
  else
    Vfhg07 <= Icc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rhhg07 <= 1'b0;
  else
    Rhhg07 <= Pcc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Njhg07 <= 1'b0;
  else
    Njhg07 <= Ddc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jlhg07 <= 1'b0;
  else
    Jlhg07 <= Kdc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fnhg07 <= 1'b0;
  else
    Fnhg07 <= Rdc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bphg07 <= 1'b0;
  else
    Bphg07 <= Ydc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xqhg07 <= 1'b0;
  else
    Xqhg07 <= Fec8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tshg07 <= 1'b0;
  else
    Tshg07 <= Tec8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Puhg07 <= 1'b0;
  else
    Puhg07 <= Afc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mwhg07 <= 1'b0;
  else
    Mwhg07 <= Hfc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jyhg07 <= 1'b0;
  else
    Jyhg07 <= Ofc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    G0ig07 <= 1'b0;
  else
    G0ig07 <= Vfc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D2ig07 <= 1'b0;
  else
    D2ig07 <= Cgc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    A4ig07 <= 1'b0;
  else
    A4ig07 <= Jgc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X5ig07 <= 1'b0;
  else
    X5ig07 <= Xgc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U7ig07 <= 1'b0;
  else
    U7ig07 <= Ehc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R9ig07 <= 1'b0;
  else
    R9ig07 <= Lhc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Obig07 <= 1'b0;
  else
    Obig07 <= Shc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ldig07 <= 1'b0;
  else
    Ldig07 <= Zhc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ifig07 <= 1'b0;
  else
    Ifig07 <= Gic8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fhig07 <= 1'b0;
  else
    Fhig07 <= Uic8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cjig07 <= 1'b0;
  else
    Cjig07 <= Bjc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zkig07 <= 1'b0;
  else
    Zkig07 <= Ijc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wmig07 <= 1'b0;
  else
    Wmig07 <= Pjc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Toig07 <= 1'b0;
  else
    Toig07 <= Wjc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qqig07 <= 1'b0;
  else
    Qqig07 <= Dkc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nsig07 <= 1'b0;
  else
    Nsig07 <= Kkc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kuig07 <= 1'b0;
  else
    Kuig07 <= Rkc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hwig07 <= 1'b0;
  else
    Hwig07 <= Y5d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Myig07 <= 1'b0;
  else
    Myig07 <= Uad8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R0jg07 <= 1'b0;
  else
    R0jg07 <= Qfd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W2jg07 <= 1'b0;
  else
    W2jg07 <= Wpd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B5jg07 <= 1'b0;
  else
    B5jg07 <= Sud8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    G7jg07 <= 1'b0;
  else
    G7jg07 <= Ozd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L9jg07 <= 1'b0;
  else
    L9jg07 <= G9e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qbjg07 <= 1'b0;
  else
    Qbjg07 <= Cee8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vdjg07 <= 1'b0;
  else
    Vdjg07 <= R3f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Agjg07 <= 1'b0;
  else
    Agjg07 <= N8f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fijg07 <= 1'b0;
  else
    Fijg07 <= Qdf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kkjg07 <= 1'b0;
  else
    Kkjg07 <= U3d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Omjg07 <= 1'b0;
  else
    Omjg07 <= Q8d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sojg07 <= 1'b0;
  else
    Sojg07 <= Mdd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wqjg07 <= 1'b0;
  else
    Wqjg07 <= Snd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Atjg07 <= 1'b0;
  else
    Atjg07 <= Osd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Evjg07 <= 1'b0;
  else
    Evjg07 <= Kxd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ixjg07 <= 1'b0;
  else
    Ixjg07 <= C7e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mzjg07 <= 1'b0;
  else
    Mzjg07 <= Ybe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q1kg07 <= 1'b0;
  else
    Q1kg07 <= N1f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U3kg07 <= 1'b0;
  else
    U3kg07 <= J6f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y5kg07 <= 1'b0;
  else
    Y5kg07 <= Uff8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    C8kg07 <= 1'b0;
  else
    C8kg07 <= Muw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cakg07 <= 1'b0;
  else
    Cakg07 <= W4d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hckg07 <= 1'b0;
  else
    Hckg07 <= S9d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mekg07 <= 1'b0;
  else
    Mekg07 <= Oed8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rgkg07 <= 1'b0;
  else
    Rgkg07 <= Uod8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wikg07 <= 1'b0;
  else
    Wikg07 <= Qtd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Blkg07 <= 1'b0;
  else
    Blkg07 <= Myd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gnkg07 <= 1'b0;
  else
    Gnkg07 <= E8e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lpkg07 <= 1'b0;
  else
    Lpkg07 <= Ade8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qrkg07 <= 1'b0;
  else
    Qrkg07 <= P2f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vtkg07 <= 1'b0;
  else
    Vtkg07 <= L7f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Awkg07 <= 1'b0;
  else
    Awkg07 <= Sef8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fykg07 <= 1'b0;
  else
    Fykg07 <= S2d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J0lg07 <= 1'b0;
  else
    J0lg07 <= O7d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N2lg07 <= 1'b0;
  else
    N2lg07 <= Kcd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R4lg07 <= 1'b0;
  else
    R4lg07 <= Qmd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V6lg07 <= 1'b0;
  else
    V6lg07 <= Mrd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z8lg07 <= 1'b0;
  else
    Z8lg07 <= Iwd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dblg07 <= 1'b0;
  else
    Dblg07 <= A6e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hdlg07 <= 1'b0;
  else
    Hdlg07 <= Wae8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lflg07 <= 1'b0;
  else
    Lflg07 <= L0f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Phlg07 <= 1'b0;
  else
    Phlg07 <= H5f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tjlg07 <= 1'b0;
  else
    Tjlg07 <= Wgf8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xllg07 <= 1'b0;
  else
    Xllg07 <= Yql7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bolg07 <= 1'b0;
  else
    Bolg07 <= Rql7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qplg07 <= 1'b0;
  else
    Qplg07 <= Kql7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hrlg07 <= 1'b0;
  else
    Hrlg07 <= Dql7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yslg07 <= 1'b0;
  else
    Yslg07 <= Vc88v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zulg07 <= 1'b0;
  else
    Zulg07 <= Jd88v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Axlg07 <= 1'b0;
  else
    Axlg07 <= Ac88v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ezlg07 <= 1'b0;
  else
    Ezlg07 <= Hc88v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    I1mg07 <= 1'b0;
  else
    I1mg07 <= Oc88v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    H3mg07 <= 1'b0;
  else
    H3mg07 <= Cd88v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    I5mg07 <= 1'b0;
  else
    I5mg07 <= Qd88v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    J7mg07 <= 1'b0;
  else
    J7mg07 <= Zdo7v6;

always @(posedge FCLK) F9mg07 <= Hx88v6;
always @(posedge FCLK) Lbmg07 <= Ax88v6;
always @(posedge FCLK) Rdmg07 <= Tw88v6;
always @(posedge FCLK) Xfmg07 <= Mw88v6;
always @(posedge FCLK) Dimg07 <= Fw88v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hkmg07 <= 1'b0;
  else
    Hkmg07 <= Wpl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ylmg07 <= 1'b0;
  else
    Ylmg07 <= Rwe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pnmg07 <= 1'b0;
  else
    Pnmg07 <= Kwe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Epmg07 <= 1'b0;
  else
    Epmg07 <= Dwe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vqmg07 <= 1'b0;
  else
    Vqmg07 <= Wve8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Msmg07 <= 1'b0;
  else
    Msmg07 <= Pve8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dumg07 <= 1'b0;
  else
    Dumg07 <= Uue8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vvmg07 <= 1'b0;
  else
    Vvmg07 <= Nue8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nxmg07 <= 1'b0;
  else
    Nxmg07 <= Gue8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fzmg07 <= 1'b0;
  else
    Fzmg07 <= Zte8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X0ng07 <= 1'b0;
  else
    X0ng07 <= Ste8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P2ng07 <= 1'b0;
  else
    P2ng07 <= Lte8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H4ng07 <= 1'b0;
  else
    H4ng07 <= Ete8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z5ng07 <= 1'b0;
  else
    Z5ng07 <= Xse8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R7ng07 <= 1'b0;
  else
    R7ng07 <= Qse8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J9ng07 <= 1'b0;
  else
    J9ng07 <= Jse8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bbng07 <= 1'b0;
  else
    Bbng07 <= Cse8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tcng07 <= 1'b0;
  else
    Tcng07 <= Vre8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Leng07 <= 1'b0;
  else
    Leng07 <= Ore8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dgng07 <= 1'b0;
  else
    Dgng07 <= Hre8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vhng07 <= 1'b0;
  else
    Vhng07 <= Are8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Njng07 <= 1'b0;
  else
    Njng07 <= Tqe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Flng07 <= 1'b0;
  else
    Flng07 <= Mqe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xmng07 <= 1'b0;
  else
    Xmng07 <= Fqe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pong07 <= 1'b0;
  else
    Pong07 <= Ype8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hqng07 <= 1'b0;
  else
    Hqng07 <= Rpe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zrng07 <= 1'b0;
  else
    Zrng07 <= Kpe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rtng07 <= 1'b0;
  else
    Rtng07 <= Dpe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jvng07 <= 1'b0;
  else
    Jvng07 <= Woe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Axng07 <= 1'b0;
  else
    Axng07 <= Poe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ryng07 <= 1'b0;
  else
    Ryng07 <= Ioe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    I0og07 <= 1'b0;
  else
    I0og07 <= Boe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z1og07 <= 1'b0;
  else
    Z1og07 <= Une8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q3og07 <= 1'b0;
  else
    Q3og07 <= Nne8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H5og07 <= 1'b0;
  else
    H5og07 <= Gne8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y6og07 <= 1'b0;
  else
    Y6og07 <= Zme8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P8og07 <= 1'b0;
  else
    P8og07 <= Sme8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gaog07 <= 1'b0;
  else
    Gaog07 <= Yv88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ncog07 <= 1'b0;
  else
    Ncog07 <= Qqo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Eeog07 <= 1'b0;
  else
    Eeog07 <= Jqo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vfog07 <= 1'b0;
  else
    Vfog07 <= Cqo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mhog07 <= 1'b0;
  else
    Mhog07 <= Vpo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Djog07 <= 1'b0;
  else
    Djog07 <= Opo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ukog07 <= 1'b0;
  else
    Ukog07 <= Hpo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lmog07 <= 1'b0;
  else
    Lmog07 <= Apo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Coog07 <= 1'b0;
  else
    Coog07 <= Too7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tpog07 <= 1'b0;
  else
    Tpog07 <= Moo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Krog07 <= 1'b0;
  else
    Krog07 <= Foo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Btog07 <= 1'b0;
  else
    Btog07 <= Yno7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tuog07 <= 1'b0;
  else
    Tuog07 <= Rno7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lwog07 <= 1'b0;
  else
    Lwog07 <= Kno7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dyog07 <= 1'b0;
  else
    Dyog07 <= Dno7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vzog07 <= 1'b0;
  else
    Vzog07 <= Wmo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N1pg07 <= 1'b0;
  else
    N1pg07 <= Pmo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F3pg07 <= 1'b0;
  else
    F3pg07 <= Imo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X4pg07 <= 1'b0;
  else
    X4pg07 <= Bmo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P6pg07 <= 1'b0;
  else
    P6pg07 <= Ulo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H8pg07 <= 1'b0;
  else
    H8pg07 <= Nlo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z9pg07 <= 1'b0;
  else
    Z9pg07 <= Glo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rbpg07 <= 1'b0;
  else
    Rbpg07 <= Zko7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jdpg07 <= 1'b0;
  else
    Jdpg07 <= Sko7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bfpg07 <= 1'b0;
  else
    Bfpg07 <= Lko7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tgpg07 <= 1'b0;
  else
    Tgpg07 <= Eko7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lipg07 <= 1'b0;
  else
    Lipg07 <= Xjo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dkpg07 <= 1'b0;
  else
    Dkpg07 <= Qjo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vlpg07 <= 1'b0;
  else
    Vlpg07 <= Jjo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nnpg07 <= 1'b0;
  else
    Nnpg07 <= Vio7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fppg07 <= 1'b0;
  else
    Fppg07 <= Oio7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xqpg07 <= 1'b0;
  else
    Xqpg07 <= Hio7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pspg07 <= 1'b0;
  else
    Pspg07 <= Ppl7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Supg07 <= 1'b0;
  else
    Supg07 <= Ipl7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xwpg07 <= 1'b0;
  else
    Xwpg07 <= Bpl7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Azpg07 <= 1'b0;
  else
    Azpg07 <= Uol7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    C1qg07 <= 1'b0;
  else
    C1qg07 <= Nol7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    G3qg07 <= 1'b0;
  else
    G3qg07 <= Gol7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    J5qg07 <= 1'b0;
  else
    J5qg07 <= Znl7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    N7qg07 <= 1'b0;
  else
    N7qg07 <= Snl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T9qg07 <= 1'b0;
  else
    T9qg07 <= Lnl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ubqg07 <= 1'b0;
  else
    Ubqg07 <= Enl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wdqg07 <= 1'b0;
  else
    Wdqg07 <= En68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yfqg07 <= 1'b0;
  else
    Yfqg07 <= Qt68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Biqg07 <= 1'b0;
  else
    Biqg07 <= Ct68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dkqg07 <= 1'b0;
  else
    Dkqg07 <= Vs68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gmqg07 <= 1'b0;
  else
    Gmqg07 <= Os68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Joqg07 <= 1'b0;
  else
    Joqg07 <= Hs68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mqqg07 <= 1'b0;
  else
    Mqqg07 <= As68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Psqg07 <= 1'b0;
  else
    Psqg07 <= Tr68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Suqg07 <= 1'b0;
  else
    Suqg07 <= Yq68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vwqg07 <= 1'b0;
  else
    Vwqg07 <= Dq68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yyqg07 <= 1'b0;
  else
    Yyqg07 <= Wp68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B1rg07 <= 1'b0;
  else
    B1rg07 <= Ip68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    E3rg07 <= 1'b0;
  else
    E3rg07 <= Uo68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H5rg07 <= 1'b0;
  else
    H5rg07 <= No68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K7rg07 <= 1'b0;
  else
    K7rg07 <= Go68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N9rg07 <= 1'b0;
  else
    N9rg07 <= Zn68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qbrg07 <= 1'b0;
  else
    Qbrg07 <= Sn68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tdrg07 <= 1'b0;
  else
    Tdrg07 <= Ln68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wfrg07 <= 1'b0;
  else
    Wfrg07 <= Xml7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yhrg07 <= 1'b0;
  else
    Yhrg07 <= Qml7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Akrg07 <= 1'b0;
  else
    Akrg07 <= Jml7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cmrg07 <= 1'b0;
  else
    Cmrg07 <= Cml7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Eorg07 <= 1'b0;
  else
    Eorg07 <= Vll7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gqrg07 <= 1'b0;
  else
    Gqrg07 <= Oll7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Isrg07 <= 1'b0;
  else
    Isrg07 <= Hll7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kurg07 <= 1'b0;
  else
    Kurg07 <= All7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mwrg07 <= 1'b0;
  else
    Mwrg07 <= Tkl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oyrg07 <= 1'b0;
  else
    Oyrg07 <= R5d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T0sg07 <= 1'b0;
  else
    T0sg07 <= Nad8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y2sg07 <= 1'b0;
  else
    Y2sg07 <= Jfd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D5sg07 <= 1'b0;
  else
    D5sg07 <= Ppd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    I7sg07 <= 1'b0;
  else
    I7sg07 <= Lud8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N9sg07 <= 1'b0;
  else
    N9sg07 <= Hzd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sbsg07 <= 1'b0;
  else
    Sbsg07 <= Z8e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xdsg07 <= 1'b0;
  else
    Xdsg07 <= Vde8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cgsg07 <= 1'b0;
  else
    Cgsg07 <= K3f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hisg07 <= 1'b0;
  else
    Hisg07 <= G8f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mksg07 <= 1'b0;
  else
    Mksg07 <= Xdf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rmsg07 <= 1'b0;
  else
    Rmsg07 <= N3d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vosg07 <= 1'b0;
  else
    Vosg07 <= J8d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zqsg07 <= 1'b0;
  else
    Zqsg07 <= Fdd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dtsg07 <= 1'b0;
  else
    Dtsg07 <= Lnd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hvsg07 <= 1'b0;
  else
    Hvsg07 <= Hsd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lxsg07 <= 1'b0;
  else
    Lxsg07 <= Dxd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pzsg07 <= 1'b0;
  else
    Pzsg07 <= V6e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T1tg07 <= 1'b0;
  else
    T1tg07 <= Rbe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X3tg07 <= 1'b0;
  else
    X3tg07 <= G1f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B6tg07 <= 1'b0;
  else
    B6tg07 <= C6f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F8tg07 <= 1'b0;
  else
    F8tg07 <= Bgf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jatg07 <= 1'b0;
  else
    Jatg07 <= Mkl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kctg07 <= 1'b0;
  else
    Kctg07 <= Fkl7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Letg07 <= 1'b0;
  else
    Letg07 <= A8y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kgtg07 <= 1'b0;
  else
    Kgtg07 <= O8y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jitg07 <= 1'b0;
  else
    Jitg07 <= V8y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Iktg07 <= 1'b0;
  else
    Iktg07 <= C9y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hmtg07 <= 1'b0;
  else
    Hmtg07 <= J9y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hotg07 <= 1'b0;
  else
    Hotg07 <= Q9y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hqtg07 <= 1'b0;
  else
    Hqtg07 <= Eay7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hstg07 <= 1'b0;
  else
    Hstg07 <= Lay7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hutg07 <= 1'b0;
  else
    Hutg07 <= Say7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hwtg07 <= 1'b0;
  else
    Hwtg07 <= Gby7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hytg07 <= 1'b0;
  else
    Hytg07 <= Wyx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    G0ug07 <= 1'b0;
  else
    G0ug07 <= Dzx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F2ug07 <= 1'b0;
  else
    F2ug07 <= Nby7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    E4ug07 <= 1'b0;
  else
    E4ug07 <= P4d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J6ug07 <= 1'b0;
  else
    J6ug07 <= L9d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O8ug07 <= 1'b0;
  else
    O8ug07 <= Hed8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Taug07 <= 1'b0;
  else
    Taug07 <= Nod8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ycug07 <= 1'b0;
  else
    Ycug07 <= Jtd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dfug07 <= 1'b0;
  else
    Dfug07 <= Fyd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ihug07 <= 1'b0;
  else
    Ihug07 <= X7e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Njug07 <= 1'b0;
  else
    Njug07 <= Tce8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Slug07 <= 1'b0;
  else
    Slug07 <= I2f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xnug07 <= 1'b0;
  else
    Xnug07 <= E7f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cqug07 <= 1'b0;
  else
    Cqug07 <= Zef8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hsug07 <= 1'b0;
  else
    Hsug07 <= Dhf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Luug07 <= 1'b0;
  else
    Luug07 <= A5f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pwug07 <= 1'b0;
  else
    Pwug07 <= E0f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tyug07 <= 1'b0;
  else
    Tyug07 <= Pae8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X0vg07 <= 1'b0;
  else
    X0vg07 <= T5e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B3vg07 <= 1'b0;
  else
    B3vg07 <= Bwd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F5vg07 <= 1'b0;
  else
    F5vg07 <= Frd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J7vg07 <= 1'b0;
  else
    J7vg07 <= Jmd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N9vg07 <= 1'b0;
  else
    N9vg07 <= Dcd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rbvg07 <= 1'b0;
  else
    Rbvg07 <= H7d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vdvg07 <= 1'b0;
  else
    Vdvg07 <= L2d8v6;

always @(posedge HCLK) Zfvg07 <= Z1e8v6;
always @(posedge HCLK) Aivg07 <= S1e8v6;
always @(posedge HCLK) Bkvg07 <= L1e8v6;
always @(posedge HCLK) Cmvg07 <= E1e8v6;
always @(posedge HCLK) Dovg07 <= X0e8v6;
always @(posedge HCLK) Eqvg07 <= Q0e8v6;
always @(posedge HCLK) Fsvg07 <= Qle8v6;
always @(posedge HCLK) Guvg07 <= Jle8v6;
always @(posedge HCLK) Hwvg07 <= Cle8v6;
always @(posedge HCLK) Iyvg07 <= Vke8v6;
always @(posedge HCLK) J0wg07 <= Oke8v6;
always @(posedge HCLK) K2wg07 <= Hke8v6;
always @(posedge HCLK) L4wg07 <= Ake8v6;
always @(posedge HCLK) M6wg07 <= Tje8v6;
always @(posedge HCLK) N8wg07 <= Bid8v6;
always @(posedge HCLK) Nawg07 <= Uhd8v6;
always @(posedge HCLK) Ocwg07 <= Nhd8v6;
always @(posedge HCLK) Pewg07 <= Ghd8v6;
always @(posedge HCLK) Qgwg07 <= Zgd8v6;
always @(posedge HCLK) Riwg07 <= Sgd8v6;
always @(posedge HCLK) Skwg07 <= Lgd8v6;
always @(posedge HCLK) Tmwg07 <= Eac8v6;
always @(posedge HCLK) Towg07 <= Lac8v6;
always @(posedge HCLK) Tqwg07 <= Sac8v6;
always @(posedge HCLK) Tswg07 <= Zac8v6;
always @(posedge HCLK) Tuwg07 <= Gbc8v6;
always @(posedge HCLK) Twwg07 <= Ubc8v6;
always @(posedge HCLK) Tywg07 <= Bcc8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T0xg07 <= 1'b1;
  else
    T0xg07 <= Djd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U2xg07 <= 1'b0;
  else
    U2xg07 <= H948v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    S5xg07 <= 1'b0;
  else
    S5xg07 <= A948v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q8xg07 <= 1'b0;
  else
    Q8xg07 <= K5d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vaxg07 <= 1'b0;
  else
    Vaxg07 <= Gad8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Adxg07 <= 1'b0;
  else
    Adxg07 <= Cfd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ffxg07 <= 1'b0;
  else
    Ffxg07 <= Ipd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Khxg07 <= 1'b0;
  else
    Khxg07 <= Eud8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pjxg07 <= 1'b0;
  else
    Pjxg07 <= Azd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ulxg07 <= 1'b0;
  else
    Ulxg07 <= S8e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Znxg07 <= 1'b0;
  else
    Znxg07 <= Ode8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Eqxg07 <= 1'b0;
  else
    Eqxg07 <= D3f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jsxg07 <= 1'b0;
  else
    Jsxg07 <= Z7f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ouxg07 <= 1'b0;
  else
    Ouxg07 <= Eef8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Twxg07 <= 1'b0;
  else
    Twxg07 <= Igf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xyxg07 <= 1'b0;
  else
    Xyxg07 <= V5f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B1yg07 <= 1'b0;
  else
    B1yg07 <= Z0f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F3yg07 <= 1'b0;
  else
    F3yg07 <= Kbe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J5yg07 <= 1'b0;
  else
    J5yg07 <= O6e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N7yg07 <= 1'b0;
  else
    N7yg07 <= Wwd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R9yg07 <= 1'b0;
  else
    R9yg07 <= Asd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vbyg07 <= 1'b0;
  else
    Vbyg07 <= End8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zdyg07 <= 1'b0;
  else
    Zdyg07 <= Ycd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dgyg07 <= 1'b0;
  else
    Dgyg07 <= C8d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hiyg07 <= 1'b0;
  else
    Hiyg07 <= G3d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lkyg07 <= 1'b0;
  else
    Lkyg07 <= Yh88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nmyg07 <= 1'b0;
  else
    Nmyg07 <= Wxc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Poyg07 <= 1'b0;
  else
    Poyg07 <= Mzc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rqyg07 <= 1'b0;
  else
    Rqyg07 <= H0d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tsyg07 <= 1'b0;
  else
    Tsyg07 <= Q1d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vuyg07 <= 1'b0;
  else
    Vuyg07 <= M6d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xwyg07 <= 1'b0;
  else
    Xwyg07 <= Ibd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zyyg07 <= 1'b0;
  else
    Zyyg07 <= Wid8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B1zg07 <= 1'b0;
  else
    B1zg07 <= Rjd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    E3zg07 <= 1'b0;
  else
    E3zg07 <= Mkd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H5zg07 <= 1'b0;
  else
    H5zg07 <= Ald8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K7zg07 <= 1'b0;
  else
    K7zg07 <= Old8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N9zg07 <= 1'b0;
  else
    N9zg07 <= Kqd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qbzg07 <= 1'b0;
  else
    Qbzg07 <= Gvd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tdzg07 <= 1'b0;
  else
    Tdzg07 <= U2e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wfzg07 <= 1'b0;
  else
    Wfzg07 <= I3e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zhzg07 <= 1'b0;
  else
    Zhzg07 <= W3e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ckzg07 <= 1'b0;
  else
    Ckzg07 <= K4e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fmzg07 <= 1'b0;
  else
    Fmzg07 <= Y4e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Iozg07 <= 1'b0;
  else
    Iozg07 <= U9e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lqzg07 <= 1'b0;
  else
    Lqzg07 <= Mje8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oszg07 <= 1'b0;
  else
    Oszg07 <= Fxe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ruzg07 <= 1'b0;
  else
    Ruzg07 <= Txe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uwzg07 <= 1'b0;
  else
    Uwzg07 <= Hye8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xyzg07 <= 1'b0;
  else
    Xyzg07 <= Vye8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    A10h07 <= 1'b0;
  else
    A10h07 <= Jze8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D30h07 <= 1'b0;
  else
    D30h07 <= F4f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    G50h07 <= 1'b0;
  else
    G50h07 <= Cdf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J70h07 <= 1'b0;
  else
    J70h07 <= Kzx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L90h07 <= 1'b0;
  else
    L90h07 <= Yzx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nb0h07 <= 1'b0;
  else
    Nb0h07 <= H1y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pd0h07 <= 1'b0;
  else
    Pd0h07 <= C2y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rf0h07 <= 1'b0;
  else
    Rf0h07 <= J2y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Th0h07 <= 1'b0;
  else
    Th0h07 <= Q2y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vj0h07 <= 1'b0;
  else
    Vj0h07 <= X2y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xl0h07 <= 1'b0;
  else
    Xl0h07 <= S3y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zn0h07 <= 1'b0;
  else
    Zn0h07 <= G4y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bq0h07 <= 1'b0;
  else
    Bq0h07 <= N4y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ds0h07 <= 1'b0;
  else
    Ds0h07 <= U4y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fu0h07 <= 1'b0;
  else
    Fu0h07 <= P5y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hw0h07 <= 1'b0;
  else
    Hw0h07 <= W5y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Iy0h07 <= 1'b0;
  else
    Iy0h07 <= D6y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J01h07 <= 1'b0;
  else
    J01h07 <= K6y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K21h07 <= 1'b0;
  else
    K21h07 <= R6y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L41h07 <= 1'b0;
  else
    L41h07 <= Y6y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M61h07 <= 1'b0;
  else
    M61h07 <= M7y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N81h07 <= 1'b0;
  else
    N81h07 <= T7y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oa1h07 <= 1'b0;
  else
    Oa1h07 <= Daf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hd1h07 <= 1'b0;
  else
    Hd1h07 <= Yaf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ag1h07 <= 1'b0;
  else
    Ag1h07 <= Mbf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ni1h07 <= 1'b0;
  else
    Ni1h07 <= X8k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ml1h07 <= 1'b0;
  else
    Ml1h07 <= Tbf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lo1h07 <= 1'b0;
  else
    Lo1h07 <= Fbf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zq1h07 <= 1'b0;
  else
    Zq1h07 <= Raf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    St1h07 <= 1'b0;
  else
    St1h07 <= Kaf8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lw1h07 <= 1'b0;
  else
    Lw1h07 <= W9f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kz1h07 <= 1'b0;
  else
    Kz1h07 <= P9f8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J22h07 <= 1'b0;
  else
    J22h07 <= Zvc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F52h07 <= 1'b0;
  else
    F52h07 <= Dyc8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    C82h07 <= 1'b0;
  else
    C82h07 <= Xd88v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    R92h07 <= 1'b0;
  else
    R92h07 <= Wq58v6;

always @(posedge HCLK) Fb2h07 <= Kr58v6;
always @(posedge HCLK) Xc2h07 <= Cu58v6;
always @(posedge HCLK) Ne2h07 <= Xu58v6;
always @(posedge HCLK) Dg2h07 <= Gw58v6;
always @(posedge HCLK) Th2h07 <= Nw58v6;
always @(posedge HCLK) Ij2h07 <= Uw58v6;
always @(posedge HCLK) Xk2h07 <= Px58v6;
always @(posedge HCLK) Mm2h07 <= Wx58v6;
always @(posedge HCLK) Bo2h07 <= Ry58v6;
always @(posedge HCLK) Qp2h07 <= Bx58v6;
always @(posedge HCLK) Fr2h07 <= Zv58v6;
always @(posedge HCLK) Vs2h07 <= Sv58v6;
always @(posedge HCLK) Lu2h07 <= Lv58v6;
always @(posedge HCLK) Bw2h07 <= Vt58v6;
always @(posedge HCLK) Rx2h07 <= Ts58v6;
always @(posedge HCLK) Hz2h07 <= Ms58v6;
always @(posedge HCLK) X03h07 <= Fs58v6;
always @(posedge HCLK) N23h07 <= Yr58v6;
always @(posedge HCLK) D43h07 <= Rr58v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    V53h07 <= 1'b0;
  else
    V53h07 <= A768v6;

always @(posedge HCLK) J73h07 <= O768v6;
always @(posedge HCLK) B93h07 <= Ga68v6;
always @(posedge HCLK) Ra3h07 <= Bb68v6;
always @(posedge HCLK) Hc3h07 <= Kc68v6;
always @(posedge HCLK) Xd3h07 <= Rc68v6;
always @(posedge HCLK) Mf3h07 <= Yc68v6;
always @(posedge HCLK) Bh3h07 <= Td68v6;
always @(posedge HCLK) Qi3h07 <= Ae68v6;
always @(posedge HCLK) Fk3h07 <= Ve68v6;
always @(posedge HCLK) Ul3h07 <= Fd68v6;
always @(posedge HCLK) Jn3h07 <= Dc68v6;
always @(posedge HCLK) Zo3h07 <= Wb68v6;
always @(posedge HCLK) Pq3h07 <= Pb68v6;
always @(posedge HCLK) Fs3h07 <= Z968v6;
always @(posedge HCLK) Vt3h07 <= X868v6;
always @(posedge HCLK) Lv3h07 <= Q868v6;
always @(posedge HCLK) Bx3h07 <= J868v6;
always @(posedge HCLK) Ry3h07 <= C868v6;
always @(posedge HCLK) H04h07 <= V768v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Z14h07 <= 1'b0;
  else
    Z14h07 <= Ol68v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    M34h07 <= 1'b0;
  else
    M34h07 <= Cv48v6;

always @(posedge HCLK) A54h07 <= Ux48v6;
always @(posedge HCLK) Q64h07 <= Py48v6;
always @(posedge HCLK) G84h07 <= Yz48v6;
always @(posedge HCLK) W94h07 <= F058v6;
always @(posedge HCLK) Lb4h07 <= M058v6;
always @(posedge HCLK) Ad4h07 <= H158v6;
always @(posedge HCLK) Pe4h07 <= O158v6;
always @(posedge HCLK) Eg4h07 <= J258v6;
always @(posedge HCLK) Th4h07 <= T058v6;
always @(posedge HCLK) Ij4h07 <= Rz48v6;
always @(posedge HCLK) Yk4h07 <= Kz48v6;
always @(posedge HCLK) Om4h07 <= Dz48v6;
always @(posedge HCLK) Eo4h07 <= Nx48v6;
always @(posedge HCLK) Up4h07 <= Lw48v6;
always @(posedge HCLK) Kr4h07 <= Ew48v6;
always @(posedge HCLK) At4h07 <= Xv48v6;
always @(posedge HCLK) Qu4h07 <= Qv48v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gw4h07 <= 1'b0;
  else
    Gw4h07 <= On48v6;

always @(posedge HCLK) Ux4h07 <= Gq48v6;
always @(posedge HCLK) Kz4h07 <= Br48v6;
always @(posedge HCLK) A15h07 <= Rs48v6;
always @(posedge HCLK) P25h07 <= Ys48v6;
always @(posedge HCLK) E45h07 <= Tt48v6;
always @(posedge HCLK) T55h07 <= Au48v6;
always @(posedge HCLK) I75h07 <= Vu48v6;
always @(posedge HCLK) X85h07 <= Ft48v6;
always @(posedge HCLK) Ma5h07 <= Ds48v6;
always @(posedge HCLK) Cc5h07 <= Wr48v6;
always @(posedge HCLK) Sd5h07 <= Pr48v6;
always @(posedge HCLK) If5h07 <= Xo48v6;
always @(posedge HCLK) Yg5h07 <= Qo48v6;
always @(posedge HCLK) Oi5h07 <= Jo48v6;
always @(posedge HCLK) Ek5h07 <= Co48v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ul5h07 <= 1'b0;
  else
    Ul5h07 <= Yy58v6;

always @(posedge HCLK) In5h07 <= Mz58v6;
always @(posedge HCLK) Ap5h07 <= E268v6;
always @(posedge HCLK) Qq5h07 <= Z268v6;
always @(posedge HCLK) Gs5h07 <= I468v6;
always @(posedge HCLK) Wt5h07 <= P468v6;
always @(posedge HCLK) Lv5h07 <= W468v6;
always @(posedge HCLK) Ax5h07 <= R568v6;
always @(posedge HCLK) Py5h07 <= Y568v6;
always @(posedge HCLK) E06h07 <= T668v6;
always @(posedge HCLK) T16h07 <= D568v6;
always @(posedge HCLK) I36h07 <= B468v6;
always @(posedge HCLK) Y46h07 <= U368v6;
always @(posedge HCLK) O66h07 <= N368v6;
always @(posedge HCLK) E86h07 <= X168v6;
always @(posedge HCLK) U96h07 <= V068v6;
always @(posedge HCLK) Kb6h07 <= O068v6;
always @(posedge HCLK) Ad6h07 <= H068v6;
always @(posedge HCLK) Qe6h07 <= A068v6;
always @(posedge HCLK) Gg6h07 <= Tz58v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yh6h07 <= 1'b0;
  else
    Yh6h07 <= Sa58v6;

always @(posedge HCLK) Mj6h07 <= Gb58v6;
always @(posedge HCLK) El6h07 <= Yd58v6;
always @(posedge HCLK) Um6h07 <= Te58v6;
always @(posedge HCLK) Ko6h07 <= Cg58v6;
always @(posedge HCLK) Aq6h07 <= Jg58v6;
always @(posedge HCLK) Pr6h07 <= Qg58v6;
always @(posedge HCLK) Et6h07 <= Lh58v6;
always @(posedge HCLK) Tu6h07 <= Sh58v6;
always @(posedge HCLK) Iw6h07 <= Ni58v6;
always @(posedge HCLK) Xx6h07 <= Xg58v6;
always @(posedge HCLK) Mz6h07 <= Vf58v6;
always @(posedge HCLK) C17h07 <= Of58v6;
always @(posedge HCLK) S27h07 <= Hf58v6;
always @(posedge HCLK) I47h07 <= Rd58v6;
always @(posedge HCLK) Y57h07 <= Pc58v6;
always @(posedge HCLK) O77h07 <= Ic58v6;
always @(posedge HCLK) E97h07 <= Bc58v6;
always @(posedge HCLK) Ua7h07 <= Ub58v6;
always @(posedge HCLK) Kc7h07 <= Nb58v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ce7h07 <= 1'b0;
  else
    Ce7h07 <= Q258v6;

always @(posedge HCLK) Qf7h07 <= W558v6;
always @(posedge HCLK) Gh7h07 <= R658v6;
always @(posedge HCLK) Wi7h07 <= A858v6;
always @(posedge HCLK) Mk7h07 <= H858v6;
always @(posedge HCLK) Bm7h07 <= O858v6;
always @(posedge HCLK) Qn7h07 <= J958v6;
always @(posedge HCLK) Fp7h07 <= Q958v6;
always @(posedge HCLK) Uq7h07 <= La58v6;
always @(posedge HCLK) Js7h07 <= V858v6;
always @(posedge HCLK) Yt7h07 <= T758v6;
always @(posedge HCLK) Ov7h07 <= M758v6;
always @(posedge HCLK) Ex7h07 <= F758v6;
always @(posedge HCLK) Uy7h07 <= P558v6;
always @(posedge HCLK) K08h07 <= N458v6;
always @(posedge HCLK) A28h07 <= G458v6;
always @(posedge HCLK) Q38h07 <= Z358v6;
always @(posedge HCLK) G58h07 <= S358v6;
always @(posedge HCLK) W68h07 <= L358v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    O88h07 <= 1'b0;
  else
    O88h07 <= Ui58v6;

always @(posedge HCLK) Ca8h07 <= Ij58v6;
always @(posedge HCLK) Ub8h07 <= Am58v6;
always @(posedge HCLK) Kd8h07 <= Vm58v6;
always @(posedge HCLK) Af8h07 <= Eo58v6;
always @(posedge HCLK) Qg8h07 <= Lo58v6;
always @(posedge HCLK) Fi8h07 <= So58v6;
always @(posedge HCLK) Uj8h07 <= Np58v6;
always @(posedge HCLK) Jl8h07 <= Up58v6;
always @(posedge HCLK) Ym8h07 <= Pq58v6;
always @(posedge HCLK) No8h07 <= Zo58v6;
always @(posedge HCLK) Cq8h07 <= Xn58v6;
always @(posedge HCLK) Sr8h07 <= Qn58v6;
always @(posedge HCLK) It8h07 <= Jn58v6;
always @(posedge HCLK) Yu8h07 <= Tl58v6;
always @(posedge HCLK) Ow8h07 <= Rk58v6;
always @(posedge HCLK) Ey8h07 <= Kk58v6;
always @(posedge HCLK) Uz8h07 <= Dk58v6;
always @(posedge HCLK) K19h07 <= Wj58v6;
always @(posedge HCLK) A39h07 <= Pj58v6;
always @(posedge HCLK) S49h07 <= Nh68v6;
always @(posedge HCLK) J69h07 <= Ii68v6;
always @(posedge HCLK) A89h07 <= Rj68v6;
always @(posedge HCLK) Q99h07 <= Yj68v6;
always @(posedge HCLK) Gb9h07 <= Fk68v6;
always @(posedge HCLK) Wc9h07 <= Al68v6;
always @(posedge HCLK) Me9h07 <= Hl68v6;
always @(posedge HCLK) Cg9h07 <= Mk68v6;
always @(posedge HCLK) Sh9h07 <= Kj68v6;
always @(posedge HCLK) Ij9h07 <= Dj68v6;
always @(posedge HCLK) Yk9h07 <= Wi68v6;
always @(posedge HCLK) Pm9h07 <= Gh68v6;
always @(posedge HCLK) Go9h07 <= Eg68v6;
always @(posedge HCLK) Xp9h07 <= Xf68v6;
always @(posedge HCLK) Or9h07 <= Qf68v6;
always @(posedge HCLK) Ft9h07 <= Jf68v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wu9h07 <= 1'b0;
  else
    Wu9h07 <= Tb88v6;

always @(posedge FCLK) Xw9h07 <= Yjl7v6;
always @(posedge FCLK) Zy9h07 <= Rjl7v6;
always @(posedge FCLK) B1ah07 <= Kjl7v6;
always @(posedge FCLK) D3ah07 <= Qjv7v6;
always @(posedge FCLK) J5ah07 <= Ekv7v6;
always @(posedge FCLK) P7ah07 <= Djl7v6;
always @(posedge FCLK) R9ah07 <= Wil7v6;
always @(posedge FCLK) Tbah07 <= Pil7v6;
always @(posedge FCLK) Vdah07 <= Mhv7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bgah07 <= 1'b0;
  else
    Bgah07 <= Iil7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hiah07 <= 1'b0;
  else
    Hiah07 <= Bil7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jkah07 <= 1'b0;
  else
    Jkah07 <= Uhl7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lmah07 <= 1'b0;
  else
    Lmah07 <= Nhl7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Noah07 <= 1'b0;
  else
    Noah07 <= Ghl7v6;

always @(posedge FCLK) Oqah07 <= Zgl7v6;
always @(posedge FCLK) Msah07 <= Sgl7v6;
always @(posedge FCLK) Luah07 <= Lgl7v6;
always @(posedge FCLK) Kwah07 <= Egl7v6;
always @(posedge FCLK) Jyah07 <= Xfl7v6;
always @(posedge FCLK) I0bh07 <= Qfl7v6;
always @(posedge FCLK) H2bh07 <= Jfl7v6;
always @(posedge FCLK) G4bh07 <= Cfl7v6;
always @(posedge FCLK) F6bh07 <= Vel7v6;
always @(posedge FCLK) E8bh07 <= Oel7v6;
always @(posedge FCLK) Dabh07 <= Hel7v6;
always @(posedge FCLK) Ccbh07 <= Ael7v6;
always @(posedge FCLK) Bebh07 <= Tdl7v6;
always @(posedge FCLK) Agbh07 <= Mdl7v6;
always @(posedge FCLK) Zhbh07 <= Fdl7v6;
always @(posedge FCLK) Yjbh07 <= Ycl7v6;
always @(posedge FCLK) Xlbh07 <= Rcl7v6;
always @(posedge FCLK) Wnbh07 <= Kcl7v6;
always @(posedge FCLK) Vpbh07 <= Dcl7v6;
always @(posedge FCLK) Urbh07 <= Wbl7v6;
always @(posedge FCLK) Ttbh07 <= Pbl7v6;
always @(posedge FCLK) Svbh07 <= Ibl7v6;
always @(posedge FCLK) Rxbh07 <= Bbl7v6;
always @(posedge FCLK) Qzbh07 <= Ual7v6;
always @(posedge FCLK) O1ch07 <= Nal7v6;
always @(posedge FCLK) M3ch07 <= Gal7v6;
always @(posedge FCLK) K5ch07 <= Z9l7v6;
always @(posedge FCLK) I7ch07 <= S9l7v6;
always @(posedge FCLK) G9ch07 <= L9l7v6;
always @(posedge FCLK) Ebch07 <= E9l7v6;
always @(posedge FCLK) Cdch07 <= X8l7v6;
always @(posedge FCLK) Afch07 <= Q8l7v6;
always @(posedge FCLK) Chch07 <= J8l7v6;
always @(posedge FCLK) Fjch07 <= C8l7v6;
always @(posedge FCLK) Ilch07 <= V7l7v6;
always @(posedge FCLK) Lnch07 <= O7l7v6;
always @(posedge FCLK) Opch07 <= H7l7v6;
always @(posedge FCLK) Rrch07 <= A7l7v6;
always @(posedge FCLK) Utch07 <= T6l7v6;
always @(posedge FCLK) Xvch07 <= M6l7v6;
always @(posedge FCLK) Aych07 <= F6l7v6;
always @(posedge FCLK) D0dh07 <= Y5l7v6;
always @(posedge FCLK) G2dh07 <= R5l7v6;
always @(posedge FCLK) J4dh07 <= K5l7v6;
always @(posedge FCLK) M6dh07 <= D5l7v6;
always @(posedge FCLK) P8dh07 <= W4l7v6;
always @(posedge FCLK) Sadh07 <= P4l7v6;
always @(posedge FCLK) Vcdh07 <= I4l7v6;
always @(posedge FCLK) Yedh07 <= B4l7v6;
always @(posedge FCLK) Bhdh07 <= U3l7v6;
always @(posedge FCLK) Ejdh07 <= N3l7v6;
always @(posedge FCLK) Hldh07 <= G3l7v6;
always @(posedge FCLK) Kndh07 <= Z2l7v6;
always @(posedge FCLK) Npdh07 <= S2l7v6;
always @(posedge FCLK) Qrdh07 <= L2l7v6;
always @(posedge FCLK) Stdh07 <= E2l7v6;
always @(posedge FCLK) Uvdh07 <= X1l7v6;
always @(posedge FCLK) Wxdh07 <= Q1l7v6;
always @(posedge FCLK) Yzdh07 <= J1l7v6;
always @(posedge FCLK) A2eh07 <= C1l7v6;
always @(posedge FCLK) C4eh07 <= V0l7v6;
always @(posedge FCLK) E6eh07 <= O0l7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    G8eh07 <= 1'b0;
  else
    G8eh07 <= H0l7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Daeh07 <= 1'b0;
  else
    Daeh07 <= A0l7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bceh07 <= 1'b0;
  else
    Bceh07 <= Tzk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zdeh07 <= 1'b0;
  else
    Zdeh07 <= Mzk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xfeh07 <= 1'b0;
  else
    Xfeh07 <= Fzk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vheh07 <= 1'b0;
  else
    Vheh07 <= Yyk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tjeh07 <= 1'b0;
  else
    Tjeh07 <= Ryk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rleh07 <= 1'b0;
  else
    Rleh07 <= Kyk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pneh07 <= 1'b0;
  else
    Pneh07 <= Dyk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Npeh07 <= 1'b0;
  else
    Npeh07 <= Wxk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lreh07 <= 1'b0;
  else
    Lreh07 <= Pxk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jteh07 <= 1'b0;
  else
    Jteh07 <= Ixk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hveh07 <= 1'b0;
  else
    Hveh07 <= Bxk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fxeh07 <= 1'b0;
  else
    Fxeh07 <= Uwk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dzeh07 <= 1'b0;
  else
    Dzeh07 <= Nwk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    A1fh07 <= 1'b0;
  else
    A1fh07 <= Gwk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    X2fh07 <= 1'b0;
  else
    X2fh07 <= Zvk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    U4fh07 <= 1'b0;
  else
    U4fh07 <= Svk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    R6fh07 <= 1'b0;
  else
    R6fh07 <= Lvk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    O8fh07 <= 1'b0;
  else
    O8fh07 <= Evk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lafh07 <= 1'b0;
  else
    Lafh07 <= Xuk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Icfh07 <= 1'b0;
  else
    Icfh07 <= Quk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fefh07 <= 1'b0;
  else
    Fefh07 <= Juk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kgfh07 <= 1'b0;
  else
    Kgfh07 <= Cuk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qifh07 <= 1'b0;
  else
    Qifh07 <= Vtk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wkfh07 <= 1'b0;
  else
    Wkfh07 <= Otk7v6;

always @(posedge FCLK) Cnfh07 <= Htk7v6;
always @(posedge FCLK) Apfh07 <= Atk7v6;
always @(posedge FCLK) Yqfh07 <= Tsk7v6;
always @(posedge FCLK) Wsfh07 <= Msk7v6;
always @(posedge FCLK) Yufh07 <= Fsk7v6;
always @(posedge FCLK) Axfh07 <= Yrk7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Czfh07 <= 1'b0;
  else
    Czfh07 <= Rrk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    H1gh07 <= 1'b0;
  else
    H1gh07 <= Krk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    N3gh07 <= 1'b0;
  else
    N3gh07 <= Drk7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    T5gh07 <= 1'b0;
  else
    T5gh07 <= Wqk7v6;

always @(posedge FCLK) Z7gh07 <= Pqk7v6;
always @(posedge FCLK) Bagh07 <= Iqk7v6;
always @(posedge FCLK) Ecgh07 <= Bqk7v6;
always @(posedge FCLK) Hegh07 <= Upk7v6;
always @(posedge FCLK) Kggh07 <= Npk7v6;
always @(posedge FCLK) Nigh07 <= Gpk7v6;
always @(posedge FCLK) Qkgh07 <= Zok7v6;
always @(posedge FCLK) Tmgh07 <= Sok7v6;
always @(posedge FCLK) Wogh07 <= Lok7v6;
always @(posedge FCLK) Zqgh07 <= Eok7v6;
always @(posedge FCLK) Ctgh07 <= Xnk7v6;
always @(posedge FCLK) Fvgh07 <= Qnk7v6;
always @(posedge FCLK) Ixgh07 <= Jnk7v6;
always @(posedge FCLK) Lzgh07 <= Cnk7v6;
always @(posedge FCLK) O1hh07 <= Vmk7v6;
always @(posedge FCLK) R3hh07 <= Omk7v6;
always @(posedge FCLK) U5hh07 <= Hmk7v6;
always @(posedge FCLK) X7hh07 <= Amk7v6;
always @(posedge FCLK) Aahh07 <= Tlk7v6;
always @(posedge FCLK) Dchh07 <= Mlk7v6;
always @(posedge FCLK) Gehh07 <= Flk7v6;
always @(posedge FCLK) Jghh07 <= Ykk7v6;
always @(posedge FCLK) Mihh07 <= Rkk7v6;
always @(posedge FCLK) Pkhh07 <= Kkk7v6;
always @(posedge FCLK) Rmhh07 <= Dkk7v6;
always @(posedge FCLK) Tohh07 <= Wjk7v6;
always @(posedge FCLK) Vqhh07 <= Pjk7v6;
always @(posedge FCLK) Xshh07 <= Ijk7v6;
always @(posedge FCLK) Zuhh07 <= Bjk7v6;
always @(posedge FCLK) Bxhh07 <= Uik7v6;
always @(posedge FCLK) Dzhh07 <= Nik7v6;
always @(posedge FCLK) F1ih07 <= Gik7v6;
always @(posedge FCLK) H3ih07 <= Zhk7v6;
always @(posedge FCLK) J5ih07 <= Shk7v6;
always @(posedge FCLK) L7ih07 <= Lhk7v6;
always @(posedge FCLK) N9ih07 <= Ehk7v6;
always @(posedge FCLK) Pbih07 <= Xgk7v6;
always @(posedge FCLK) Rdih07 <= Qgk7v6;
always @(posedge FCLK) Tfih07 <= Jgk7v6;
always @(posedge FCLK) Vhih07 <= Cgk7v6;
always @(posedge FCLK) Yjih07 <= Vfk7v6;
always @(posedge FCLK) Bmih07 <= Ofk7v6;
always @(posedge FCLK) Eoih07 <= Hfk7v6;
always @(posedge FCLK) Hqih07 <= Afk7v6;
always @(posedge FCLK) Ksih07 <= Tek7v6;
always @(posedge FCLK) Nuih07 <= Mek7v6;
always @(posedge FCLK) Qwih07 <= Fek7v6;
always @(posedge FCLK) Tyih07 <= Ydk7v6;
always @(posedge FCLK) W0jh07 <= Rdk7v6;
always @(posedge FCLK) Z2jh07 <= Kdk7v6;
always @(posedge FCLK) C5jh07 <= Ddk7v6;
always @(posedge FCLK) F7jh07 <= Wck7v6;
always @(posedge FCLK) I9jh07 <= Pck7v6;
always @(posedge FCLK) Lbjh07 <= Ick7v6;
always @(posedge FCLK) Odjh07 <= Bck7v6;
always @(posedge FCLK) Rfjh07 <= Ubk7v6;
always @(posedge FCLK) Uhjh07 <= Nbk7v6;
always @(posedge FCLK) Xjjh07 <= Gbk7v6;
always @(posedge FCLK) Amjh07 <= Zak7v6;
always @(posedge FCLK) Dojh07 <= Sak7v6;
always @(posedge FCLK) Gqjh07 <= Lak7v6;
always @(posedge FCLK) Jsjh07 <= Eak7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lujh07 <= 1'b0;
  else
    Lujh07 <= X9k7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qwjh07 <= 1'b0;
  else
    Qwjh07 <= Q9k7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wyjh07 <= 1'b0;
  else
    Wyjh07 <= J9k7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    C1kh07 <= 1'b0;
  else
    C1kh07 <= C9k7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    I3kh07 <= 1'b0;
  else
    I3kh07 <= V8k7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Q5kh07 <= 1'b0;
  else
    Q5kh07 <= O8k7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    C8kh07 <= 1'b0;
  else
    C8kh07 <= H8k7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Oakh07 <= 1'b0;
  else
    Oakh07 <= A8k7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Adkh07 <= 1'b0;
  else
    Adkh07 <= T7k7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mfkh07 <= 1'b0;
  else
    Mfkh07 <= M7k7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Uhkh07 <= 1'b0;
  else
    Uhkh07 <= F7k7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ckkh07 <= 1'b0;
  else
    Ckkh07 <= Zt78v6;

always @(posedge HCLK) Ylkh07 <= Y6k7v6;
always @(posedge HCLK) Nnkh07 <= R6k7v6;
always @(posedge HCLK) Fqkh07 <= K6k7v6;
always @(posedge HCLK) Xskh07 <= D6k7v6;
always @(posedge HCLK) Pvkh07 <= W5k7v6;
always @(posedge HCLK) Hykh07 <= P5k7v6;
always @(posedge HCLK) Z0lh07 <= I5k7v6;
always @(posedge HCLK) R3lh07 <= B5k7v6;
always @(posedge HCLK) J6lh07 <= U4k7v6;
always @(posedge HCLK) B9lh07 <= N4k7v6;
always @(posedge HCLK) Tblh07 <= G4k7v6;
always @(posedge HCLK) Kelh07 <= Z3k7v6;
always @(posedge HCLK) Bhlh07 <= S3k7v6;
always @(posedge HCLK) Sjlh07 <= L3k7v6;
always @(posedge HCLK) Jmlh07 <= E3k7v6;
always @(posedge HCLK) Aplh07 <= X2k7v6;
always @(posedge HCLK) Rrlh07 <= Q2k7v6;
always @(posedge HCLK) Iulh07 <= J2k7v6;
always @(posedge HCLK) Zwlh07 <= C2k7v6;
always @(posedge HCLK) Qzlh07 <= V1k7v6;
always @(posedge HCLK) Z1mh07 <= O1k7v6;
always @(posedge HCLK) I4mh07 <= H1k7v6;
always @(posedge HCLK) Q6mh07 <= A1k7v6;
always @(posedge HCLK) Y8mh07 <= T0k7v6;
always @(posedge HCLK) Gbmh07 <= M0k7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pdmh07 <= 1'b0;
  else
    Pdmh07 <= F0k7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yfmh07 <= 1'b0;
  else
    Yfmh07 <= E8l8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rhmh07 <= 1'b0;
  else
    Rhmh07 <= Yzj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wjmh07 <= 1'b0;
  else
    Wjmh07 <= Rzj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bmmh07 <= 1'b0;
  else
    Bmmh07 <= Kzj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gomh07 <= 1'b0;
  else
    Gomh07 <= Dzj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lqmh07 <= 1'b0;
  else
    Lqmh07 <= Wyj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qsmh07 <= 1'b0;
  else
    Qsmh07 <= Pyj7v6;

always @(posedge HCLK) Vumh07 <= Iyj7v6;
always @(posedge HCLK) Dxmh07 <= Byj7v6;
always @(posedge HCLK) Lzmh07 <= Uxj7v6;
always @(posedge HCLK) T1nh07 <= Nxj7v6;
always @(posedge HCLK) B4nh07 <= Gxj7v6;
always @(posedge HCLK) J6nh07 <= Zwj7v6;
always @(posedge HCLK) R8nh07 <= Swj7v6;
always @(posedge HCLK) Zanh07 <= Lwj7v6;
always @(posedge HCLK) Idnh07 <= Ewj7v6;
always @(posedge HCLK) Rfnh07 <= Xvj7v6;
always @(posedge HCLK) Ainh07 <= Qvj7v6;
always @(posedge HCLK) Jknh07 <= Jvj7v6;
always @(posedge HCLK) Smnh07 <= Cvj7v6;
always @(posedge HCLK) Bpnh07 <= Vuj7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jrnh07 <= 1'b1;
  else
    Jrnh07 <= Ouj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Etnh07 <= 1'b0;
  else
    Etnh07 <= Huj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zunh07 <= 1'b0;
  else
    Zunh07 <= Auj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Uwnh07 <= 1'b0;
  else
    Uwnh07 <= Ttj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pynh07 <= 1'b0;
  else
    Pynh07 <= Mtj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    K0oh07 <= 1'b0;
  else
    K0oh07 <= Ftj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F2oh07 <= 1'b0;
  else
    F2oh07 <= Ysj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    U3oh07 <= 1'b0;
  else
    U3oh07 <= Vr78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    P5oh07 <= 1'b1;
  else
    P5oh07 <= Rsj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    G7oh07 <= 1'b0;
  else
    G7oh07 <= C477v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    B9oh07 <= 1'b0;
  else
    B9oh07 <= Vxu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kboh07 <= 1'b1;
  else
    Kboh07 <= Osk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Idoh07 <= 1'b1;
  else
    Idoh07 <= Suk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gfoh07 <= 1'b1;
  else
    Gfoh07 <= Vsk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ehoh07 <= 1'b1;
  else
    Ehoh07 <= Ctk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cjoh07 <= 1'b1;
  else
    Cjoh07 <= Jtk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Aloh07 <= 1'b1;
  else
    Aloh07 <= Qtk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ymoh07 <= 1'b1;
  else
    Ymoh07 <= Xtk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wooh07 <= 1'b1;
  else
    Wooh07 <= Euk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Uqoh07 <= 1'b1;
  else
    Uqoh07 <= Luk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ssoh07 <= 1'b0;
  else
    Ssoh07 <= Yjd8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ruoh07 <= 1'b0;
  else
    Ruoh07 <= Sa77v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pwoh07 <= 1'b0;
  else
    Pwoh07 <= Ru77v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wyoh07 <= 1'b0;
  else
    Wyoh07 <= Ksj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    W0ph07 <= 1'b0;
  else
    W0ph07 <= Dsj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    U2ph07 <= 1'b1;
  else
    U2ph07 <= Wrj7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R4ph07 <= 1'b0;
  else
    R4ph07 <= Qyu7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T6ph07 <= 1'b0;
  else
    T6ph07 <= Xyu7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W8ph07 <= 1'b0;
  else
    W8ph07 <= F848v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bbph07 <= 1'b0;
  else
    Bbph07 <= M848v6;

always @(posedge FCLK) Gdph07 <= Prj7v6;
always @(posedge FCLK) Qfph07 <= Y748v6;
always @(posedge FCLK) Aiph07 <= R748v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kkph07 <= 1'b0;
  else
    Kkph07 <= S3adt6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Emph07 <= 1'b0;
  else
    Emph07 <= T848v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Joph07 <= 1'b0;
  else
    Joph07 <= Kwl8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hqph07 <= 1'b0;
  else
    Hqph07 <= Tfx7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lsph07 <= 1'b0;
  else
    Lsph07 <= Lua7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vuph07 <= 1'b0;
  else
    Vuph07 <= Gsa7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ixph07 <= 1'b0;
  else
    Ixph07 <= Pma7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pzph07 <= 1'b0;
  else
    Pzph07 <= J2b7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    R1qh07 <= 1'b0;
  else
    R1qh07 <= Y5a7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Z3qh07 <= 1'b0;
  else
    Z3qh07 <= Mqa7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F6qh07 <= 1'b0;
  else
    F6qh07 <= Dwl8v6;

always @(posedge FCLK) D8qh07 <= Irj7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Oaqh07 <= 1'b0;
  else
    Oaqh07 <= Rex7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Scqh07 <= 1'b0;
  else
    Scqh07 <= Zxymz6[8];

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zeqh07 <= 1'b0;
  else
    Zeqh07 <= Ezu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dhqh07 <= 1'b1;
  else
    Dhqh07 <= Wy67v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ejqh07 <= 1'b0;
  else
    Ejqh07 <= Jyu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zkqh07 <= 1'b0;
  else
    Zkqh07 <= Drymz6[1];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fnqh07 <= 1'b0;
  else
    Fnqh07 <= Frc7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Woqh07 <= 1'b0;
  else
    Woqh07 <= Cyu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Uqqh07 <= 1'b0;
  else
    Uqqh07 <= Br77v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vsqh07 <= 1'b0;
  else
    Vsqh07 <= Brj7v6;

always @(posedge HCLK) Nuqh07 <= Uqj7v6;
always @(posedge HCLK) Lwqh07 <= Nqj7v6;
always @(posedge HCLK) Kyqh07 <= Gqj7v6;
always @(posedge HCLK) J0rh07 <= Zpj7v6;
always @(posedge HCLK) I2rh07 <= Spj7v6;
always @(posedge HCLK) H4rh07 <= Lpj7v6;
always @(posedge HCLK) G6rh07 <= Epj7v6;
always @(posedge HCLK) F8rh07 <= Xoj7v6;
always @(posedge HCLK) Earh07 <= Qoj7v6;
always @(posedge HCLK) Dcrh07 <= Joj7v6;
always @(posedge HCLK) Cerh07 <= Coj7v6;
always @(posedge HCLK) Bgrh07 <= Vnj7v6;
always @(posedge HCLK) Airh07 <= Onj7v6;
always @(posedge HCLK) Zjrh07 <= Hnj7v6;
always @(posedge HCLK) Ylrh07 <= Anj7v6;
always @(posedge HCLK) Xnrh07 <= Tmj7v6;
always @(posedge HCLK) Wprh07 <= Mmj7v6;
always @(posedge HCLK) Vrrh07 <= Fmj7v6;
always @(posedge HCLK) Gxps07 <= Ylj7v6;
always @(posedge HCLK) Fzps07 <= Rlj7v6;
always @(posedge HCLK) E1qs07 <= Klj7v6;
always @(posedge HCLK) D3qs07 <= Dlj7v6;
always @(posedge HCLK) C5qs07 <= Wkj7v6;
always @(posedge HCLK) B7qs07 <= Pkj7v6;
always @(posedge HCLK) A9qs07 <= Ikj7v6;
always @(posedge HCLK) Zaqs07 <= Bkj7v6;
always @(posedge HCLK) Ycqs07 <= Ujj7v6;
always @(posedge HCLK) Xeqs07 <= Njj7v6;
always @(posedge HCLK) Wgqs07 <= Gjj7v6;
always @(posedge HCLK) Viqs07 <= Zij7v6;
always @(posedge HCLK) Ukqs07 <= Sij7v6;
always @(posedge HCLK) Tmqs07 <= Lij7v6;
always @(posedge HCLK) Soqs07 <= Eij7v6;
always @(posedge HCLK) Rqqs07 <= Xhj7v6;
always @(posedge HCLK) Qsqs07 <= Qhj7v6;
always @(posedge HCLK) Puqs07 <= Jhj7v6;
always @(posedge HCLK) Owqs07 <= Chj7v6;
always @(posedge HCLK) Nyqs07 <= Vgj7v6;
always @(posedge HCLK) M0rs07 <= Ogj7v6;
always @(posedge HCLK) L2rs07 <= Hgj7v6;
always @(posedge HCLK) K4rs07 <= Agj7v6;
always @(posedge HCLK) I6rs07 <= Tfj7v6;
always @(posedge HCLK) G8rs07 <= Mfj7v6;
always @(posedge HCLK) Ears07 <= Ffj7v6;
always @(posedge HCLK) Ccrs07 <= Yej7v6;
always @(posedge HCLK) Aers07 <= Rej7v6;
always @(posedge HCLK) Yfrs07 <= Kej7v6;
always @(posedge HCLK) Whrs07 <= Dej7v6;
always @(posedge HCLK) Ujrs07 <= Wdj7v6;
always @(posedge HCLK) Dmrs07 <= Pdj7v6;
always @(posedge HCLK) Mors07 <= Idj7v6;
always @(posedge HCLK) Vqrs07 <= Bdj7v6;
always @(posedge HCLK) Etrs07 <= Ucj7v6;
always @(posedge HCLK) Nvrs07 <= Ncj7v6;
always @(posedge HCLK) Wxrs07 <= Gcj7v6;
always @(posedge HCLK) F0ss07 <= Zbj7v6;
always @(posedge HCLK) O2ss07 <= Sbj7v6;
always @(posedge HCLK) X4ss07 <= Lbj7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    L7ss07 <= 1'b0;
  else
    L7ss07 <= Twu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    G9ss07 <= 1'b0;
  else
    G9ss07 <= Hxu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bbss07 <= 1'b0;
  else
    Bbss07 <= Oxu7v6;

always @(posedge HCLK) Wcss07 <= Ebj7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tess07 <= 1'b0;
  else
    Tess07 <= Ce78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ngss07 <= 1'b0;
  else
    Ngss07 <= Qe78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hiss07 <= 1'b0;
  else
    Hiss07 <= Xe78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bkss07 <= 1'b0;
  else
    Bkss07 <= Sf78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cmss07 <= 1'b1;
  else
    Cmss07 <= Hk78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Aoss07 <= 1'b0;
  else
    Aoss07 <= Ak78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ypss07 <= 1'b0;
  else
    Ypss07 <= Ok78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vrss07 <= 1'b0;
  else
    Vrss07 <= Cl78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Stss07 <= 1'b0;
  else
    Stss07 <= Xl78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pvss07 <= 1'b0;
  else
    Pvss07 <= Em78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mxss07 <= 1'b0;
  else
    Mxss07 <= Zm78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kzss07 <= 1'b0;
  else
    Kzss07 <= Gn78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    I1ts07 <= 1'b0;
  else
    I1ts07 <= Nn78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    G3ts07 <= 1'b0;
  else
    G3ts07 <= Un78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    C5ts07 <= 1'b0;
  else
    C5ts07 <= Nyd7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    P7ts07 <= 1'b0;
  else
    P7ts07 <= N6h7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Cats07 <= 1'b0;
  else
    Cats07 <= M7e7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Fcts07 <= 1'b0;
  else
    Fcts07 <= Fj78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Dets07 <= 1'b0;
  else
    Dets07 <= Yi78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Bgts07 <= 1'b0;
  else
    Bgts07 <= Ri78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Zhts07 <= 1'b0;
  else
    Zhts07 <= Ki78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Xjts07 <= 1'b0;
  else
    Xjts07 <= Di78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Vlts07 <= 1'b0;
  else
    Vlts07 <= Wh78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Tnts07 <= 1'b0;
  else
    Tnts07 <= Ph78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Rpts07 <= 1'b0;
  else
    Rpts07 <= Ih78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Prts07 <= 1'b0;
  else
    Prts07 <= Bh78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Ntts07 <= 1'b0;
  else
    Ntts07 <= Ug78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Mvts07 <= 1'b0;
  else
    Mvts07 <= Ng78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Lxts07 <= 1'b0;
  else
    Lxts07 <= Gg78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kzts07 <= 1'b0;
  else
    Kzts07 <= Bo78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    H1us07 <= 1'b0;
  else
    H1us07 <= Sm78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    E3us07 <= 1'b1;
  else
    E3us07 <= Zf78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    D5us07 <= 1'b0;
  else
    D5us07 <= Io78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F7us07 <= 1'b0;
  else
    F7us07 <= Po78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    C9us07 <= 1'b1;
  else
    C9us07 <= Wo78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ebus07 <= 1'b0;
  else
    Ebus07 <= Lf78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fdus07 <= 1'b0;
  else
    Fdus07 <= Ef78v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gfus07 <= 1'b0;
  else
    Gfus07 <= Qur7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Thus07 <= 1'b0;
  else
    Thus07 <= Ja1nz6[0];

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Mkus07 <= 1'b0;
  else
    Mkus07 <= Brg7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fnus07 <= 1'b0;
  else
    Fnus07 <= Xaj7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lous07 <= 1'b1;
  else
    Lous07 <= Ysx7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bqus07 <= 1'b1;
  else
    Bqus07 <= Qaj7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Prus07 <= 1'b0;
  else
    Prus07 <= Jaj7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ntus07 <= 1'b0;
  else
    Ntus07 <= Caj7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mvus07 <= 1'b0;
  else
    Mvus07 <= Amr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kxus07 <= 1'b0;
  else
    Kxus07 <= Dbl8v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Xzus07 <= 1'b0;
  else
    Xzus07 <= U81nz6[0];

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Q2vs07 <= 1'b0;
  else
    Q2vs07 <= Uyg7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    J5vs07 <= 1'b0;
  else
    J5vs07 <= Ahp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    H7vs07 <= 1'b0;
  else
    H7vs07 <= Cip7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F9vs07 <= 1'b0;
  else
    F9vs07 <= Ejp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dbvs07 <= 1'b0;
  else
    Dbvs07 <= Gkp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bdvs07 <= 1'b0;
  else
    Bdvs07 <= Ilp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zevs07 <= 1'b0;
  else
    Zevs07 <= Pal8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xgvs07 <= 1'b0;
  else
    Xgvs07 <= Hhp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vivs07 <= 1'b0;
  else
    Vivs07 <= Jip7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tkvs07 <= 1'b0;
  else
    Tkvs07 <= Ljp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rmvs07 <= 1'b0;
  else
    Rmvs07 <= Nkp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Povs07 <= 1'b0;
  else
    Povs07 <= Plp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Nqvs07 <= 1'b0;
  else
    Nqvs07 <= Bal8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lsvs07 <= 1'b0;
  else
    Lsvs07 <= N9l8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Juvs07 <= 1'b0;
  else
    Juvs07 <= U9l8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hwvs07 <= 1'b0;
  else
    Hwvs07 <= Vd78v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Uyvs07 <= 1'b0;
  else
    Uyvs07 <= U81nz6[2];

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    N1ws07 <= 1'b0;
  else
    N1ws07 <= Y3h7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    G4ws07 <= 1'b0;
  else
    G4ws07 <= V9j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    X5ws07 <= 1'b0;
  else
    X5ws07 <= O9j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    O7ws07 <= 1'b0;
  else
    O7ws07 <= H9j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F9ws07 <= 1'b0;
  else
    F9ws07 <= A9j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Waws07 <= 1'b0;
  else
    Waws07 <= T8j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ncws07 <= 1'b0;
  else
    Ncws07 <= M8j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Eews07 <= 1'b0;
  else
    Eews07 <= F8j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wfws07 <= 1'b0;
  else
    Wfws07 <= Y7j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yhws07 <= 1'b0;
  else
    Yhws07 <= R7j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qjws07 <= 1'b0;
  else
    Qjws07 <= K7j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ilws07 <= 1'b0;
  else
    Ilws07 <= D7j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lnws07 <= 1'b0;
  else
    Lnws07 <= W6j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hpws07 <= 1'b0;
  else
    Hpws07 <= P6j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Drws07 <= 1'b0;
  else
    Drws07 <= I6j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Atws07 <= 1'b0;
  else
    Atws07 <= B6j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xuws07 <= 1'b0;
  else
    Xuws07 <= U5j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Uwws07 <= 1'b0;
  else
    Uwws07 <= N5j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tyws07 <= 1'b0;
  else
    Tyws07 <= G5j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    S0xs07 <= 1'b0;
  else
    S0xs07 <= Z4j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    R2xs07 <= 1'b0;
  else
    R2xs07 <= S4j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Q4xs07 <= 1'b0;
  else
    Q4xs07 <= L4j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    P6xs07 <= 1'b0;
  else
    P6xs07 <= E4j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    O8xs07 <= 1'b0;
  else
    O8xs07 <= X3j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Naxs07 <= 1'b0;
  else
    Naxs07 <= Q3j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mcxs07 <= 1'b0;
  else
    Mcxs07 <= J3j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lexs07 <= 1'b0;
  else
    Lexs07 <= C3j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kgxs07 <= 1'b0;
  else
    Kgxs07 <= V2j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jixs07 <= 1'b0;
  else
    Jixs07 <= O2j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ikxs07 <= 1'b0;
  else
    Ikxs07 <= H2j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hmxs07 <= 1'b0;
  else
    Hmxs07 <= A2j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Goxs07 <= 1'b0;
  else
    Goxs07 <= T1j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fqxs07 <= 1'b0;
  else
    Fqxs07 <= M1j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Esxs07 <= 1'b0;
  else
    Esxs07 <= F1j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Duxs07 <= 1'b0;
  else
    Duxs07 <= Y0j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cwxs07 <= 1'b0;
  else
    Cwxs07 <= R0j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Byxs07 <= 1'b0;
  else
    Byxs07 <= K0j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    A0ys07 <= 1'b0;
  else
    A0ys07 <= D0j7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Z1ys07 <= 1'b0;
  else
    Z1ys07 <= Wzi7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y3ys07 <= 1'b0;
  else
    Y3ys07 <= P4k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V6ys07 <= 1'b0;
  else
    V6ys07 <= Rcs7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y9ys07 <= 1'b0;
  else
    Y9ys07 <= Kcs7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bdys07 <= 1'b0;
  else
    Bdys07 <= Pbs7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Egys07 <= 1'b0;
  else
    Egys07 <= Z9s7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ijys07 <= 1'b0;
  else
    Ijys07 <= L9s7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mmys07 <= 1'b0;
  else
    Mmys07 <= E9s7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qpys07 <= 1'b0;
  else
    Qpys07 <= X8s7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Usys07 <= 1'b0;
  else
    Usys07 <= V7s7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yvys07 <= 1'b0;
  else
    Yvys07 <= T6s7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Czys07 <= 1'b0;
  else
    Czys07 <= M6s7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    G2zs07 <= 1'b0;
  else
    G2zs07 <= T7j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D5zs07 <= 1'b0;
  else
    D5zs07 <= Nok8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M7zs07 <= 1'b0;
  else
    M7zs07 <= Svy7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W9zs07 <= 1'b0;
  else
    W9zs07 <= Gwy7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gczs07 <= 1'b0;
  else
    Gczs07 <= Dyy7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qezs07 <= 1'b0;
  else
    Qezs07 <= Ryy7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ahzs07 <= 1'b0;
  else
    Ahzs07 <= Tzy7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kjzs07 <= 1'b0;
  else
    Kjzs07 <= H0z7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ulzs07 <= 1'b0;
  else
    Ulzs07 <= X1z7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Eozs07 <= 1'b0;
  else
    Eozs07 <= L2z7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oqzs07 <= 1'b0;
  else
    Oqzs07 <= N3z7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yszs07 <= 1'b0;
  else
    Yszs07 <= B4z7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hvzs07 <= 1'b0;
  else
    Hvzs07 <= P4z7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rxzs07 <= 1'b0;
  else
    Rxzs07 <= D5z7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B00t07 <= 1'b0;
  else
    B00t07 <= R5z7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L20t07 <= 1'b0;
  else
    L20t07 <= I738v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V40t07 <= 1'b0;
  else
    V40t07 <= P738v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F70t07 <= 1'b0;
  else
    F70t07 <= Kck8v6;

always @(posedge HCLK) O90t07 <= Ddy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lc0t07 <= 1'b0;
  else
    Lc0t07 <= Fyk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ve0t07 <= 1'b0;
  else
    Ve0t07 <= Aui8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sh0t07 <= 1'b0;
  else
    Sh0t07 <= Agi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dk0t07 <= 1'b0;
  else
    Dk0t07 <= Nk38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gm0t07 <= 1'b0;
  else
    Gm0t07 <= Uk38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lo0t07 <= 1'b0;
  else
    Lo0t07 <= B3l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kr0t07 <= 1'b0;
  else
    Kr0t07 <= Uvs7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ju0t07 <= 1'b0;
  else
    Ju0t07 <= Bws7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ix0t07 <= 1'b0;
  else
    Ix0t07 <= Chi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L01t07 <= 1'b0;
  else
    L01t07 <= Y838v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M31t07 <= 1'b0;
  else
    M31t07 <= Jhi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J61t07 <= 1'b0;
  else
    J61t07 <= Rei8v6;

always @(posedge HCLK) G91t07 <= F1i8v6;
always @(posedge HCLK) Lb1t07 <= R0i8v6;
always @(posedge HCLK) Qd1t07 <= Cbp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tg1t07 <= 1'b0;
  else
    Tg1t07 <= Pzi7v6;

always @(posedge FCLK) Qi1t07 <= Izi7v6;
always @(posedge FCLK) Sk1t07 <= Bzi7v6;
always @(posedge FCLK) Um1t07 <= Uyi7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wo1t07 <= 1'b0;
  else
    Wo1t07 <= Nyi7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cr1t07 <= 1'b0;
  else
    Cr1t07 <= Da88v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jt1t07 <= 1'b0;
  else
    Jt1t07 <= Gyi7v6;

always @(posedge FCLK) Pv1t07 <= Zxi7v6;
always @(posedge FCLK) Nx1t07 <= Sxi7v6;
always @(posedge FCLK) Lz1t07 <= Lxi7v6;
always @(posedge FCLK) N12t07 <= Exi7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    P32t07 <= 1'b0;
  else
    P32t07 <= Xwi7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    R52t07 <= 1'b0;
  else
    R52t07 <= Ohw7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Z72t07 <= 1'b0;
  else
    Z72t07 <= Kfw7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ba2t07 <= 1'b0;
  else
    Ba2t07 <= Ahw7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ac2t07 <= 1'b0;
  else
    Ac2t07 <= Qwi7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ge2t07 <= 1'b0;
  else
    Ge2t07 <= Ra88v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fg2t07 <= 1'b0;
  else
    Fg2t07 <= Ya88v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Li2t07 <= 1'b0;
  else
    Li2t07 <= Ka88v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tk2t07 <= 1'b0;
  else
    Tk2t07 <= Dfw7v6;

always @(posedge FCLK) Vm2t07 <= Jwi7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xo2t07 <= 1'b0;
  else
    Xo2t07 <= W988v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Er2t07 <= 1'b0;
  else
    Er2t07 <= Cwi7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    It2t07 <= 1'b0;
  else
    It2t07 <= Vvi7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pv2t07 <= 1'b0;
  else
    Pv2t07 <= Mzj8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ox2t07 <= 1'b0;
  else
    Ox2t07 <= Ovi7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qz2t07 <= 1'b0;
  else
    Qz2t07 <= Od78v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    J23t07 <= 1'b0;
  else
    J23t07 <= Hd78v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    K33t07 <= 1'b0;
  else
    K33t07 <= Hcget6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J43t07 <= 1'b0;
  else
    J43t07 <= Hvi7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K63t07 <= 1'b0;
  else
    K63t07 <= Avi7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q83t07 <= 1'b0;
  else
    Q83t07 <= Tui7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pa3t07 <= 1'b0;
  else
    Pa3t07 <= Mui7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pc3t07 <= 1'b0;
  else
    Pc3t07 <= Fui7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qe3t07 <= 1'b0;
  else
    Qe3t07 <= Yti7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ug3t07 <= 1'b0;
  else
    Ug3t07 <= Rti7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ni3t07 <= 1'b0;
  else
    Ni3t07 <= Kti7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kk3t07 <= 1'b0;
  else
    Kk3t07 <= Dti7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jm3t07 <= 1'b0;
  else
    Jm3t07 <= Wsi7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Io3t07 <= 1'b0;
  else
    Io3t07 <= Psi7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hq3t07 <= 1'b0;
  else
    Hq3t07 <= Isi7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gs3t07 <= 1'b0;
  else
    Gs3t07 <= Bsi7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fu3t07 <= 1'b0;
  else
    Fu3t07 <= Uri7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ew3t07 <= 1'b0;
  else
    Ew3t07 <= Nri7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dy3t07 <= 1'b0;
  else
    Dy3t07 <= Gri7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    C04t07 <= 1'b0;
  else
    C04t07 <= Zqi7v6;

always @(posedge HCLK) H24t07 <= Sqi7v6;
always @(posedge HCLK) Q44t07 <= Lqi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y64t07 <= 1'b0;
  else
    Y64t07 <= Mi88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V94t07 <= 1'b0;
  else
    V94t07 <= Ti88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sc4t07 <= 1'b1;
  else
    Sc4t07 <= Gwc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pf4t07 <= 1'b0;
  else
    Pf4t07 <= Nwc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mi4t07 <= 1'b0;
  else
    Mi4t07 <= Wcc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ik4t07 <= 1'b0;
  else
    Ik4t07 <= Hw98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zn4t07 <= 1'b0;
  else
    Zn4t07 <= Zr98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qr4t07 <= 1'b0;
  else
    Qr4t07 <= Yn98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hv4t07 <= 1'b0;
  else
    Hv4t07 <= Mh98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vy4t07 <= 1'b0;
  else
    Vy4t07 <= F9a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N25t07 <= 1'b0;
  else
    N25t07 <= Nda8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F65t07 <= 1'b0;
  else
    F65t07 <= Vha8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X95t07 <= 1'b0;
  else
    X95t07 <= Dma8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pd5t07 <= 1'b0;
  else
    Pd5t07 <= X4a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hh5t07 <= 1'b0;
  else
    Hh5t07 <= R7b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tk5t07 <= 1'b0;
  else
    Tk5t07 <= Zbb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fo5t07 <= 1'b0;
  else
    Fo5t07 <= Hgb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rr5t07 <= 1'b0;
  else
    Rr5t07 <= Pkb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dv5t07 <= 1'b0;
  else
    Dv5t07 <= J3b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Py5t07 <= 1'b0;
  else
    Py5t07 <= Bza8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B26t07 <= 1'b0;
  else
    B26t07 <= Tua8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N56t07 <= 1'b0;
  else
    N56t07 <= Vb98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z86t07 <= 1'b0;
  else
    Z86t07 <= Zd98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lc6t07 <= 1'b0;
  else
    Lc6t07 <= Fh98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xf6t07 <= 1'b0;
  else
    Xf6t07 <= Lk98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jj6t07 <= 1'b0;
  else
    Jj6t07 <= Rn98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vm6t07 <= 1'b0;
  else
    Vm6t07 <= Sr98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hq6t07 <= 1'b0;
  else
    Hq6t07 <= Aw98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tt6t07 <= 1'b0;
  else
    Tt6t07 <= R998v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fx6t07 <= 1'b0;
  else
    Fx6t07 <= K1a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R07t07 <= 1'b0;
  else
    R07t07 <= Q4a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D47t07 <= 1'b0;
  else
    D47t07 <= Wla8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P77t07 <= 1'b0;
  else
    P77t07 <= Oha8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bb7t07 <= 1'b0;
  else
    Bb7t07 <= Gda8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ne7t07 <= 1'b0;
  else
    Ne7t07 <= Y8a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zh7t07 <= 1'b0;
  else
    Zh7t07 <= Mua8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ll7t07 <= 1'b0;
  else
    Ll7t07 <= Uya8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xo7t07 <= 1'b0;
  else
    Xo7t07 <= C3b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Js7t07 <= 1'b0;
  else
    Js7t07 <= Ikb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uv7t07 <= 1'b0;
  else
    Uv7t07 <= Agb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gz7t07 <= 1'b0;
  else
    Gz7t07 <= Sbb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    S28t07 <= 1'b0;
  else
    S28t07 <= K7b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    E68t07 <= 1'b0;
  else
    E68t07 <= Gxb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P98t07 <= 1'b0;
  else
    P98t07 <= Aub8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ad8t07 <= 1'b0;
  else
    Ad8t07 <= Wrb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lg8t07 <= 1'b0;
  else
    Lg8t07 <= C9c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tj8t07 <= 1'b0;
  else
    Tj8t07 <= Y6c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gn8t07 <= 1'b0;
  else
    Gn8t07 <= Q2c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tq8t07 <= 1'b0;
  else
    Tq8t07 <= M0c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gu8t07 <= 1'b0;
  else
    Gu8t07 <= Nxb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tx8t07 <= 1'b0;
  else
    Tx8t07 <= Vw98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K19t07 <= 1'b0;
  else
    K19t07 <= Ns98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B59t07 <= 1'b0;
  else
    B59t07 <= Mo98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    S89t07 <= 1'b0;
  else
    S89t07 <= Ai98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gc9t07 <= 1'b0;
  else
    Gc9t07 <= T9a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yf9t07 <= 1'b0;
  else
    Yf9t07 <= Bea8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qj9t07 <= 1'b0;
  else
    Qj9t07 <= Jia8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    In9t07 <= 1'b0;
  else
    In9t07 <= Rma8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ar9t07 <= 1'b0;
  else
    Ar9t07 <= L5a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Su9t07 <= 1'b0;
  else
    Su9t07 <= F8b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ey9t07 <= 1'b0;
  else
    Ey9t07 <= Ncb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q1at07 <= 1'b0;
  else
    Q1at07 <= Vgb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    C5at07 <= 1'b0;
  else
    C5at07 <= Dlb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O8at07 <= 1'b0;
  else
    O8at07 <= X3b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Acat07 <= 1'b0;
  else
    Acat07 <= Pza8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mfat07 <= 1'b0;
  else
    Mfat07 <= Hva8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yiat07 <= 1'b0;
  else
    Yiat07 <= Cc98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kmat07 <= 1'b0;
  else
    Kmat07 <= Ge98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wpat07 <= 1'b0;
  else
    Wpat07 <= Th98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Itat07 <= 1'b0;
  else
    Itat07 <= Sk98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uwat07 <= 1'b0;
  else
    Uwat07 <= Fo98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    G0bt07 <= 1'b0;
  else
    G0bt07 <= Gs98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    S3bt07 <= 1'b0;
  else
    S3bt07 <= Ow98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    E7bt07 <= 1'b0;
  else
    E7bt07 <= Y998v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qabt07 <= 1'b0;
  else
    Qabt07 <= R1a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cebt07 <= 1'b0;
  else
    Cebt07 <= E5a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ohbt07 <= 1'b0;
  else
    Ohbt07 <= Kma8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Albt07 <= 1'b0;
  else
    Albt07 <= Cia8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mobt07 <= 1'b0;
  else
    Mobt07 <= Uda8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yrbt07 <= 1'b0;
  else
    Yrbt07 <= M9a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kvbt07 <= 1'b0;
  else
    Kvbt07 <= Ava8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wybt07 <= 1'b0;
  else
    Wybt07 <= Iza8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    I2ct07 <= 1'b0;
  else
    I2ct07 <= Q3b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U5ct07 <= 1'b0;
  else
    U5ct07 <= Wkb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F9ct07 <= 1'b0;
  else
    F9ct07 <= Ogb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rcct07 <= 1'b0;
  else
    Rcct07 <= Gcb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dgct07 <= 1'b0;
  else
    Dgct07 <= Y7b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pjct07 <= 1'b0;
  else
    Pjct07 <= Uxb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Anct07 <= 1'b0;
  else
    Anct07 <= Hub8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lqct07 <= 1'b0;
  else
    Lqct07 <= Dsb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wtct07 <= 1'b0;
  else
    Wtct07 <= J9c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Exct07 <= 1'b0;
  else
    Exct07 <= F7c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R0dt07 <= 1'b0;
  else
    R0dt07 <= X2c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    E4dt07 <= 1'b0;
  else
    E4dt07 <= T0c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R7dt07 <= 1'b0;
  else
    R7dt07 <= Byb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ebdt07 <= 1'b0;
  else
    Ebdt07 <= Jx98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vedt07 <= 1'b0;
  else
    Vedt07 <= Bt98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Midt07 <= 1'b0;
  else
    Midt07 <= Ap98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dmdt07 <= 1'b0;
  else
    Dmdt07 <= Oi98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rpdt07 <= 1'b0;
  else
    Rpdt07 <= Haa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jtdt07 <= 1'b0;
  else
    Jtdt07 <= Pea8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bxdt07 <= 1'b0;
  else
    Bxdt07 <= Xia8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T0et07 <= 1'b0;
  else
    T0et07 <= Fna8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L4et07 <= 1'b0;
  else
    L4et07 <= Z5a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D8et07 <= 1'b0;
  else
    D8et07 <= T8b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pbet07 <= 1'b0;
  else
    Pbet07 <= Bdb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bfet07 <= 1'b0;
  else
    Bfet07 <= Jhb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Niet07 <= 1'b0;
  else
    Niet07 <= Rlb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zlet07 <= 1'b0;
  else
    Zlet07 <= L4b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lpet07 <= 1'b0;
  else
    Lpet07 <= D0b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xset07 <= 1'b0;
  else
    Xset07 <= Vva8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jwet07 <= 1'b0;
  else
    Jwet07 <= Jc98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vzet07 <= 1'b0;
  else
    Vzet07 <= Ne98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H3ft07 <= 1'b0;
  else
    H3ft07 <= Hi98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T6ft07 <= 1'b0;
  else
    T6ft07 <= Zk98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Faft07 <= 1'b0;
  else
    Faft07 <= To98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rdft07 <= 1'b0;
  else
    Rdft07 <= Us98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dhft07 <= 1'b0;
  else
    Dhft07 <= Cx98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pkft07 <= 1'b0;
  else
    Pkft07 <= Fa98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Boft07 <= 1'b0;
  else
    Boft07 <= Y1a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nrft07 <= 1'b0;
  else
    Nrft07 <= S5a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zuft07 <= 1'b0;
  else
    Zuft07 <= Yma8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lyft07 <= 1'b0;
  else
    Lyft07 <= Qia8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X1gt07 <= 1'b0;
  else
    X1gt07 <= Iea8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J5gt07 <= 1'b0;
  else
    J5gt07 <= Aaa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V8gt07 <= 1'b0;
  else
    V8gt07 <= Ova8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hcgt07 <= 1'b0;
  else
    Hcgt07 <= Wza8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tfgt07 <= 1'b0;
  else
    Tfgt07 <= E4b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fjgt07 <= 1'b0;
  else
    Fjgt07 <= Klb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qmgt07 <= 1'b0;
  else
    Qmgt07 <= Chb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cqgt07 <= 1'b0;
  else
    Cqgt07 <= Ucb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Otgt07 <= 1'b0;
  else
    Otgt07 <= M8b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Axgt07 <= 1'b0;
  else
    Axgt07 <= Iyb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L0ht07 <= 1'b0;
  else
    L0ht07 <= Oub8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W3ht07 <= 1'b0;
  else
    W3ht07 <= Ksb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H7ht07 <= 1'b0;
  else
    H7ht07 <= Q9c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Paht07 <= 1'b0;
  else
    Paht07 <= M7c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ceht07 <= 1'b0;
  else
    Ceht07 <= E3c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Phht07 <= 1'b0;
  else
    Phht07 <= A1c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Clht07 <= 1'b0;
  else
    Clht07 <= Pyb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Poht07 <= 1'b0;
  else
    Poht07 <= Xx98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gsht07 <= 1'b0;
  else
    Gsht07 <= Pt98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xvht07 <= 1'b0;
  else
    Xvht07 <= Op98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ozht07 <= 1'b0;
  else
    Ozht07 <= Cj98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    C3it07 <= 1'b0;
  else
    C3it07 <= Vaa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U6it07 <= 1'b0;
  else
    U6it07 <= Dfa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mait07 <= 1'b0;
  else
    Mait07 <= Lja8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Eeit07 <= 1'b0;
  else
    Eeit07 <= Tna8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Whit07 <= 1'b0;
  else
    Whit07 <= N6a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Olit07 <= 1'b0;
  else
    Olit07 <= H9b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Apit07 <= 1'b0;
  else
    Apit07 <= Pdb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Msit07 <= 1'b0;
  else
    Msit07 <= Xhb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yvit07 <= 1'b0;
  else
    Yvit07 <= Fmb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kzit07 <= 1'b0;
  else
    Kzit07 <= Z4b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W2jt07 <= 1'b0;
  else
    W2jt07 <= R0b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    I6jt07 <= 1'b0;
  else
    I6jt07 <= Jwa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U9jt07 <= 1'b0;
  else
    U9jt07 <= Qc98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gdjt07 <= 1'b0;
  else
    Gdjt07 <= Ue98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sgjt07 <= 1'b0;
  else
    Sgjt07 <= Vi98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ekjt07 <= 1'b0;
  else
    Ekjt07 <= Gl98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qnjt07 <= 1'b0;
  else
    Qnjt07 <= Hp98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Crjt07 <= 1'b0;
  else
    Crjt07 <= It98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oujt07 <= 1'b0;
  else
    Oujt07 <= Qx98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ayjt07 <= 1'b0;
  else
    Ayjt07 <= Ma98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M1kt07 <= 1'b0;
  else
    M1kt07 <= F2a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y4kt07 <= 1'b0;
  else
    Y4kt07 <= G6a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K8kt07 <= 1'b0;
  else
    K8kt07 <= Mna8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wbkt07 <= 1'b0;
  else
    Wbkt07 <= Eja8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ifkt07 <= 1'b0;
  else
    Ifkt07 <= Wea8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uikt07 <= 1'b0;
  else
    Uikt07 <= Oaa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gmkt07 <= 1'b0;
  else
    Gmkt07 <= Cwa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Spkt07 <= 1'b0;
  else
    Spkt07 <= K0b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Etkt07 <= 1'b0;
  else
    Etkt07 <= S4b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qwkt07 <= 1'b0;
  else
    Qwkt07 <= Ylb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B0lt07 <= 1'b0;
  else
    B0lt07 <= Qhb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N3lt07 <= 1'b0;
  else
    N3lt07 <= Idb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z6lt07 <= 1'b0;
  else
    Z6lt07 <= A9b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lalt07 <= 1'b0;
  else
    Lalt07 <= Wyb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wdlt07 <= 1'b0;
  else
    Wdlt07 <= Vub8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hhlt07 <= 1'b0;
  else
    Hhlt07 <= Rsb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sklt07 <= 1'b0;
  else
    Sklt07 <= X9c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Aolt07 <= 1'b0;
  else
    Aolt07 <= T7c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nrlt07 <= 1'b0;
  else
    Nrlt07 <= L3c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Avlt07 <= 1'b0;
  else
    Avlt07 <= H1c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nylt07 <= 1'b0;
  else
    Nylt07 <= Dzb8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    A2mt07 <= 1'b0;
  else
    A2mt07 <= Je78v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U3mt07 <= 1'b0;
  else
    U3mt07 <= F7y7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    V5mt07 <= 1'b0;
  else
    V5mt07 <= Axu7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q7mt07 <= 1'b0;
  else
    Q7mt07 <= Yyc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pamt07 <= 1'b0;
  else
    Pamt07 <= Kyc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Scmt07 <= 1'b0;
  else
    Scmt07 <= Ryc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uemt07 <= 1'b0;
  else
    Uemt07 <= Fi88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rhmt07 <= 1'b0;
  else
    Rhmt07 <= Fv98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ilmt07 <= 1'b0;
  else
    Ilmt07 <= Xq98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zomt07 <= 1'b0;
  else
    Zomt07 <= Wm98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qsmt07 <= 1'b0;
  else
    Qsmt07 <= Kg98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ewmt07 <= 1'b0;
  else
    Ewmt07 <= D8a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wzmt07 <= 1'b0;
  else
    Wzmt07 <= Lca8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O3nt07 <= 1'b0;
  else
    O3nt07 <= Tga8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    G7nt07 <= 1'b0;
  else
    G7nt07 <= Bla8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yant07 <= 1'b0;
  else
    Yant07 <= V3a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qent07 <= 1'b0;
  else
    Qent07 <= P6b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cint07 <= 1'b0;
  else
    Cint07 <= Xab8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Olnt07 <= 1'b0;
  else
    Olnt07 <= Ffb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Apnt07 <= 1'b0;
  else
    Apnt07 <= Njb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Msnt07 <= 1'b0;
  else
    Msnt07 <= H2b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yvnt07 <= 1'b0;
  else
    Yvnt07 <= Zxa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kznt07 <= 1'b0;
  else
    Kznt07 <= Rta8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W2ot07 <= 1'b0;
  else
    W2ot07 <= Hb98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    I6ot07 <= 1'b0;
  else
    I6ot07 <= Ld98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U9ot07 <= 1'b0;
  else
    U9ot07 <= Dg98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gdot07 <= 1'b0;
  else
    Gdot07 <= Xj98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sgot07 <= 1'b0;
  else
    Sgot07 <= Pm98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ekot07 <= 1'b0;
  else
    Ekot07 <= Qq98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qnot07 <= 1'b0;
  else
    Qnot07 <= Yu98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Crot07 <= 1'b0;
  else
    Crot07 <= D998v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ouot07 <= 1'b0;
  else
    Ouot07 <= W0a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ayot07 <= 1'b0;
  else
    Ayot07 <= O3a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M1pt07 <= 1'b0;
  else
    M1pt07 <= Uka8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y4pt07 <= 1'b0;
  else
    Y4pt07 <= Mga8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K8pt07 <= 1'b0;
  else
    K8pt07 <= Eca8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wbpt07 <= 1'b0;
  else
    Wbpt07 <= W7a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ifpt07 <= 1'b0;
  else
    Ifpt07 <= Kta8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uipt07 <= 1'b0;
  else
    Uipt07 <= Sxa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gmpt07 <= 1'b0;
  else
    Gmpt07 <= A2b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sppt07 <= 1'b0;
  else
    Sppt07 <= Gjb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dtpt07 <= 1'b0;
  else
    Dtpt07 <= Yeb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pwpt07 <= 1'b0;
  else
    Pwpt07 <= Qab8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B0qt07 <= 1'b0;
  else
    B0qt07 <= I6b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N3qt07 <= 1'b0;
  else
    N3qt07 <= Ewb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y6qt07 <= 1'b0;
  else
    Y6qt07 <= Mtb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jaqt07 <= 1'b0;
  else
    Jaqt07 <= Irb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Udqt07 <= 1'b0;
  else
    Udqt07 <= O8c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Chqt07 <= 1'b0;
  else
    Chqt07 <= K6c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pkqt07 <= 1'b0;
  else
    Pkqt07 <= C2c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Coqt07 <= 1'b0;
  else
    Coqt07 <= Yzb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Prqt07 <= 1'b0;
  else
    Prqt07 <= Lwb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cvqt07 <= 1'b0;
  else
    Cvqt07 <= Uwc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zxqt07 <= 1'b0;
  else
    Zxqt07 <= Tv98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q1rt07 <= 1'b0;
  else
    Q1rt07 <= Lr98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H5rt07 <= 1'b0;
  else
    H5rt07 <= Kn98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y8rt07 <= 1'b0;
  else
    Y8rt07 <= Yg98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mcrt07 <= 1'b0;
  else
    Mcrt07 <= R8a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Egrt07 <= 1'b0;
  else
    Egrt07 <= Zca8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wjrt07 <= 1'b0;
  else
    Wjrt07 <= Hha8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Onrt07 <= 1'b0;
  else
    Onrt07 <= Pla8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Grrt07 <= 1'b0;
  else
    Grrt07 <= J4a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yurt07 <= 1'b0;
  else
    Yurt07 <= D7b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kyrt07 <= 1'b0;
  else
    Kyrt07 <= Lbb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W1st07 <= 1'b0;
  else
    W1st07 <= Tfb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    I5st07 <= 1'b0;
  else
    I5st07 <= Bkb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U8st07 <= 1'b0;
  else
    U8st07 <= V2b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gcst07 <= 1'b0;
  else
    Gcst07 <= Nya8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sfst07 <= 1'b0;
  else
    Sfst07 <= Fua8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ejst07 <= 1'b0;
  else
    Ejst07 <= Ob98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qmst07 <= 1'b0;
  else
    Qmst07 <= Sd98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cqst07 <= 1'b0;
  else
    Cqst07 <= Rg98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Otst07 <= 1'b0;
  else
    Otst07 <= Ek98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Axst07 <= 1'b0;
  else
    Axst07 <= Dn98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M0tt07 <= 1'b0;
  else
    M0tt07 <= Er98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y3tt07 <= 1'b0;
  else
    Y3tt07 <= Mv98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K7tt07 <= 1'b0;
  else
    K7tt07 <= K998v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Watt07 <= 1'b0;
  else
    Watt07 <= D1a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Iett07 <= 1'b0;
  else
    Iett07 <= C4a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uhtt07 <= 1'b0;
  else
    Uhtt07 <= Ila8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gltt07 <= 1'b0;
  else
    Gltt07 <= Aha8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sott07 <= 1'b0;
  else
    Sott07 <= Sca8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Estt07 <= 1'b0;
  else
    Estt07 <= K8a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qvtt07 <= 1'b0;
  else
    Qvtt07 <= Yta8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cztt07 <= 1'b0;
  else
    Cztt07 <= Gya8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O2ut07 <= 1'b0;
  else
    O2ut07 <= O2b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    A6ut07 <= 1'b0;
  else
    A6ut07 <= Ujb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L9ut07 <= 1'b0;
  else
    L9ut07 <= Mfb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xcut07 <= 1'b0;
  else
    Xcut07 <= Ebb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jgut07 <= 1'b0;
  else
    Jgut07 <= W6b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vjut07 <= 1'b0;
  else
    Vjut07 <= Swb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gnut07 <= 1'b0;
  else
    Gnut07 <= Ttb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rqut07 <= 1'b0;
  else
    Rqut07 <= Prb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cuut07 <= 1'b0;
  else
    Cuut07 <= V8c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kxut07 <= 1'b0;
  else
    Kxut07 <= R6c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X0vt07 <= 1'b0;
  else
    X0vt07 <= J2c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K4vt07 <= 1'b0;
  else
    K4vt07 <= F0c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X7vt07 <= 1'b0;
  else
    X7vt07 <= Zwb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kbvt07 <= 1'b0;
  else
    Kbvt07 <= Bxc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hevt07 <= 1'b0;
  else
    Hevt07 <= Ru98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yhvt07 <= 1'b0;
  else
    Yhvt07 <= Jq98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Plvt07 <= 1'b0;
  else
    Plvt07 <= Im98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gpvt07 <= 1'b0;
  else
    Gpvt07 <= Wf98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Usvt07 <= 1'b0;
  else
    Usvt07 <= P7a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mwvt07 <= 1'b0;
  else
    Mwvt07 <= Xba8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    E0wt07 <= 1'b0;
  else
    E0wt07 <= Fga8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W3wt07 <= 1'b0;
  else
    W3wt07 <= Nka8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O7wt07 <= 1'b0;
  else
    O7wt07 <= H3a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gbwt07 <= 1'b0;
  else
    Gbwt07 <= B6b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sewt07 <= 1'b0;
  else
    Sewt07 <= Jab8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Eiwt07 <= 1'b0;
  else
    Eiwt07 <= Reb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qlwt07 <= 1'b0;
  else
    Qlwt07 <= Zib8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cpwt07 <= 1'b0;
  else
    Cpwt07 <= T1b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oswt07 <= 1'b0;
  else
    Oswt07 <= Lxa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Awwt07 <= 1'b0;
  else
    Awwt07 <= Dta8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mzwt07 <= 1'b0;
  else
    Mzwt07 <= Ab98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y2xt07 <= 1'b0;
  else
    Y2xt07 <= Ed98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K6xt07 <= 1'b0;
  else
    K6xt07 <= Pf98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W9xt07 <= 1'b0;
  else
    W9xt07 <= Qj98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Idxt07 <= 1'b0;
  else
    Idxt07 <= Bm98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ugxt07 <= 1'b0;
  else
    Ugxt07 <= Cq98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gkxt07 <= 1'b0;
  else
    Gkxt07 <= Ku98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Snxt07 <= 1'b0;
  else
    Snxt07 <= W898v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Erxt07 <= 1'b0;
  else
    Erxt07 <= P0a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Quxt07 <= 1'b0;
  else
    Quxt07 <= A3a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cyxt07 <= 1'b0;
  else
    Cyxt07 <= Gka8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O1yt07 <= 1'b0;
  else
    O1yt07 <= Yfa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    A5yt07 <= 1'b0;
  else
    A5yt07 <= Qba8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M8yt07 <= 1'b0;
  else
    M8yt07 <= I7a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ybyt07 <= 1'b0;
  else
    Ybyt07 <= Wsa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kfyt07 <= 1'b0;
  else
    Kfyt07 <= Exa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wiyt07 <= 1'b0;
  else
    Wiyt07 <= M1b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Imyt07 <= 1'b0;
  else
    Imyt07 <= Sib8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tpyt07 <= 1'b0;
  else
    Tpyt07 <= Keb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ftyt07 <= 1'b0;
  else
    Ftyt07 <= Cab8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rwyt07 <= 1'b0;
  else
    Rwyt07 <= U5b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D0zt07 <= 1'b0;
  else
    D0zt07 <= Qvb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O3zt07 <= 1'b0;
  else
    O3zt07 <= Ftb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z6zt07 <= 1'b0;
  else
    Z6zt07 <= Brb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kazt07 <= 1'b0;
  else
    Kazt07 <= H8c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sdzt07 <= 1'b0;
  else
    Sdzt07 <= D6c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fhzt07 <= 1'b0;
  else
    Fhzt07 <= V1c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Skzt07 <= 1'b0;
  else
    Skzt07 <= Xvb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fozt07 <= 1'b0;
  else
    Fozt07 <= Ixc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Crzt07 <= 1'b0;
  else
    Crzt07 <= Du98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tuzt07 <= 1'b0;
  else
    Tuzt07 <= Vp98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kyzt07 <= 1'b0;
  else
    Kyzt07 <= Ul98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B20u07 <= 1'b0;
  else
    B20u07 <= If98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P50u07 <= 1'b0;
  else
    P50u07 <= Zja8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H90u07 <= 1'b0;
  else
    H90u07 <= Rfa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zc0u07 <= 1'b0;
  else
    Zc0u07 <= Jba8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rg0u07 <= 1'b0;
  else
    Rg0u07 <= B7a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jk0u07 <= 1'b0;
  else
    Jk0u07 <= T2a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bo0u07 <= 1'b0;
  else
    Bo0u07 <= N5b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nr0u07 <= 1'b0;
  else
    Nr0u07 <= V9b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zu0u07 <= 1'b0;
  else
    Zu0u07 <= Deb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ly0u07 <= 1'b0;
  else
    Ly0u07 <= Lib8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X11u07 <= 1'b0;
  else
    X11u07 <= F1b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J51u07 <= 1'b0;
  else
    J51u07 <= Xwa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V81u07 <= 1'b0;
  else
    V81u07 <= Psa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hc1u07 <= 1'b0;
  else
    Hc1u07 <= A8c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pf1u07 <= 1'b0;
  else
    Pf1u07 <= W5c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cj1u07 <= 1'b0;
  else
    Cj1u07 <= O1c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pm1u07 <= 1'b0;
  else
    Pm1u07 <= Jvb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cq1u07 <= 1'b0;
  else
    Cq1u07 <= I0a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ot1u07 <= 1'b0;
  else
    Ot1u07 <= M2a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ax1u07 <= 1'b0;
  else
    Ax1u07 <= Sja8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M02u07 <= 1'b0;
  else
    M02u07 <= Cba8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y32u07 <= 1'b0;
  else
    Y32u07 <= U6a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K72u07 <= 1'b0;
  else
    K72u07 <= Isa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wa2u07 <= 1'b0;
  else
    Wa2u07 <= Qwa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ie2u07 <= 1'b0;
  else
    Ie2u07 <= Y0b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uh2u07 <= 1'b0;
  else
    Uh2u07 <= Eib8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fl2u07 <= 1'b0;
  else
    Fl2u07 <= Wdb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ro2u07 <= 1'b0;
  else
    Ro2u07 <= O9b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ds2u07 <= 1'b0;
  else
    Ds2u07 <= G5b8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pv2u07 <= 1'b0;
  else
    Pv2u07 <= Cvb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Az2u07 <= 1'b0;
  else
    Az2u07 <= Ysb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L23u07 <= 1'b0;
  else
    L23u07 <= Uqb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W53u07 <= 1'b0;
  else
    W53u07 <= Ta98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    I93u07 <= 1'b0;
  else
    I93u07 <= Xc98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uc3u07 <= 1'b0;
  else
    Uc3u07 <= Bf98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gg3u07 <= 1'b0;
  else
    Gg3u07 <= Jj98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sj3u07 <= 1'b0;
  else
    Sj3u07 <= Nl98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    En3u07 <= 1'b0;
  else
    En3u07 <= Wt98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qq3u07 <= 1'b0;
  else
    Qq3u07 <= Q8k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cu3u07 <= 1'b0;
  else
    Cu3u07 <= P898v6;

always @(posedge HCLK) Ox3u07 <= Nbc8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oz3u07 <= 1'b0;
  else
    Oz3u07 <= P5c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B34u07 <= 1'b0;
  else
    B34u07 <= I5c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O64u07 <= 1'b0;
  else
    O64u07 <= B5c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ba4u07 <= 1'b0;
  else
    Ba4u07 <= U4c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Od4u07 <= 1'b0;
  else
    Od4u07 <= N4c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bh4u07 <= 1'b0;
  else
    Bh4u07 <= G4c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ok4u07 <= 1'b0;
  else
    Ok4u07 <= Z3c8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bo4u07 <= 1'b0;
  else
    Bo4u07 <= S3c8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Or4u07 <= 1'b0;
  else
    Or4u07 <= Vk78v6;

always @(posedge HCLK) Lt4u07 <= H768v6;
always @(posedge HCLK) Av4u07 <= Fz58v6;
always @(posedge HCLK) Pw4u07 <= Dr58v6;
always @(posedge HCLK) Ey4u07 <= Bj58v6;
always @(posedge HCLK) Tz4u07 <= Za58v6;
always @(posedge HCLK) I15u07 <= X258v6;
always @(posedge HCLK) X25u07 <= Jv48v6;
always @(posedge HCLK) M45u07 <= Vn48v6;
always @(posedge FCLK) B65u07 <= Xjv7v6;
always @(posedge FCLK) H85u07 <= Thv7v6;
always @(posedge HCLK) Na5u07 <= Zoy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uc5u07 <= 1'b0;
  else
    Uc5u07 <= Xmk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ef5u07 <= 1'b0;
  else
    Ef5u07 <= R5s7v6;

always @(posedge HCLK) Ii5u07 <= Soy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pk5u07 <= 1'b0;
  else
    Pk5u07 <= I3l8v6;

always @(posedge HCLK) Zm5u07 <= Dky7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xp5u07 <= 1'b0;
  else
    Xp5u07 <= K5s7v6;

always @(posedge HCLK) Bt5u07 <= Loy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Iv5u07 <= 1'b0;
  else
    Iv5u07 <= Hzk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sx5u07 <= 1'b0;
  else
    Sx5u07 <= D5s7v6;

always @(posedge HCLK) W06u07 <= Eoy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D36u07 <= 1'b0;
  else
    D36u07 <= K1p7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    I66u07 <= 1'b0;
  else
    I66u07 <= Nzo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N96u07 <= 1'b0;
  else
    N96u07 <= Syo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tc6u07 <= 1'b0;
  else
    Tc6u07 <= Lyo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zf6u07 <= 1'b0;
  else
    Zf6u07 <= Eyo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fj6u07 <= 1'b0;
  else
    Fj6u07 <= Xxo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lm6u07 <= 1'b0;
  else
    Lm6u07 <= Jxo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rp6u07 <= 1'b0;
  else
    Rp6u07 <= Hwo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xs6u07 <= 1'b0;
  else
    Xs6u07 <= Fvo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dw6u07 <= 1'b0;
  else
    Dw6u07 <= Yuo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jz6u07 <= 1'b0;
  else
    Jz6u07 <= Ruo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P27u07 <= 1'b0;
  else
    P27u07 <= Kuo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V57u07 <= 1'b0;
  else
    V57u07 <= Duo7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B97u07 <= 1'b0;
  else
    B97u07 <= W4s7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fc7u07 <= 1'b0;
  else
    Fc7u07 <= Lqw7v6;

always @(posedge FCLK) Fe7u07 <= Eqi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qg7u07 <= 1'b0;
  else
    Qg7u07 <= Jiw7v6;

always @(posedge FCLK) Qi7u07 <= Xpi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bl7u07 <= 1'b0;
  else
    Bl7u07 <= Qiw7v6;

always @(posedge FCLK) Bn7u07 <= Qpi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mp7u07 <= 1'b0;
  else
    Mp7u07 <= Xiw7v6;

always @(posedge FCLK) Mr7u07 <= Jpi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xt7u07 <= 1'b0;
  else
    Xt7u07 <= Ejw7v6;

always @(posedge FCLK) Xv7u07 <= Cpi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Iy7u07 <= 1'b0;
  else
    Iy7u07 <= Ljw7v6;

always @(posedge FCLK) I08u07 <= Voi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T28u07 <= 1'b0;
  else
    T28u07 <= Sjw7v6;

always @(posedge FCLK) T48u07 <= Ooi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    E78u07 <= 1'b0;
  else
    E78u07 <= Zjw7v6;

always @(posedge FCLK) E98u07 <= Hoi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pb8u07 <= 1'b0;
  else
    Pb8u07 <= Gkw7v6;

always @(posedge FCLK) Pd8u07 <= Aoi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ag8u07 <= 1'b0;
  else
    Ag8u07 <= Nkw7v6;

always @(posedge FCLK) Bi8u07 <= Tni7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nk8u07 <= 1'b0;
  else
    Nk8u07 <= Ukw7v6;

always @(posedge FCLK) Om8u07 <= Mni7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ap8u07 <= 1'b0;
  else
    Ap8u07 <= Blw7v6;

always @(posedge FCLK) Br8u07 <= Fni7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nt8u07 <= 1'b0;
  else
    Nt8u07 <= Ilw7v6;

always @(posedge FCLK) Ov8u07 <= Ymi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ay8u07 <= 1'b0;
  else
    Ay8u07 <= Plw7v6;

always @(posedge FCLK) B09u07 <= Rmi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N29u07 <= 1'b0;
  else
    N29u07 <= Wlw7v6;

always @(posedge FCLK) O49u07 <= Kmi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    A79u07 <= 1'b0;
  else
    A79u07 <= Dmw7v6;

always @(posedge FCLK) B99u07 <= Dmi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nb9u07 <= 1'b0;
  else
    Nb9u07 <= Kmw7v6;

always @(posedge FCLK) Od9u07 <= Wli7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ag9u07 <= 1'b0;
  else
    Ag9u07 <= Rmw7v6;

always @(posedge FCLK) Bi9u07 <= Pli7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nk9u07 <= 1'b0;
  else
    Nk9u07 <= Ymw7v6;

always @(posedge FCLK) Om9u07 <= Ili7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ap9u07 <= 1'b0;
  else
    Ap9u07 <= Fnw7v6;

always @(posedge FCLK) Br9u07 <= Bli7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nt9u07 <= 1'b0;
  else
    Nt9u07 <= Mnw7v6;

always @(posedge FCLK) Ov9u07 <= Uki7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ay9u07 <= 1'b0;
  else
    Ay9u07 <= Tnw7v6;

always @(posedge FCLK) B0au07 <= Nki7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N2au07 <= 1'b0;
  else
    N2au07 <= Aow7v6;

always @(posedge FCLK) O4au07 <= Gki7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    A7au07 <= 1'b0;
  else
    A7au07 <= How7v6;

always @(posedge FCLK) B9au07 <= Zji7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nbau07 <= 1'b0;
  else
    Nbau07 <= Oow7v6;

always @(posedge FCLK) Odau07 <= Sji7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Agau07 <= 1'b0;
  else
    Agau07 <= Vow7v6;

always @(posedge FCLK) Biau07 <= Lji7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nkau07 <= 1'b0;
  else
    Nkau07 <= Cpw7v6;

always @(posedge FCLK) Omau07 <= Eji7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Apau07 <= 1'b0;
  else
    Apau07 <= Jpw7v6;

always @(posedge FCLK) Brau07 <= Xii7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ntau07 <= 1'b0;
  else
    Ntau07 <= Qpw7v6;

always @(posedge FCLK) Ovau07 <= Qii7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ayau07 <= 1'b0;
  else
    Ayau07 <= Xpw7v6;

always @(posedge FCLK) B0bu07 <= Jii7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N2bu07 <= 1'b0;
  else
    N2bu07 <= Eqw7v6;

always @(posedge FCLK) O4bu07 <= Cii7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    A7bu07 <= 1'b0;
  else
    A7bu07 <= I7zmz6[31];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    A9bu07 <= 1'b0;
  else
    A9bu07 <= I7zmz6[1];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zabu07 <= 1'b0;
  else
    Zabu07 <= L5zmz6[1];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ldbu07 <= 1'b0;
  else
    Ldbu07 <= L5zmz6[1];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Sfbu07 <= 1'b0;
  else
    Sfbu07 <= I7zmz6[2];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rhbu07 <= 1'b0;
  else
    Rhbu07 <= L5zmz6[2];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dkbu07 <= 1'b0;
  else
    Dkbu07 <= L5zmz6[2];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kmbu07 <= 1'b0;
  else
    Kmbu07 <= I7zmz6[3];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jobu07 <= 1'b0;
  else
    Jobu07 <= L5zmz6[3];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vqbu07 <= 1'b0;
  else
    Vqbu07 <= L5zmz6[3];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ctbu07 <= 1'b0;
  else
    Ctbu07 <= I7zmz6[4];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bvbu07 <= 1'b0;
  else
    Bvbu07 <= L5zmz6[4];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Nxbu07 <= 1'b0;
  else
    Nxbu07 <= L5zmz6[4];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Uzbu07 <= 1'b0;
  else
    Uzbu07 <= I7zmz6[5];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    T1cu07 <= 1'b0;
  else
    T1cu07 <= L5zmz6[5];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F4cu07 <= 1'b0;
  else
    F4cu07 <= L5zmz6[5];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    M6cu07 <= 1'b0;
  else
    M6cu07 <= I7zmz6[6];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    L8cu07 <= 1'b0;
  else
    L8cu07 <= L5zmz6[6];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xacu07 <= 1'b0;
  else
    Xacu07 <= L5zmz6[6];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Edcu07 <= 1'b0;
  else
    Edcu07 <= I7zmz6[7];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dfcu07 <= 1'b0;
  else
    Dfcu07 <= L5zmz6[7];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Phcu07 <= 1'b0;
  else
    Phcu07 <= I7zmz6[8];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ojcu07 <= 1'b0;
  else
    Ojcu07 <= L5zmz6[8];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Amcu07 <= 1'b0;
  else
    Amcu07 <= I7zmz6[9];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zncu07 <= 1'b0;
  else
    Zncu07 <= L5zmz6[9];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lqcu07 <= 1'b0;
  else
    Lqcu07 <= I7zmz6[10];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lscu07 <= 1'b0;
  else
    Lscu07 <= L5zmz6[10];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yucu07 <= 1'b0;
  else
    Yucu07 <= I7zmz6[11];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ywcu07 <= 1'b0;
  else
    Ywcu07 <= L5zmz6[11];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lzcu07 <= 1'b0;
  else
    Lzcu07 <= I7zmz6[12];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    L1du07 <= 1'b0;
  else
    L1du07 <= L5zmz6[12];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Y3du07 <= 1'b0;
  else
    Y3du07 <= I7zmz6[13];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Y5du07 <= 1'b0;
  else
    Y5du07 <= L5zmz6[13];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    L8du07 <= 1'b0;
  else
    L8du07 <= I7zmz6[14];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ladu07 <= 1'b0;
  else
    Ladu07 <= L5zmz6[14];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ycdu07 <= 1'b0;
  else
    Ycdu07 <= I7zmz6[15];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yedu07 <= 1'b0;
  else
    Yedu07 <= L5zmz6[15];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lhdu07 <= 1'b0;
  else
    Lhdu07 <= I7zmz6[16];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ljdu07 <= 1'b0;
  else
    Ljdu07 <= L5zmz6[16];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yldu07 <= 1'b0;
  else
    Yldu07 <= I7zmz6[17];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yndu07 <= 1'b0;
  else
    Yndu07 <= L5zmz6[17];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lqdu07 <= 1'b0;
  else
    Lqdu07 <= I7zmz6[18];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lsdu07 <= 1'b0;
  else
    Lsdu07 <= L5zmz6[18];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yudu07 <= 1'b0;
  else
    Yudu07 <= I7zmz6[19];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ywdu07 <= 1'b0;
  else
    Ywdu07 <= L5zmz6[19];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lzdu07 <= 1'b0;
  else
    Lzdu07 <= I7zmz6[20];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    L1eu07 <= 1'b0;
  else
    L1eu07 <= Tct8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Y3eu07 <= 1'b0;
  else
    Y3eu07 <= I7zmz6[21];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Y5eu07 <= 1'b0;
  else
    Y5eu07 <= L5zmz6[21];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    L8eu07 <= 1'b0;
  else
    L8eu07 <= I7zmz6[22];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Laeu07 <= 1'b0;
  else
    Laeu07 <= L5zmz6[22];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yceu07 <= 1'b0;
  else
    Yceu07 <= I7zmz6[23];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yeeu07 <= 1'b0;
  else
    Yeeu07 <= L5zmz6[23];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lheu07 <= 1'b0;
  else
    Lheu07 <= I7zmz6[24];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ljeu07 <= 1'b0;
  else
    Ljeu07 <= L5zmz6[24];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yleu07 <= 1'b0;
  else
    Yleu07 <= I7zmz6[25];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yneu07 <= 1'b0;
  else
    Yneu07 <= L5zmz6[25];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lqeu07 <= 1'b0;
  else
    Lqeu07 <= I7zmz6[26];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lseu07 <= 1'b0;
  else
    Lseu07 <= L5zmz6[26];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yueu07 <= 1'b0;
  else
    Yueu07 <= I7zmz6[27];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yweu07 <= 1'b0;
  else
    Yweu07 <= L5zmz6[27];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lzeu07 <= 1'b0;
  else
    Lzeu07 <= I7zmz6[28];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    L1fu07 <= 1'b0;
  else
    L1fu07 <= L5zmz6[28];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Y3fu07 <= 1'b0;
  else
    Y3fu07 <= I7zmz6[29];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Y5fu07 <= 1'b0;
  else
    Y5fu07 <= L5zmz6[29];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    L8fu07 <= 1'b0;
  else
    L8fu07 <= I7zmz6[30];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lafu07 <= 1'b0;
  else
    Lafu07 <= L5zmz6[30];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ycfu07 <= 1'b0;
  else
    Ycfu07 <= L5zmz6[31];

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lffu07 <= 1'b0;
  else
    Lffu07 <= Ipk8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mhfu07 <= 1'b0;
  else
    Mhfu07 <= Bmv7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ljfu07 <= 1'b0;
  else
    Ljfu07 <= Fb88v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rlfu07 <= 1'b0;
  else
    Rlfu07 <= Mb88v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rnfu07 <= 1'b0;
  else
    Rnfu07 <= P988v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zpfu07 <= 1'b0;
  else
    Zpfu07 <= Pew7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bsfu07 <= 1'b0;
  else
    Bsfu07 <= Mgw7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cufu07 <= 1'b0;
  else
    Cufu07 <= Ciw7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dwfu07 <= 1'b0;
  else
    Dwfu07 <= Fgw7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Eyfu07 <= 1'b0;
  else
    Eyfu07 <= J4w7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    D0gu07 <= 1'b0;
  else
    D0gu07 <= Yfw7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    D2gu07 <= 1'b0;
  else
    D2gu07 <= Rfw7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    L4gu07 <= 1'b0;
  else
    L4gu07 <= Wew7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    N6gu07 <= 1'b0;
  else
    N6gu07 <= Vhi7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O9gu07 <= 1'b0;
  else
    O9gu07 <= Zb48v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pbgu07 <= 1'b0;
  else
    Pbgu07 <= Bcy7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ndgu07 <= 1'b0;
  else
    Ndgu07 <= Uby7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ofgu07 <= 1'b0;
  else
    Ofgu07 <= Rka7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Uhgu07 <= 1'b0;
  else
    Uhgu07 <= W3a7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Akgu07 <= 1'b0;
  else
    Akgu07 <= T6k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Imgu07 <= 1'b0;
  else
    Imgu07 <= M6k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qogu07 <= 1'b0;
  else
    Qogu07 <= Ohi7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Uqgu07 <= 1'b0;
  else
    Uqgu07 <= Hhi7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xsgu07 <= 1'b0;
  else
    Xsgu07 <= Ahi7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wugu07 <= 1'b0;
  else
    Wugu07 <= Tgi7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vwgu07 <= 1'b0;
  else
    Vwgu07 <= Cy97v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Azgu07 <= 1'b0;
  else
    Azgu07 <= Edo7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    D1hu07 <= 1'b0;
  else
    D1hu07 <= P7b7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    E3hu07 <= 1'b0;
  else
    E3hu07 <= Vca7v6;

always @(posedge HCLK) H5hu07 <= Aqu7v6;
always @(posedge HCLK) K7hu07 <= Tpu7v6;
always @(posedge HCLK) N9hu07 <= Mpu7v6;
always @(posedge HCLK) Rbhu07 <= Fpu7v6;
always @(posedge HCLK) Vdhu07 <= You7v6;
always @(posedge HCLK) Zfhu07 <= Rou7v6;
always @(posedge HCLK) Dihu07 <= Kou7v6;
always @(posedge HCLK) Hkhu07 <= Dou7v6;
always @(posedge HCLK) Lmhu07 <= Wnu7v6;
always @(posedge HCLK) Pohu07 <= Pnu7v6;
always @(posedge HCLK) Tqhu07 <= Inu7v6;
always @(posedge HCLK) Xshu07 <= Bnu7v6;
always @(posedge HCLK) Bvhu07 <= Umu7v6;
always @(posedge HCLK) Fxhu07 <= Nmu7v6;
always @(posedge HCLK) Jzhu07 <= Gmu7v6;
always @(posedge HCLK) N1iu07 <= Zlu7v6;
always @(posedge HCLK) R3iu07 <= Slu7v6;
always @(posedge HCLK) V5iu07 <= Llu7v6;
always @(posedge HCLK) Z7iu07 <= Elu7v6;
always @(posedge HCLK) Daiu07 <= Xku7v6;
always @(posedge HCLK) Hciu07 <= Qku7v6;
always @(posedge HCLK) Leiu07 <= Jku7v6;
always @(posedge HCLK) Pgiu07 <= Cku7v6;
always @(posedge HCLK) Tiiu07 <= Vju7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xkiu07 <= 1'b0;
  else
    Xkiu07 <= T1zmz6[15];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fniu07 <= 1'b0;
  else
    Fniu07 <= T1zmz6[23];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Npiu07 <= 1'b0;
  else
    Npiu07 <= T1zmz6[31];

always @(posedge HCLK) Vriu07 <= Oju7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ytiu07 <= 1'b0;
  else
    Ytiu07 <= T1zmz6[10];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gwiu07 <= 1'b0;
  else
    Gwiu07 <= T1zmz6[11];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Oyiu07 <= 1'b0;
  else
    Oyiu07 <= T1zmz6[12];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    W0ju07 <= 1'b0;
  else
    W0ju07 <= T1zmz6[13];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    E3ju07 <= 1'b0;
  else
    E3ju07 <= T1zmz6[16];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    M5ju07 <= 1'b0;
  else
    M5ju07 <= T1zmz6[17];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    U7ju07 <= 1'b0;
  else
    U7ju07 <= T1zmz6[18];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Caju07 <= 1'b0;
  else
    Caju07 <= T1zmz6[19];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kcju07 <= 1'b0;
  else
    Kcju07 <= T1zmz6[20];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Seju07 <= 1'b0;
  else
    Seju07 <= T1zmz6[21];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ahju07 <= 1'b0;
  else
    Ahju07 <= T1zmz6[24];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ijju07 <= 1'b0;
  else
    Ijju07 <= T1zmz6[25];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qlju07 <= 1'b0;
  else
    Qlju07 <= T1zmz6[26];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ynju07 <= 1'b0;
  else
    Ynju07 <= T1zmz6[27];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gqju07 <= 1'b0;
  else
    Gqju07 <= T1zmz6[28];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Osju07 <= 1'b0;
  else
    Osju07 <= T1zmz6[29];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wuju07 <= 1'b0;
  else
    Wuju07 <= T1zmz6[34];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Exju07 <= 1'b0;
  else
    Exju07 <= T1zmz6[35];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mzju07 <= 1'b0;
  else
    Mzju07 <= T1zmz6[8];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    T1ku07 <= 1'b0;
  else
    T1ku07 <= T1zmz6[9];

always @(posedge HCLK) A4ku07 <= Mgi7v6;
always @(posedge HCLK) J6ku07 <= Fgi7v6;
always @(posedge HCLK) A9ku07 <= Yfi7v6;
always @(posedge HCLK) Ibku07 <= Gtu7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gdku07 <= 1'b0;
  else
    Gdku07 <= Hsk8v6;

always @(posedge HCLK) Afku07 <= Rvu7v6;
always @(posedge HCLK) Zgku07 <= Kvu7v6;
always @(posedge HCLK) Xiku07 <= Dvu7v6;
always @(posedge HCLK) Vkku07 <= Wuu7v6;
always @(posedge HCLK) Tmku07 <= Puu7v6;
always @(posedge HCLK) Roku07 <= Iuu7v6;
always @(posedge HCLK) Pqku07 <= Buu7v6;
always @(posedge HCLK) Nsku07 <= Utu7v6;
always @(posedge HCLK) Luku07 <= Ntu7v6;
always @(posedge HCLK) Jwku07 <= Zsu7v6;
always @(posedge HCLK) Hyku07 <= Ssu7v6;
always @(posedge HCLK) G0lu07 <= Lsu7v6;
always @(posedge HCLK) F2lu07 <= Esu7v6;
always @(posedge HCLK) E4lu07 <= Xru7v6;
always @(posedge HCLK) D6lu07 <= Qru7v6;
always @(posedge HCLK) C8lu07 <= Rfi7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ualu07 <= 1'b0;
  else
    Ualu07 <= Mec8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qclu07 <= 1'b0;
  else
    Qclu07 <= H8y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pelu07 <= 1'b0;
  else
    Pelu07 <= I5y7v6;

always @(posedge HCLK) Qglu07 <= Iid8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qilu07 <= 1'b0;
  else
    Qilu07 <= Xfd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tklu07 <= 1'b0;
  else
    Tklu07 <= Egd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vmlu07 <= 1'b0;
  else
    Vmlu07 <= Nqb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hqlu07 <= 1'b0;
  else
    Hqlu07 <= Gqb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Stlu07 <= 1'b0;
  else
    Stlu07 <= Zpb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Exlu07 <= 1'b0;
  else
    Exlu07 <= Spb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P0mu07 <= 1'b0;
  else
    P0mu07 <= Lpb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B4mu07 <= 1'b0;
  else
    B4mu07 <= Epb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M7mu07 <= 1'b0;
  else
    M7mu07 <= Xob8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yamu07 <= 1'b0;
  else
    Yamu07 <= Qob8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jemu07 <= 1'b0;
  else
    Jemu07 <= Job8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vhmu07 <= 1'b0;
  else
    Vhmu07 <= Cob8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Glmu07 <= 1'b0;
  else
    Glmu07 <= Vnb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Somu07 <= 1'b0;
  else
    Somu07 <= Onb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dsmu07 <= 1'b0;
  else
    Dsmu07 <= Hnb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pvmu07 <= 1'b0;
  else
    Pvmu07 <= Anb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Azmu07 <= 1'b0;
  else
    Azmu07 <= Tmb8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M2nu07 <= 1'b0;
  else
    M2nu07 <= Mmb8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    X5nu07 <= 1'b0;
  else
    X5nu07 <= Lm78v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    U7nu07 <= 1'b0;
  else
    U7nu07 <= Jt68v6;

always @(posedge HCLK) W9nu07 <= Tk68v6;
always @(posedge HCLK) Mbnu07 <= Md68v6;
always @(posedge HCLK) Bdnu07 <= K568v6;
always @(posedge HCLK) Qenu07 <= Ix58v6;
always @(posedge HCLK) Fgnu07 <= Gp58v6;
always @(posedge HCLK) Uhnu07 <= Eh58v6;
always @(posedge HCLK) Jjnu07 <= C958v6;
always @(posedge HCLK) Yknu07 <= A158v6;
always @(posedge HCLK) Nmnu07 <= Mt48v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Conu07 <= 1'b0;
  else
    Conu07 <= Uas7v6;

always @(posedge HCLK) Frnu07 <= Uz28v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wtnu07 <= 1'b0;
  else
    Wtnu07 <= Bbs7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ee9917 <= 1'b0;
  else
    Ee9917 <= Ixy7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ng9917 <= 1'b0;
  else
    Ng9917 <= B0p7v6;

always @(posedge HCLK) Sj9917 <= Nz28v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jm9917 <= 1'b0;
  else
    Jm9917 <= Ibs7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mp9917 <= 1'b0;
  else
    Mp9917 <= Fzy7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vr9917 <= 1'b0;
  else
    Vr9917 <= I0p7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Av9917 <= 1'b0;
  else
    Av9917 <= Vlk8v6;

always @(posedge HCLK) Ix9917 <= Zy28v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zz9917 <= 1'b0;
  else
    Zz9917 <= Pbk8v6;

always @(posedge HCLK) I2a917 <= Sy28v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z4a917 <= 1'b0;
  else
    Z4a917 <= Dcs7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    C8a917 <= 1'b0;
  else
    C8a917 <= J1z7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Laa917 <= 1'b0;
  else
    Laa917 <= Juc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hda917 <= 1'b0;
  else
    Hda917 <= Vtc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dga917 <= 1'b0;
  else
    Dga917 <= Htc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zia917 <= 1'b0;
  else
    Zia917 <= Atc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vla917 <= 1'b0;
  else
    Vla917 <= Tsc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Roa917 <= 1'b0;
  else
    Roa917 <= Fsc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nra917 <= 1'b0;
  else
    Nra917 <= Kfi7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mta917 <= 1'b0;
  else
    Mta917 <= Dfi7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mva917 <= 1'b0;
  else
    Mva917 <= Wei7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rxa917 <= 1'b0;
  else
    Rxa917 <= Jnc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vza917 <= 1'b0;
  else
    Vza917 <= Rrc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y1b917 <= 1'b0;
  else
    Y1b917 <= Ykc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    W3b917 <= 1'b0;
  else
    W3b917 <= Pei7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    X6b917 <= 1'b0;
  else
    X6b917 <= Flc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    A9b917 <= 1'b0;
  else
    A9b917 <= Krc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dbb917 <= 1'b0;
  else
    Dbb917 <= Drc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gdb917 <= 1'b0;
  else
    Gdb917 <= Wqc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jfb917 <= 1'b0;
  else
    Jfb917 <= Pqc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mhb917 <= 1'b0;
  else
    Mhb917 <= Iqc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pjb917 <= 1'b0;
  else
    Pjb917 <= Bqc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Slb917 <= 1'b0;
  else
    Slb917 <= Upc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vnb917 <= 1'b0;
  else
    Vnb917 <= Npc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ypb917 <= 1'b0;
  else
    Ypb917 <= Gpc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bsb917 <= 1'b0;
  else
    Bsb917 <= Zoc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fub917 <= 1'b0;
  else
    Fub917 <= Soc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jwb917 <= 1'b0;
  else
    Jwb917 <= Loc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nyb917 <= 1'b0;
  else
    Nyb917 <= Eoc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    R0c917 <= 1'b0;
  else
    R0c917 <= Xnc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    V2c917 <= 1'b0;
  else
    V2c917 <= Qnc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z4c917 <= 1'b0;
  else
    Z4c917 <= Cnc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    D7c917 <= 1'b0;
  else
    D7c917 <= Vmc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    H9c917 <= 1'b0;
  else
    H9c917 <= Omc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lbc917 <= 1'b0;
  else
    Lbc917 <= Hmc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pdc917 <= 1'b0;
  else
    Pdc917 <= Amc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tfc917 <= 1'b0;
  else
    Tfc917 <= Tlc8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xhc917 <= 1'b0;
  else
    Xhc917 <= Mlc8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bkc917 <= 1'b0;
  else
    Bkc917 <= Iei7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Slc917 <= 1'b0;
  else
    Slc917 <= Bei7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rnc917 <= 1'b0;
  else
    Rnc917 <= Udi7v6;

always @(posedge HCLK) Mpc917 <= Ndi7v6;
always @(posedge HCLK) Vrc917 <= Gdi7v6;
always @(posedge HCLK) Muc917 <= Zci7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Uwc917 <= 1'b0;
  else
    Uwc917 <= Ty77v6;

always @(posedge HCLK) Vyc917 <= Sci7v6;
always @(posedge HCLK) N1d917 <= Lci7v6;
always @(posedge HCLK) C4d917 <= Eci7v6;
always @(posedge HCLK) R6d917 <= Xbi7v6;
always @(posedge HCLK) G9d917 <= Qbi7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vbd917 <= 1'b1;
  else
    Vbd917 <= Zu68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ydd917 <= 1'b0;
  else
    Ydd917 <= N548v6;

always @(posedge FCLK) Dgd917 <= Jbi7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Nid917 <= 1'b0;
  else
    Nid917 <= Vgx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rkd917 <= 1'b0;
  else
    Rkd917 <= U548v6;

always @(posedge FCLK) Wmd917 <= Cbi7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gpd917 <= 1'b0;
  else
    Gpd917 <= Yex7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Krd917 <= 1'b0;
  else
    Krd917 <= Zxymz6[7];

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rtd917 <= 1'b0;
  else
    Rtd917 <= B648v6;

always @(posedge FCLK) Wvd917 <= Vai7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gyd917 <= 1'b0;
  else
    Gyd917 <= Ffx7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    K0e917 <= 1'b0;
  else
    K0e917 <= Zxymz6[6];

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R2e917 <= 1'b0;
  else
    R2e917 <= I648v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W4e917 <= 1'b0;
  else
    W4e917 <= Y048v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    V7e917 <= 1'b0;
  else
    V7e917 <= R048v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uae917 <= 1'b0;
  else
    Uae917 <= G548v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sde917 <= 1'b0;
  else
    Sde917 <= Z448v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qge917 <= 1'b0;
  else
    Qge917 <= C348v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pje917 <= 1'b0;
  else
    Pje917 <= V248v6;

always @(posedge FCLK) Ome917 <= Oai7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yoe917 <= 1'b0;
  else
    Yoe917 <= Mfx7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cre917 <= 1'b0;
  else
    Cre917 <= Zxymz6[5];

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jte917 <= 1'b0;
  else
    Jte917 <= W648v6;

always @(posedge FCLK) Ove917 <= Hai7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yxe917 <= 1'b0;
  else
    Yxe917 <= Agx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    C0f917 <= 1'b0;
  else
    C0f917 <= K748v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H2f917 <= 1'b0;
  else
    H2f917 <= A2x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    G5f917 <= 1'b0;
  else
    G5f917 <= T1x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F8f917 <= 1'b0;
  else
    F8f917 <= I6x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ebf917 <= 1'b0;
  else
    Ebf917 <= B6x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Def917 <= 1'b0;
  else
    Def917 <= Qax7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Chf917 <= 1'b0;
  else
    Chf917 <= Jax7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bkf917 <= 1'b0;
  else
    Bkf917 <= Dex7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zmf917 <= 1'b0;
  else
    Zmf917 <= O0d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wof917 <= 1'b0;
  else
    Wof917 <= Ws38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vrf917 <= 1'b0;
  else
    Vrf917 <= Ps38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uuf917 <= 1'b0;
  else
    Uuf917 <= Av38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Txf917 <= 1'b0;
  else
    Txf917 <= Tu38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    S0g917 <= 1'b0;
  else
    S0g917 <= Ex38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    R3g917 <= 1'b0;
  else
    R3g917 <= Xw38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q6g917 <= 1'b0;
  else
    Q6g917 <= O2x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    P9g917 <= 1'b0;
  else
    P9g917 <= H2x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ocg917 <= 1'b0;
  else
    Ocg917 <= W6x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nfg917 <= 1'b0;
  else
    Nfg917 <= P6x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mig917 <= 1'b0;
  else
    Mig917 <= Ebx7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Llg917 <= 1'b0;
  else
    Llg917 <= Xax7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kog917 <= 1'b0;
  else
    Kog917 <= S4x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jrg917 <= 1'b0;
  else
    Jrg917 <= L4x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Iug917 <= 1'b0;
  else
    Iug917 <= A9x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hxg917 <= 1'b0;
  else
    Hxg917 <= Idx7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    F0h917 <= 1'b0;
  else
    F0h917 <= Bdx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D3h917 <= 1'b0;
  else
    D3h917 <= Y0x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    C6h917 <= 1'b0;
  else
    C6h917 <= R0x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B9h917 <= 1'b0;
  else
    B9h917 <= O9x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ach917 <= 1'b0;
  else
    Ach917 <= H9x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zeh917 <= 1'b0;
  else
    Zeh917 <= G5x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yhh917 <= 1'b0;
  else
    Yhh917 <= Z4x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xkh917 <= 1'b0;
  else
    Xkh917 <= Kt38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wnh917 <= 1'b0;
  else
    Wnh917 <= Dt38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vqh917 <= 1'b0;
  else
    Vqh917 <= Ov38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uth917 <= 1'b0;
  else
    Uth917 <= Hv38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Twh917 <= 1'b0;
  else
    Twh917 <= Sx38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Szh917 <= 1'b0;
  else
    Szh917 <= Lx38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R2i917 <= 1'b0;
  else
    R2i917 <= Q3x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q5i917 <= 1'b0;
  else
    Q5i917 <= J3x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P8i917 <= 1'b0;
  else
    P8i917 <= Y7x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Obi917 <= 1'b0;
  else
    Obi917 <= R7x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nei917 <= 1'b0;
  else
    Nei917 <= Gcx7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mhi917 <= 1'b0;
  else
    Mhi917 <= Zbx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lki917 <= 1'b0;
  else
    Lki917 <= Ovw7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kni917 <= 1'b0;
  else
    Kni917 <= Hvw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jqi917 <= 1'b0;
  else
    Jqi917 <= Cax7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Iti917 <= 1'b0;
  else
    Iti917 <= V9x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hwi917 <= 1'b0;
  else
    Hwi917 <= U5x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gzi917 <= 1'b0;
  else
    Gzi917 <= N5x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F2j917 <= 1'b0;
  else
    F2j917 <= M1x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    E5j917 <= 1'b0;
  else
    E5j917 <= F1x7v6;

always @(posedge FCLK) D8j917 <= Aai7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Naj917 <= 1'b0;
  else
    Naj917 <= Ogx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rcj917 <= 1'b0;
  else
    Rcj917 <= Cfk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qfj917 <= 1'b0;
  else
    Qfj917 <= Vek8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pij917 <= 1'b0;
  else
    Pij917 <= Egk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Olj917 <= 1'b0;
  else
    Olj917 <= Rtw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Noj917 <= 1'b0;
  else
    Noj917 <= Rqk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lrj917 <= 1'b0;
  else
    Lrj917 <= Su68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qtj917 <= 1'b0;
  else
    Qtj917 <= Lu68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vvj917 <= 1'b0;
  else
    Vvj917 <= Eu68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ayj917 <= 1'b0;
  else
    Ayj917 <= Xt68v6;

always @(posedge HCLK) F0k917 <= G2e8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    G2k917 <= 1'b0;
  else
    G2k917 <= C0e8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J4k917 <= 1'b0;
  else
    J4k917 <= Vzd8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M6k917 <= 1'b0;
  else
    M6k917 <= Qgc8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J8k917 <= 1'b0;
  else
    J8k917 <= Bsa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bck917 <= 1'b0;
  else
    Bck917 <= Ura8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nfk917 <= 1'b0;
  else
    Nfk917 <= Nra8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fjk917 <= 1'b0;
  else
    Fjk917 <= Gra8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Rmk917 <= 1'b0;
  else
    Rmk917 <= Zqa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jqk917 <= 1'b0;
  else
    Jqk917 <= Sqa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vtk917 <= 1'b0;
  else
    Vtk917 <= Lqa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nxk917 <= 1'b0;
  else
    Nxk917 <= Eqa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z0l917 <= 1'b0;
  else
    Z0l917 <= Xpa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R4l917 <= 1'b0;
  else
    R4l917 <= Qpa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D8l917 <= 1'b0;
  else
    D8l917 <= Jpa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vbl917 <= 1'b0;
  else
    Vbl917 <= Cpa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hfl917 <= 1'b0;
  else
    Hfl917 <= Voa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zil917 <= 1'b0;
  else
    Zil917 <= Ooa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lml917 <= 1'b0;
  else
    Lml917 <= Hoa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dql917 <= 1'b0;
  else
    Dql917 <= Aoa8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ptl917 <= 1'b0;
  else
    Ptl917 <= Fr68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Svl917 <= 1'b0;
  else
    Svl917 <= Qxo7v6;

always @(posedge HCLK) Yyl917 <= Pi68v6;
always @(posedge HCLK) P0m917 <= Ib68v6;
always @(posedge HCLK) F2m917 <= G368v6;
always @(posedge HCLK) V3m917 <= Ev58v6;
always @(posedge HCLK) L5m917 <= Cn58v6;
always @(posedge HCLK) B7m917 <= Af58v6;
always @(posedge HCLK) R8m917 <= Y658v6;
always @(posedge HCLK) Ham917 <= Wy48v6;
always @(posedge HCLK) Xbm917 <= Ir48v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ndm917 <= 1'b0;
  else
    Ndm917 <= X9y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nfm917 <= 1'b0;
  else
    Nfm917 <= E3y7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Phm917 <= 1'b0;
  else
    Phm917 <= Pvnet6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ikm917 <= 1'b0;
  else
    Ikm917 <= Grw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Emm917 <= 1'b0;
  else
    Emm917 <= Xee8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hom917 <= 1'b0;
  else
    Hom917 <= Efe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lqm917 <= 1'b0;
  else
    Lqm917 <= Lfe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Psm917 <= 1'b0;
  else
    Psm917 <= Sfe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tum917 <= 1'b0;
  else
    Tum917 <= Zfe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xwm917 <= 1'b0;
  else
    Xwm917 <= Gge8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bzm917 <= 1'b0;
  else
    Bzm917 <= Nge8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    F1n917 <= 1'b0;
  else
    F1n917 <= Uge8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J3n917 <= 1'b0;
  else
    J3n917 <= Bhe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O5n917 <= 1'b0;
  else
    O5n917 <= Ihe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T7n917 <= 1'b0;
  else
    T7n917 <= Phe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y9n917 <= 1'b0;
  else
    Y9n917 <= Whe8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Dcn917 <= 1'b0;
  else
    Dcn917 <= Die8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ien917 <= 1'b0;
  else
    Ien917 <= Kie8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ngn917 <= 1'b0;
  else
    Ngn917 <= Rie8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sin917 <= 1'b0;
  else
    Sin917 <= Yie8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xkn917 <= 1'b0;
  else
    Xkn917 <= Qee8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ann917 <= 1'b0;
  else
    Ann917 <= Jee8v6;

always @(posedge HCLK) Dpn917 <= J0e8v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ern917 <= 1'b0;
  else
    Ern917 <= Nic8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Btn917 <= 1'b0;
  else
    Btn917 <= B0a8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nwn917 <= 1'b0;
  else
    Nwn917 <= Uz98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zzn917 <= 1'b0;
  else
    Zzn917 <= Nz98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L3o917 <= 1'b0;
  else
    L3o917 <= Gz98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X6o917 <= 1'b0;
  else
    X6o917 <= Zy98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jao917 <= 1'b0;
  else
    Jao917 <= Sy98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vdo917 <= 1'b0;
  else
    Vdo917 <= Ly98v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hho917 <= 1'b0;
  else
    Hho917 <= Ey98v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tko917 <= 1'b0;
  else
    Tko917 <= D388v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vmo917 <= 1'b0;
  else
    Vmo917 <= I988v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Woo917 <= 1'b0;
  else
    Woo917 <= B988v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xqo917 <= 1'b0;
  else
    Xqo917 <= U888v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yso917 <= 1'b0;
  else
    Yso917 <= N888v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zuo917 <= 1'b0;
  else
    Zuo917 <= G888v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Axo917 <= 1'b0;
  else
    Axo917 <= Z788v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bzo917 <= 1'b0;
  else
    Bzo917 <= S788v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    C1p917 <= 1'b0;
  else
    C1p917 <= L788v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    D3p917 <= 1'b0;
  else
    D3p917 <= E788v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    E5p917 <= 1'b0;
  else
    E5p917 <= X688v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F7p917 <= 1'b0;
  else
    F7p917 <= Q688v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    H9p917 <= 1'b0;
  else
    H9p917 <= T9i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Nbp917 <= 1'b0;
  else
    Nbp917 <= Wv78v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Udp917 <= 1'b0;
  else
    Udp917 <= Pv78v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bgp917 <= 1'b0;
  else
    Bgp917 <= Iv78v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Iip917 <= 1'b0;
  else
    Iip917 <= Bv78v6;

always @(posedge FCLK) Pkp917 <= Lwq7v6;
always @(posedge FCLK) Dnp917 <= Uu78v6;
always @(posedge FCLK) Spp917 <= B8v7v6;
always @(posedge FCLK) Bsp917 <= I8v7v6;
always @(posedge FCLK) Kup917 <= P8v7v6;
always @(posedge FCLK) Twp917 <= W8v7v6;
always @(posedge FCLK) Czp917 <= D9v7v6;
always @(posedge FCLK) L1q917 <= K9v7v6;
always @(posedge FCLK) U3q917 <= R9v7v6;
always @(posedge FCLK) D6q917 <= Y9v7v6;
always @(posedge FCLK) M8q917 <= Fav7v6;
always @(posedge FCLK) Vaq917 <= Mav7v6;
always @(posedge FCLK) Edq917 <= Tav7v6;
always @(posedge FCLK) Nfq917 <= Abv7v6;
always @(posedge FCLK) Whq917 <= Hbv7v6;
always @(posedge FCLK) Fkq917 <= Obv7v6;
always @(posedge FCLK) Omq917 <= Vbv7v6;
always @(posedge FCLK) Xoq917 <= Ccv7v6;
always @(posedge FCLK) Grq917 <= Jcv7v6;
always @(posedge FCLK) Ptq917 <= Qcv7v6;
always @(posedge FCLK) Yvq917 <= Xcv7v6;
always @(posedge FCLK) Hyq917 <= Edv7v6;
always @(posedge FCLK) Q0r917 <= Ldv7v6;
always @(posedge FCLK) Z2r917 <= Sdv7v6;
always @(posedge FCLK) I5r917 <= Zdv7v6;
always @(posedge FCLK) Q7r917 <= Gev7v6;
always @(posedge FCLK) Y9r917 <= Nev7v6;
always @(posedge FCLK) Gcr917 <= Uev7v6;
always @(posedge FCLK) Oer917 <= Bfv7v6;
always @(posedge FCLK) Wgr917 <= Ifv7v6;
always @(posedge FCLK) Ejr917 <= Pfv7v6;
always @(posedge FCLK) Mlr917 <= Wfv7v6;
always @(posedge FCLK) Unr917 <= Dgv7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cqr917 <= 1'b0;
  else
    Cqr917 <= J688v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Esr917 <= 1'b0;
  else
    Esr917 <= C688v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gur917 <= 1'b0;
  else
    Gur917 <= V588v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Iwr917 <= 1'b0;
  else
    Iwr917 <= O588v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kyr917 <= 1'b0;
  else
    Kyr917 <= H588v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    M0s917 <= 1'b0;
  else
    M0s917 <= A588v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    O2s917 <= 1'b0;
  else
    O2s917 <= T488v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Q4s917 <= 1'b0;
  else
    Q4s917 <= M488v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    S6s917 <= 1'b0;
  else
    S6s917 <= F488v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    U8s917 <= 1'b0;
  else
    U8s917 <= Y388v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Was917 <= 1'b0;
  else
    Was917 <= R388v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ycs917 <= 1'b0;
  else
    Ycs917 <= K388v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Afs917 <= 1'b0;
  else
    Afs917 <= P288v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Chs917 <= 1'b0;
  else
    Chs917 <= I288v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ejs917 <= 1'b0;
  else
    Ejs917 <= B288v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gls917 <= 1'b0;
  else
    Gls917 <= U188v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ins917 <= 1'b0;
  else
    Ins917 <= M9i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lps917 <= 1'b0;
  else
    Lps917 <= Dw78v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Krs917 <= 1'b0;
  else
    Krs917 <= Nbr7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ats917 <= 1'b0;
  else
    Ats917 <= Gbr7v6;

always @(posedge FCLK) Tus917 <= F7r7v6;
always @(posedge FCLK) Qws917 <= O8r7v6;
always @(posedge FCLK) Nys917 <= V8r7v6;
always @(posedge FCLK) K0t917 <= J9r7v6;
always @(posedge FCLK) G2t917 <= Q9r7v6;
always @(posedge FCLK) C4t917 <= X9r7v6;
always @(posedge FCLK) Y5t917 <= Ear7v6;
always @(posedge FCLK) U7t917 <= Lar7v6;
always @(posedge FCLK) Q9t917 <= Sar7v6;
always @(posedge FCLK) Mbt917 <= Zar7v6;
always @(posedge FCLK) Idt917 <= P5r7v6;
always @(posedge FCLK) Fft917 <= I5r7v6;
always @(posedge FCLK) Cht917 <= B5r7v6;
always @(posedge FCLK) Zit917 <= T0r7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vkt917 <= 1'b0;
  else
    Vkt917 <= Boe7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Tmt917 <= 1'b0;
  else
    Tmt917 <= G1e7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Ipt917 <= 1'b0;
  else
    Ipt917 <= Cmg7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Xrt917 <= 1'b1;
  else
    Xrt917 <= Rte7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qtt917 <= 1'b0;
  else
    Qtt917 <= I6e7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bwt917 <= 1'b0;
  else
    Bwt917 <= Iyf7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Myt917 <= 1'b0;
  else
    Myt917 <= Zpe7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    K0u917 <= 1'b0;
  else
    K0u917 <= L8l8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    X2u917 <= 1'b0;
  else
    X2u917 <= Md1nz6[2];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    N5u917 <= 1'b0;
  else
    N5u917 <= X7g7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    D8u917 <= 1'b0;
  else
    D8u917 <= S8l8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qau917 <= 1'b0;
  else
    Qau917 <= Md1nz6[1];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gdu917 <= 1'b0;
  else
    Gdu917 <= L5g7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Wfu917 <= 1'b0;
  else
    Wfu917 <= Z8l8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jiu917 <= 1'b0;
  else
    Jiu917 <= Md1nz6[0];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zku917 <= 1'b0;
  else
    Zku917 <= Z2g7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Pnu917 <= 1'b0;
  else
    Pnu917 <= F9i7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Opu917 <= 1'b0;
  else
    Opu917 <= Y8i7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Mru917 <= 1'b0;
  else
    Mru917 <= Gpr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ktu917 <= 1'b0;
  else
    Ktu917 <= B5e7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yvu917 <= 1'b0;
  else
    Yvu917 <= P0g7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Myu917 <= 1'b0;
  else
    Myu917 <= Ame7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    N0v917 <= 1'b0;
  else
    N0v917 <= Xzd7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    F3v917 <= 1'b0;
  else
    F3v917 <= Nog7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    X5v917 <= 1'b0;
  else
    X5v917 <= R8i7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    R7v917 <= 1'b1;
  else
    R7v917 <= Zor7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    J9v917 <= 1'b0;
  else
    J9v917 <= K8i7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Ebv917 <= 1'b0;
  else
    Ebv917 <= Omr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rdv917 <= 1'b0;
  else
    Rdv917 <= Yb1nz6[2];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hgv917 <= 1'b0;
  else
    Hgv917 <= Hfg7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Xiv917 <= 1'b0;
  else
    Xiv917 <= Vmr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Klv917 <= 1'b0;
  else
    Klv917 <= Yb1nz6[1];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Aov917 <= 1'b0;
  else
    Aov917 <= Vcg7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Qqv917 <= 1'b0;
  else
    Qqv917 <= Cnr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dtv917 <= 1'b0;
  else
    Dtv917 <= Yb1nz6[0];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tvv917 <= 1'b0;
  else
    Tvv917 <= Jag7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Jyv917 <= 1'b0;
  else
    Jyv917 <= Yrr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    J0w917 <= 1'b1;
  else
    J0w917 <= Rrr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    G2w917 <= 1'b0;
  else
    G2w917 <= Msr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    G4w917 <= 1'b0;
  else
    G4w917 <= D8i7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    D6w917 <= 1'b0;
  else
    D6w917 <= W7i7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    A8w917 <= 1'b0;
  else
    A8w917 <= P7i7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    X9w917 <= 1'b0;
  else
    X9w917 <= I7i7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Rbw917 <= 1'b0;
  else
    Rbw917 <= Pqr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Ndw917 <= 1'b0;
  else
    Ndw917 <= Iqr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Jfw917 <= 1'b0;
  else
    Jfw917 <= Bqr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Fhw917 <= 1'b0;
  else
    Fhw917 <= Upr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Bjw917 <= 1'b0;
  else
    Bjw917 <= Npr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Ykw917 <= 1'b0;
  else
    Ykw917 <= B7i7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Smw917 <= 1'b0;
  else
    Smw917 <= Lor7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Pow917 <= 1'b0;
  else
    Pow917 <= Eor7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Qqw917 <= 1'b0;
  else
    Qqw917 <= Xnr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Rsw917 <= 1'b0;
  else
    Rsw917 <= Qnr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Suw917 <= 1'b0;
  else
    Suw917 <= Jnr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Tww917 <= 1'b0;
  else
    Tww917 <= U6i7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Oyw917 <= 1'b0;
  else
    Oyw917 <= Krr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    O0x917 <= 1'b0;
  else
    O0x917 <= Drr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    O2x917 <= 1'b0;
  else
    O2x917 <= Fsr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    O4x917 <= 1'b1;
  else
    O4x917 <= Wqr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    T6x917 <= 1'b0;
  else
    T6x917 <= M2e7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    E9x917 <= 1'b0;
  else
    E9x917 <= Vjg7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pbx917 <= 1'b0;
  else
    Pbx917 <= Hmr7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mdx917 <= 1'b1;
  else
    Mdx917 <= Pjr7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Efx917 <= 1'b1;
  else
    Efx917 <= Zhr7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dhx917 <= 1'b1;
  else
    Dhx917 <= Gir7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cjx917 <= 1'b1;
  else
    Cjx917 <= Nir7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Blx917 <= 1'b1;
  else
    Blx917 <= Uir7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Anx917 <= 1'b1;
  else
    Anx917 <= Bjr7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Zox917 <= 1'b0;
  else
    Zox917 <= N6i7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Wqx917 <= 1'b1;
  else
    Wqx917 <= Sor7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Osx917 <= 1'b0;
  else
    Osx917 <= G6i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jux917 <= 1'b0;
  else
    Jux917 <= N188v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lwx917 <= 1'b0;
  else
    Lwx917 <= G188v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Nyx917 <= 1'b0;
  else
    Nyx917 <= Z088v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    P0y917 <= 1'b0;
  else
    P0y917 <= Mr68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    S2y917 <= 1'b0;
  else
    S2y917 <= Tvo7v6;

always @(posedge HCLK) Y5y917 <= Sg68v6;
always @(posedge HCLK) P7y917 <= L968v6;
always @(posedge HCLK) F9y917 <= J168v6;
always @(posedge HCLK) Vay917 <= Ht58v6;
always @(posedge HCLK) Lcy917 <= Fl58v6;
always @(posedge HCLK) Bey917 <= Dd58v6;
always @(posedge HCLK) Rfy917 <= B558v6;
always @(posedge HCLK) Hhy917 <= Zw48v6;
always @(posedge HCLK) Xiy917 <= Lp48v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nky917 <= 1'b0;
  else
    Nky917 <= L3y7v6;

always @(posedge FCLK) Pmy917 <= E3r7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Moy917 <= 1'b0;
  else
    Moy917 <= Ntf8v6;

always @(posedge SWCLKTCK or negedge Sz9dt6)
  if(~Sz9dt6)
    Hqy917 <= 1'b0;
  else
    Hqy917 <= Gtf8v6;

always @(posedge C3a7z6 or negedge Sz9dt6)
  if(~Sz9dt6)
    Zry917 <= 1'b0;
  else
    Zry917 <= Lt57v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lty917 <= 1'b0;
  else
    Lty917 <= Jp38v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ovy917 <= 1'b0;
  else
    Ovy917 <= Hhw7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Uxy917 <= 1'b0;
  else
    Uxy917 <= Iew7v6;

always @(posedge FCLK) A0z917 <= Bew7v6;
always @(posedge FCLK) N2z917 <= Udw7v6;
always @(posedge FCLK) A5z917 <= Ndw7v6;
always @(posedge FCLK) N7z917 <= Zcw7v6;
always @(posedge FCLK) Aaz917 <= Scw7v6;
always @(posedge FCLK) Ncz917 <= Ecw7v6;
always @(posedge FCLK) Afz917 <= Xbw7v6;
always @(posedge FCLK) Nhz917 <= Qbw7v6;
always @(posedge FCLK) Bkz917 <= Jbw7v6;
always @(posedge FCLK) Pmz917 <= Vaw7v6;
always @(posedge FCLK) Dpz917 <= Oaw7v6;
always @(posedge FCLK) Rrz917 <= Aaw7v6;
always @(posedge FCLK) Fuz917 <= T9w7v6;
always @(posedge FCLK) Twz917 <= M9w7v6;
always @(posedge FCLK) Hzz917 <= F9w7v6;
always @(posedge FCLK) V10a17 <= R8w7v6;
always @(posedge FCLK) J40a17 <= K8w7v6;
always @(posedge FCLK) X60a17 <= W7w7v6;
always @(posedge FCLK) L90a17 <= P7w7v6;
always @(posedge FCLK) Zb0a17 <= I7w7v6;
always @(posedge FCLK) Ne0a17 <= B7w7v6;
always @(posedge FCLK) Bh0a17 <= N6w7v6;
always @(posedge FCLK) Pj0a17 <= G6w7v6;
always @(posedge FCLK) Dm0a17 <= Z5w7v6;
always @(posedge FCLK) Qo0a17 <= S5w7v6;
always @(posedge FCLK) Dr0a17 <= L5w7v6;
always @(posedge FCLK) Ot0a17 <= E5w7v6;
always @(posedge FCLK) Bw0a17 <= X4w7v6;
always @(posedge FCLK) Oy0a17 <= Q4w7v6;
always @(posedge HCLK) B11a17 <= Ito7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R31a17 <= 1'b0;
  else
    R31a17 <= Zgddt6;

always @(posedge HCLK) N61a17 <= C4p7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R91a17 <= 1'b0;
  else
    R91a17 <= Cjo7v6;

always @(posedge FCLK) Jb1a17 <= U6w7v6;
always @(posedge FCLK) Xd1a17 <= Y8w7v6;
always @(posedge FCLK) Lg1a17 <= Cbw7v6;
always @(posedge FCLK) Zi1a17 <= Gdw7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ml1a17 <= 1'b0;
  else
    Ml1a17 <= Wbs7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Po1a17 <= 1'b0;
  else
    Po1a17 <= Gr38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Or1a17 <= 1'b0;
  else
    Or1a17 <= Zq38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nu1a17 <= 1'b0;
  else
    Nu1a17 <= Sq38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mx1a17 <= 1'b0;
  else
    Mx1a17 <= Lq38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L02a17 <= 1'b0;
  else
    L02a17 <= Wzw7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    K32a17 <= 1'b0;
  else
    K32a17 <= Pzw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J62a17 <= 1'b0;
  else
    J62a17 <= Uyw7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    I92a17 <= 1'b0;
  else
    I92a17 <= Nyw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hc2a17 <= 1'b0;
  else
    Hc2a17 <= Kjk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gf2a17 <= 1'b0;
  else
    Gf2a17 <= Q8s7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ki2a17 <= 1'b0;
  else
    Ki2a17 <= K0x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jl2a17 <= 1'b0;
  else
    Jl2a17 <= D0x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Io2a17 <= 1'b0;
  else
    Io2a17 <= E4x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hr2a17 <= 1'b0;
  else
    Hr2a17 <= X3x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gu2a17 <= 1'b0;
  else
    Gu2a17 <= M8x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fx2a17 <= 1'b0;
  else
    Fx2a17 <= F8x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    E03a17 <= 1'b0;
  else
    E03a17 <= Ucx7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    D33a17 <= 1'b0;
  else
    D33a17 <= Ncx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    C63a17 <= 1'b0;
  else
    C63a17 <= Gy38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    B93a17 <= 1'b0;
  else
    B93a17 <= Zx38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ac3a17 <= 1'b0;
  else
    Ac3a17 <= K048v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ze3a17 <= 1'b0;
  else
    Ze3a17 <= D048v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yh3a17 <= 1'b0;
  else
    Yh3a17 <= O248v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xk3a17 <= 1'b0;
  else
    Xk3a17 <= H248v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wn3a17 <= 1'b0;
  else
    Wn3a17 <= S448v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vq3a17 <= 1'b0;
  else
    Vq3a17 <= L448v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ut3a17 <= 1'b0;
  else
    Ut3a17 <= Izw7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tw3a17 <= 1'b0;
  else
    Tw3a17 <= Bzw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sz3a17 <= 1'b0;
  else
    Sz3a17 <= C3x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    R24a17 <= 1'b0;
  else
    R24a17 <= V2x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q54a17 <= 1'b0;
  else
    Q54a17 <= K7x7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    P84a17 <= 1'b0;
  else
    P84a17 <= D7x7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ob4a17 <= 1'b0;
  else
    Ob4a17 <= Sbx7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ne4a17 <= 1'b0;
  else
    Ne4a17 <= Lbx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mh4a17 <= 1'b0;
  else
    Mh4a17 <= Gyw7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lk4a17 <= 1'b0;
  else
    Lk4a17 <= Zxw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kn4a17 <= 1'b0;
  else
    Kn4a17 <= Wz38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jq4a17 <= 1'b0;
  else
    Jq4a17 <= Pz38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    It4a17 <= 1'b0;
  else
    It4a17 <= A248v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hw4a17 <= 1'b0;
  else
    Hw4a17 <= T148v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gz4a17 <= 1'b0;
  else
    Gz4a17 <= E448v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    F25a17 <= 1'b0;
  else
    F25a17 <= X348v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    E55a17 <= 1'b0;
  else
    E55a17 <= Zgk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    C85a17 <= 1'b0;
  else
    C85a17 <= Sxw7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bb5a17 <= 1'b0;
  else
    Bb5a17 <= Lxw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ae5a17 <= 1'b0;
  else
    Ae5a17 <= Is38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Zg5a17 <= 1'b0;
  else
    Zg5a17 <= Bs38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yj5a17 <= 1'b0;
  else
    Yj5a17 <= Qw38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xm5a17 <= 1'b0;
  else
    Xm5a17 <= Mu38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wp5a17 <= 1'b0;
  else
    Wp5a17 <= Fu38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vs5a17 <= 1'b0;
  else
    Vs5a17 <= Exw7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uv5a17 <= 1'b0;
  else
    Uv5a17 <= Xww7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ty5a17 <= 1'b0;
  else
    Ty5a17 <= Iz38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    S16a17 <= 1'b0;
  else
    S16a17 <= Bz38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R46a17 <= 1'b0;
  else
    R46a17 <= Q348v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q76a17 <= 1'b0;
  else
    Q76a17 <= J348v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pa6a17 <= 1'b0;
  else
    Pa6a17 <= M148v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Od6a17 <= 1'b0;
  else
    Od6a17 <= F148v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ng6a17 <= 1'b0;
  else
    Ng6a17 <= Ghk8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lj6a17 <= 1'b0;
  else
    Lj6a17 <= Nhk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jm6a17 <= 1'b0;
  else
    Jm6a17 <= Qww7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ip6a17 <= 1'b0;
  else
    Ip6a17 <= Ur38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hs6a17 <= 1'b0;
  else
    Hs6a17 <= Nr38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gv6a17 <= 1'b0;
  else
    Gv6a17 <= Yt38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fy6a17 <= 1'b0;
  else
    Fy6a17 <= Rt38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    E17a17 <= 1'b0;
  else
    E17a17 <= Wik8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    I37a17 <= 1'b0;
  else
    I37a17 <= Cw38v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    H67a17 <= 1'b0;
  else
    H67a17 <= Vv38v6;

always @(posedge FCLK) G97a17 <= Z5i7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qb7a17 <= 1'b0;
  else
    Qb7a17 <= Hgx7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ud7a17 <= 1'b0;
  else
    Ud7a17 <= Zxymz6[4];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bg7a17 <= 1'b0;
  else
    Bg7a17 <= Rwa7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ei7a17 <= 1'b0;
  else
    Ei7a17 <= W8zmz6[1];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ik7a17 <= 1'b0;
  else
    Ik7a17 <= Jc87v6;

always @(posedge HCLK) Gm7a17 <= Jru7v6;
always @(posedge HCLK) Fo7a17 <= Cru7v6;
always @(posedge HCLK) Eq7a17 <= Vqu7v6;
always @(posedge HCLK) Ds7a17 <= Oqu7v6;
always @(posedge HCLK) Cu7a17 <= Hqu7v6;
always @(posedge HCLK) Bw7a17 <= Yxk8v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zx7a17 <= 1'b0;
  else
    Zx7a17 <= G287v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tz7a17 <= 1'b0;
  else
    Tz7a17 <= T1zmz6[33];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    B28a17 <= 1'b0;
  else
    B28a17 <= K9a7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    A48a17 <= 1'b0;
  else
    A48a17 <= Oga7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    O68a17 <= 1'b0;
  else
    O68a17 <= Hju7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    O88a17 <= 1'b0;
  else
    O88a17 <= Aju7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ma8a17 <= 1'b0;
  else
    Ma8a17 <= Tiu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kc8a17 <= 1'b0;
  else
    Kc8a17 <= Miu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ie8a17 <= 1'b0;
  else
    Ie8a17 <= Fiu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gg8a17 <= 1'b0;
  else
    Gg8a17 <= Yhu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ei8a17 <= 1'b0;
  else
    Ei8a17 <= Wgu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ck8a17 <= 1'b0;
  else
    Ck8a17 <= Dhu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Am8a17 <= 1'b0;
  else
    Am8a17 <= Pgu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yn8a17 <= 1'b0;
  else
    Yn8a17 <= Khu7v6;

always @(posedge HCLK) Wp8a17 <= Oha7z6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Nr8a17 <= 1'b0;
  else
    Nr8a17 <= Igu7v6;

always @(posedge HCLK) Mt8a17 <= Gha7z6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dv8a17 <= 1'b0;
  else
    Dv8a17 <= Bgu7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cx8a17 <= 1'b0;
  else
    Cx8a17 <= T1zmz6[32];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kz8a17 <= 1'b0;
  else
    Kz8a17 <= Qea7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    M19a17 <= 1'b0;
  else
    M19a17 <= Ufu7v6;

always @(posedge HCLK) L39a17 <= Acu7v6;
always @(posedge HCLK) I59a17 <= P9u7v6;
always @(posedge HCLK) F79a17 <= Hcu7v6;
always @(posedge HCLK) C99a17 <= W9u7v6;
always @(posedge HCLK) Za9a17 <= Mho7v6;
always @(posedge HCLK) Qc9a17 <= Rbt7v6;
always @(posedge HCLK) Ne9a17 <= Ybt7v6;
always @(posedge HCLK) Kg9a17 <= Fct7v6;
always @(posedge HCLK) Hi9a17 <= N1u7v6;
always @(posedge HCLK) Ek9a17 <= U1u7v6;
always @(posedge HCLK) Bm9a17 <= B2u7v6;
always @(posedge HCLK) Yn9a17 <= Pot7v6;
always @(posedge HCLK) Vp9a17 <= Wot7v6;
always @(posedge HCLK) Sr9a17 <= Dpt7v6;
always @(posedge HCLK) Pt9a17 <= Leu7v6;
always @(posedge HCLK) Mv9a17 <= Seu7v6;
always @(posedge HCLK) Jx9a17 <= Zeu7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gz9a17 <= 1'b0;
  else
    Gz9a17 <= Zxymz6[3];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    N1aa17 <= 1'b0;
  else
    N1aa17 <= Zxymz6[0];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    U3aa17 <= 1'b0;
  else
    U3aa17 <= Zxymz6[1];

always @(posedge HCLK) B6aa17 <= P3t7v6;
always @(posedge HCLK) Y7aa17 <= W3t7v6;
always @(posedge HCLK) V9aa17 <= D4t7v6;
always @(posedge HCLK) Sbaa17 <= Ltt7v6;
always @(posedge HCLK) Pdaa17 <= Stt7v6;
always @(posedge HCLK) Mfaa17 <= Ztt7v6;
always @(posedge HCLK) Jhaa17 <= Bat7v6;
always @(posedge HCLK) Gjaa17 <= Iat7v6;
always @(posedge HCLK) Dlaa17 <= Pat7v6;
always @(posedge HCLK) Anaa17 <= Xzt7v6;
always @(posedge HCLK) Xoaa17 <= E0u7v6;
always @(posedge HCLK) Uqaa17 <= L0u7v6;
always @(posedge HCLK) Rsaa17 <= Ngt7v6;
always @(posedge HCLK) Ouaa17 <= Ugt7v6;
always @(posedge HCLK) Lwaa17 <= Bht7v6;
always @(posedge HCLK) Iyaa17 <= J6u7v6;
always @(posedge HCLK) F0ba17 <= Q6u7v6;
always @(posedge HCLK) C2ba17 <= X6u7v6;
always @(posedge HCLK) Z3ba17 <= Zmt7v6;
always @(posedge HCLK) W5ba17 <= Gnt7v6;
always @(posedge HCLK) T7ba17 <= Nnt7v6;
always @(posedge HCLK) Q9ba17 <= Vcu7v6;
always @(posedge HCLK) Nbba17 <= Cdu7v6;
always @(posedge HCLK) Kdba17 <= Jdu7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hfba17 <= 1'b0;
  else
    Hfba17 <= Zxymz6[2];

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ohba17 <= 1'b0;
  else
    Ohba17 <= Gas7v6;

always @(posedge FCLK) Skba17 <= J2r7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pmba17 <= 1'b0;
  else
    Pmba17 <= C8s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tpba17 <= 1'b0;
  else
    Tpba17 <= Svr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rrba17 <= 1'b0;
  else
    Rrba17 <= Tsr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ptba17 <= 1'b0;
  else
    Ptba17 <= Nvk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pvba17 <= 1'b0;
  else
    Pvba17 <= Gvk8v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pxba17 <= 1'b0;
  else
    Pxba17 <= T1zmz6[30];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xzba17 <= 1'b0;
  else
    Xzba17 <= T1zmz6[22];

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F2ca17 <= 1'b0;
  else
    F2ca17 <= T1zmz6[14];

always @(posedge HCLK) N4ca17 <= U2t7v6;
always @(posedge HCLK) K6ca17 <= B3t7v6;
always @(posedge HCLK) H8ca17 <= I3t7v6;
always @(posedge HCLK) Eaca17 <= Qst7v6;
always @(posedge HCLK) Bcca17 <= Xst7v6;
always @(posedge HCLK) Ydca17 <= Ett7v6;
always @(posedge HCLK) Vfca17 <= G9t7v6;
always @(posedge HCLK) Shca17 <= N9t7v6;
always @(posedge HCLK) Pjca17 <= U9t7v6;
always @(posedge HCLK) Mlca17 <= Czt7v6;
always @(posedge HCLK) Jnca17 <= Jzt7v6;
always @(posedge HCLK) Gpca17 <= Qzt7v6;
always @(posedge HCLK) Drca17 <= Sft7v6;
always @(posedge HCLK) Atca17 <= Zft7v6;
always @(posedge HCLK) Xuca17 <= Ggt7v6;
always @(posedge HCLK) Uwca17 <= O5u7v6;
always @(posedge HCLK) Ryca17 <= V5u7v6;
always @(posedge HCLK) O0da17 <= C6u7v6;
always @(posedge HCLK) L2da17 <= Emt7v6;
always @(posedge HCLK) I4da17 <= Lmt7v6;
always @(posedge HCLK) F6da17 <= Smt7v6;
always @(posedge HCLK) C8da17 <= K4t7v6;
always @(posedge HCLK) Z9da17 <= R4t7v6;
always @(posedge HCLK) Wbda17 <= Y4t7v6;
always @(posedge HCLK) Tdda17 <= Gut7v6;
always @(posedge HCLK) Qfda17 <= Nut7v6;
always @(posedge HCLK) Nhda17 <= Uut7v6;
always @(posedge HCLK) Kjda17 <= Wat7v6;
always @(posedge HCLK) Hlda17 <= Dbt7v6;
always @(posedge HCLK) Enda17 <= Kbt7v6;
always @(posedge HCLK) Bpda17 <= S0u7v6;
always @(posedge HCLK) Yqda17 <= Z0u7v6;
always @(posedge HCLK) Vsda17 <= G1u7v6;
always @(posedge HCLK) Suda17 <= Iht7v6;
always @(posedge HCLK) Pwda17 <= Pht7v6;
always @(posedge HCLK) Myda17 <= Wht7v6;
always @(posedge HCLK) J0ea17 <= E7u7v6;
always @(posedge HCLK) G2ea17 <= L7u7v6;
always @(posedge HCLK) D4ea17 <= S7u7v6;
always @(posedge HCLK) A6ea17 <= Unt7v6;
always @(posedge HCLK) X7ea17 <= Bot7v6;
always @(posedge HCLK) U9ea17 <= Iot7v6;
always @(posedge HCLK) Rbea17 <= Qdu7v6;
always @(posedge HCLK) Odea17 <= Xdu7v6;
always @(posedge HCLK) Lfea17 <= Eeu7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ihea17 <= 1'b0;
  else
    Ihea17 <= E2s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Djea17 <= 1'b0;
  else
    Djea17 <= X1s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Blea17 <= 1'b0;
  else
    Blea17 <= Tzr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zmea17 <= 1'b0;
  else
    Zmea17 <= Pxr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xoea17 <= 1'b0;
  else
    Xoea17 <= Pfo7v6;

always @(posedge HCLK) Xqea17 <= F787v6;
always @(posedge HCLK) Tsea17 <= F9p7v6;
always @(posedge HCLK) Wvea17 <= Pis7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kyea17 <= 1'b0;
  else
    Kyea17 <= Aes7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    J1fa17 <= 1'b0;
  else
    J1fa17 <= Mds7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    I4fa17 <= 1'b0;
  else
    I4fa17 <= Tds7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H7fa17 <= 1'b0;
  else
    H7fa17 <= Kzb8v6;

always @(posedge FCLK) Uafa17 <= Jz78v6;
always @(posedge FCLK) Bdfa17 <= L088v6;
always @(posedge FCLK) Iffa17 <= E088v6;
always @(posedge FCLK) Phfa17 <= Xz78v6;
always @(posedge FCLK) Wjfa17 <= Qz78v6;
always @(posedge FCLK) Dmfa17 <= Cz78v6;
always @(posedge FCLK) Kofa17 <= Vy78v6;
always @(posedge FCLK) Rqfa17 <= Oy78v6;
always @(posedge FCLK) Ysfa17 <= Swq7v6;
always @(posedge FCLK) Mvfa17 <= Fx78v6;
always @(posedge FCLK) Uxfa17 <= Ay78v6;
always @(posedge FCLK) C0ga17 <= Tx78v6;
always @(posedge FCLK) K2ga17 <= Mx78v6;
always @(posedge FCLK) S4ga17 <= Yw78v6;
always @(posedge FCLK) A7ga17 <= Rw78v6;
always @(posedge FCLK) I9ga17 <= Kw78v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qbga17 <= 1'b0;
  else
    Qbga17 <= Jl78v6;

always @(posedge HCLK) Ndga17 <= Oe68v6;
always @(posedge HCLK) Cfga17 <= M668v6;
always @(posedge HCLK) Rgga17 <= Ky58v6;
always @(posedge HCLK) Giga17 <= Iq58v6;
always @(posedge HCLK) Vjga17 <= Gi58v6;
always @(posedge HCLK) Klga17 <= Ea58v6;
always @(posedge HCLK) Zmga17 <= C258v6;
always @(posedge HCLK) Ooga17 <= Ou48v6;
always @(posedge FCLK) Dqga17 <= Jjv7v6;
always @(posedge FCLK) Jsga17 <= Fhv7v6;
always @(posedge FCLK) Puga17 <= H8r7v6;
always @(posedge HCLK) Mwga17 <= S5i7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bzga17 <= 1'b0;
  else
    Bzga17 <= Phd7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V0ha17 <= 1'b0;
  else
    V0ha17 <= Mwu7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V2ha17 <= 1'b0;
  else
    V2ha17 <= Byx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X5ha17 <= 1'b0;
  else
    X5ha17 <= Uxx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z8ha17 <= 1'b0;
  else
    Z8ha17 <= Azs7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qbha17 <= 1'b0;
  else
    Qbha17 <= Yck8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ieha17 <= 1'b0;
  else
    Ieha17 <= Iri8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ahha17 <= 1'b0;
  else
    Ahha17 <= Ksi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sjha17 <= 1'b0;
  else
    Sjha17 <= Uqi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Omha17 <= 1'b0;
  else
    Omha17 <= Pri8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gpha17 <= 1'b0;
  else
    Gpha17 <= Wri8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yrha17 <= 1'b0;
  else
    Yrha17 <= Dsi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Quha17 <= 1'b0;
  else
    Quha17 <= Bri8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mxha17 <= 1'b0;
  else
    Mxha17 <= Rm38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L0ia17 <= 1'b0;
  else
    L0ia17 <= Ym38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K3ia17 <= 1'b0;
  else
    K3ia17 <= Fn38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J6ia17 <= 1'b0;
  else
    J6ia17 <= Mn38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    I9ia17 <= 1'b0;
  else
    I9ia17 <= Tn38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hcia17 <= 1'b0;
  else
    Hcia17 <= Ao38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Gfia17 <= 1'b0;
  else
    Gfia17 <= Oo38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fiia17 <= 1'b0;
  else
    Fiia17 <= Ho38v6;

always @(posedge HCLK) Elia17 <= Lfl8v6;
always @(posedge HCLK) Ynia17 <= Fg38v6;
always @(posedge HCLK) Sqia17 <= Yf38v6;
always @(posedge HCLK) Ntia17 <= Rf38v6;
always @(posedge HCLK) Iwia17 <= Kf38v6;
always @(posedge HCLK) Dzia17 <= Df38v6;
always @(posedge HCLK) Y1ja17 <= We38v6;
always @(posedge HCLK) T4ja17 <= Pe38v6;
always @(posedge HCLK) O7ja17 <= Ie38v6;
always @(posedge HCLK) Jaja17 <= Mdk8v6;
always @(posedge HCLK) Hdja17 <= Msy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fgja17 <= 1'b0;
  else
    Fgja17 <= C1d8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ejja17 <= 1'b0;
  else
    Ejja17 <= Cmk8v6;

always @(posedge HCLK) Mlja17 <= C1z7v6;
always @(posedge HCLK) Vnja17 <= Pxy7v6;
always @(posedge HCLK) Sqja17 <= Sqw7v6;
always @(posedge HCLK) Ptja17 <= Jny7v6;
always @(posedge HCLK) Mwja17 <= Rry7v6;
always @(posedge HCLK) Jzja17 <= Yry7v6;
always @(posedge HCLK) G2ka17 <= Fsy7v6;
always @(posedge HCLK) D5ka17 <= Aty7v6;
always @(posedge HCLK) A8ka17 <= Vty7v6;
always @(posedge HCLK) Xaka17 <= Juy7v6;
always @(posedge HCLK) Vdka17 <= Upy7v6;
always @(posedge HCLK) Tgka17 <= Bqy7v6;
always @(posedge HCLK) Qjka17 <= Iqy7v6;
always @(posedge HCLK) Nmka17 <= Cny7v6;
always @(posedge HCLK) Lpka17 <= Wqy7v6;
always @(posedge HCLK) Jska17 <= Kry7v6;
always @(posedge HCLK) Hvka17 <= Tsy7v6;
always @(posedge HCLK) Fyka17 <= Oty7v6;
always @(posedge HCLK) D1la17 <= Pqy7v6;
always @(posedge HCLK) B4la17 <= Vmy7v6;
always @(posedge HCLK) Z6la17 <= Dry7v6;
always @(posedge HCLK) X9la17 <= Evy7v6;
always @(posedge HCLK) Vcla17 <= Hty7v6;
always @(posedge HCLK) Tfla17 <= Cuy7v6;
always @(posedge HCLK) Rila17 <= Npy7v6;
always @(posedge HCLK) Plla17 <= Uwy7v6;
always @(posedge HCLK) Nola17 <= Bxy7v6;
always @(posedge HCLK) Lrla17 <= Dck8v6;
always @(posedge HCLK) Jula17 <= Quy7v6;
always @(posedge HCLK) Hxla17 <= Xuy7v6;
always @(posedge HCLK) F0ma17 <= Njx7v6;
always @(posedge HCLK) Z2ma17 <= Gjx7v6;
always @(posedge HCLK) T5ma17 <= Zix7v6;
always @(posedge HCLK) N8ma17 <= Six7v6;
always @(posedge HCLK) Ibma17 <= Lix7v6;
always @(posedge HCLK) Dema17 <= Eix7v6;
always @(posedge HCLK) Ygma17 <= Xhx7v6;
always @(posedge HCLK) Tjma17 <= Qhx7v6;
always @(posedge HCLK) Omma17 <= Jhx7v6;
always @(posedge HCLK) Jpma17 <= Rck8v6;
always @(posedge HCLK) Gsma17 <= Eii8v6;
always @(posedge HCLK) Dvma17 <= Lii8v6;
always @(posedge HCLK) Ayma17 <= Sii8v6;
always @(posedge HCLK) X0na17 <= Zii8v6;
always @(posedge HCLK) U3na17 <= Gji8v6;
always @(posedge HCLK) R6na17 <= Nji8v6;
always @(posedge HCLK) O9na17 <= Uji8v6;
always @(posedge HCLK) Lcna17 <= Bki8v6;
always @(posedge HCLK) Ifna17 <= Iki8v6;
always @(posedge HCLK) Fina17 <= Pki8v6;
always @(posedge HCLK) Dlna17 <= Wki8v6;
always @(posedge HCLK) Bona17 <= Dli8v6;
always @(posedge HCLK) Zqna17 <= Kli8v6;
always @(posedge HCLK) Xtna17 <= Rli8v6;
always @(posedge HCLK) Vwna17 <= Yli8v6;
always @(posedge HCLK) Tzna17 <= Fmi8v6;
always @(posedge HCLK) R2oa17 <= Mmi8v6;
always @(posedge HCLK) P5oa17 <= Tmi8v6;
always @(posedge HCLK) N8oa17 <= Ani8v6;
always @(posedge HCLK) Lboa17 <= Hni8v6;
always @(posedge HCLK) Jeoa17 <= Oni8v6;
always @(posedge HCLK) Hhoa17 <= Vni8v6;
always @(posedge HCLK) Fkoa17 <= Coi8v6;
always @(posedge HCLK) Dnoa17 <= Joi8v6;
always @(posedge HCLK) Bqoa17 <= Qoi8v6;
always @(posedge HCLK) Zsoa17 <= Xoi8v6;
always @(posedge HCLK) Xvoa17 <= Epi8v6;
always @(posedge HCLK) Vyoa17 <= Lpi8v6;
always @(posedge HCLK) T1pa17 <= Wbk8v6;
always @(posedge HCLK) R4pa17 <= Ydy7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O7pa17 <= 1'b0;
  else
    O7pa17 <= Okl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oapa17 <= 1'b0;
  else
    Oapa17 <= P0p7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tdpa17 <= 1'b0;
  else
    Tdpa17 <= Lnk8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Agpa17 <= 1'b0;
  else
    Agpa17 <= Gxx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kipa17 <= 1'b0;
  else
    Kipa17 <= Lwx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ukpa17 <= 1'b0;
  else
    Ukpa17 <= Swx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Enpa17 <= 1'b0;
  else
    Enpa17 <= Nxx7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oppa17 <= 1'b0;
  else
    Oppa17 <= Tuw7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Mspa17 <= 1'b0;
  else
    Mspa17 <= Avw7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kvpa17 <= 1'b0;
  else
    Kvpa17 <= S1get6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pxpa17 <= 1'b0;
  else
    Pxpa17 <= Xai8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    M0qa17 <= 1'b0;
  else
    M0qa17 <= Nlv7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O2qa17 <= 1'b0;
  else
    O2qa17 <= Bve8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    G4qa17 <= 1'b0;
  else
    G4qa17 <= Q7l8v6;

always @(posedge FCLK) I6qa17 <= Glv7v6;
always @(posedge FCLK) S8qa17 <= Zkv7v6;
always @(posedge FCLK) Jbqa17 <= Skv7v6;
always @(posedge FCLK) Aeqa17 <= U7v7v6;
always @(posedge FCLK) Lgqa17 <= N7v7v6;
always @(posedge FCLK) Wiqa17 <= G7v7v6;
always @(posedge FCLK) Hlqa17 <= Z6v7v6;
always @(posedge FCLK) Snqa17 <= S6v7v6;
always @(posedge FCLK) Dqqa17 <= L6v7v6;
always @(posedge FCLK) Osqa17 <= E6v7v6;
always @(posedge FCLK) Zuqa17 <= X5v7v6;
always @(posedge FCLK) Kxqa17 <= Q5v7v6;
always @(posedge FCLK) Vzqa17 <= J5v7v6;
always @(posedge FCLK) G2ra17 <= C5v7v6;
always @(posedge FCLK) S4ra17 <= V4v7v6;
always @(posedge FCLK) E7ra17 <= O4v7v6;
always @(posedge FCLK) Q9ra17 <= H4v7v6;
always @(posedge FCLK) Ccra17 <= A4v7v6;
always @(posedge FCLK) Oera17 <= T3v7v6;
always @(posedge FCLK) Ahra17 <= M3v7v6;
always @(posedge FCLK) Mjra17 <= F3v7v6;
always @(posedge FCLK) Ylra17 <= Y2v7v6;
always @(posedge FCLK) Kora17 <= R2v7v6;
always @(posedge FCLK) Wqra17 <= K2v7v6;
always @(posedge FCLK) Itra17 <= D2v7v6;
always @(posedge FCLK) Uvra17 <= W1v7v6;
always @(posedge FCLK) Gyra17 <= P1v7v6;
always @(posedge FCLK) S0sa17 <= I1v7v6;
always @(posedge FCLK) E3sa17 <= B1v7v6;
always @(posedge FCLK) Q5sa17 <= U0v7v6;
always @(posedge FCLK) C8sa17 <= N0v7v6;
always @(posedge FCLK) Oasa17 <= G0v7v6;
always @(posedge FCLK) Adsa17 <= Zzu7v6;
always @(posedge FCLK) Mfsa17 <= Szu7v6;
always @(posedge FCLK) Yhsa17 <= Lzu7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kksa17 <= 1'b0;
  else
    Kksa17 <= Yzq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rnsa17 <= 1'b0;
  else
    Rnsa17 <= Wyq7v6;

always @(posedge FCLK) Arsa17 <= Shr7v6;
always @(posedge FCLK) Tssa17 <= Xgr7v6;
always @(posedge FCLK) Musa17 <= Qgr7v6;
always @(posedge FCLK) Fwsa17 <= Jgr7v6;
always @(posedge FCLK) Yxsa17 <= Cgr7v6;
always @(posedge FCLK) Rzsa17 <= Vfr7v6;
always @(posedge FCLK) K1ta17 <= Ofr7v6;
always @(posedge FCLK) D3ta17 <= Hfr7v6;
always @(posedge FCLK) W4ta17 <= Afr7v6;
always @(posedge FCLK) P6ta17 <= Ter7v6;
always @(posedge FCLK) I8ta17 <= Mer7v6;
always @(posedge FCLK) Cata17 <= Fer7v6;
always @(posedge FCLK) Wbta17 <= Ydr7v6;
always @(posedge FCLK) Qdta17 <= Rdr7v6;
always @(posedge FCLK) Kfta17 <= Kdr7v6;
always @(posedge FCLK) Ehta17 <= Ddr7v6;
always @(posedge FCLK) Yita17 <= Wcr7v6;
always @(posedge FCLK) Skta17 <= Pcr7v6;
always @(posedge FCLK) Mmta17 <= Icr7v6;
always @(posedge FCLK) Gota17 <= Lhr7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Aqta17 <= 1'b1;
  else
    Aqta17 <= Mup7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Trta17 <= 1'b0;
  else
    Trta17 <= Fho7v6;

always @(posedge FCLK) Qtta17 <= D7q7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ivta17 <= 1'b0;
  else
    Ivta17 <= W6q7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bxta17 <= 1'b0;
  else
    Bxta17 <= Fcl8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yyta17 <= 1'b0;
  else
    Yyta17 <= D847v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Q0ua17 <= 1'b0;
  else
    Q0ua17 <= L5i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    L2ua17 <= 1'b0;
  else
    L2ua17 <= E5i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    H4ua17 <= 1'b0;
  else
    H4ua17 <= X4i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    D6ua17 <= 1'b0;
  else
    D6ua17 <= Q4i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Z7ua17 <= 1'b0;
  else
    Z7ua17 <= J4i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    V9ua17 <= 1'b0;
  else
    V9ua17 <= C4i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rbua17 <= 1'b0;
  else
    Rbua17 <= V3i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ndua17 <= 1'b0;
  else
    Ndua17 <= O3i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jfua17 <= 1'b0;
  else
    Jfua17 <= H3i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fhua17 <= 1'b0;
  else
    Fhua17 <= A3i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bjua17 <= 1'b0;
  else
    Bjua17 <= T2i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xkua17 <= 1'b0;
  else
    Xkua17 <= M2i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tmua17 <= 1'b0;
  else
    Tmua17 <= F2i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Poua17 <= 1'b0;
  else
    Poua17 <= Y1i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lqua17 <= 1'b0;
  else
    Lqua17 <= R1i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hsua17 <= 1'b0;
  else
    Hsua17 <= K1i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Duua17 <= 1'b0;
  else
    Duua17 <= D1i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zvua17 <= 1'b0;
  else
    Zvua17 <= W0i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vxua17 <= 1'b0;
  else
    Vxua17 <= P0i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rzua17 <= 1'b0;
  else
    Rzua17 <= I0i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    N1va17 <= 1'b0;
  else
    N1va17 <= B0i7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    J3va17 <= 1'b0;
  else
    J3va17 <= Uzh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F5va17 <= 1'b0;
  else
    F5va17 <= Nzh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    B7va17 <= 1'b0;
  else
    B7va17 <= Gzh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    X8va17 <= 1'b0;
  else
    X8va17 <= Zyh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tava17 <= 1'b0;
  else
    Tava17 <= Syh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pcva17 <= 1'b0;
  else
    Pcva17 <= Lyh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Leva17 <= 1'b0;
  else
    Leva17 <= Eyh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Hgva17 <= 1'b0;
  else
    Hgva17 <= Xxh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Diva17 <= 1'b0;
  else
    Diva17 <= Qxh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zjva17 <= 1'b0;
  else
    Zjva17 <= Jxh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vlva17 <= 1'b0;
  else
    Vlva17 <= Cxh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rnva17 <= 1'b0;
  else
    Rnva17 <= Vwh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Npva17 <= 1'b0;
  else
    Npva17 <= Owh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jrva17 <= 1'b0;
  else
    Jrva17 <= Hwh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ftva17 <= 1'b0;
  else
    Ftva17 <= Awh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bvva17 <= 1'b0;
  else
    Bvva17 <= Tvh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xwva17 <= 1'b0;
  else
    Xwva17 <= Mvh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tyva17 <= 1'b0;
  else
    Tyva17 <= Fvh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    P0wa17 <= 1'b0;
  else
    P0wa17 <= Yuh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    K2wa17 <= 1'b0;
  else
    K2wa17 <= Ruh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    F4wa17 <= 1'b0;
  else
    F4wa17 <= Kuh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    A6wa17 <= 1'b0;
  else
    A6wa17 <= Duh7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    V7wa17 <= 1'b0;
  else
    V7wa17 <= Wth7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Q9wa17 <= 1'b0;
  else
    Q9wa17 <= Pth7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lbwa17 <= 1'b0;
  else
    Lbwa17 <= Ith7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gdwa17 <= 1'b0;
  else
    Gdwa17 <= Bth7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Bfwa17 <= 1'b0;
  else
    Bfwa17 <= Ush7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wgwa17 <= 1'b0;
  else
    Wgwa17 <= X447v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Oiwa17 <= 1'b0;
  else
    Oiwa17 <= I6q7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mkwa17 <= 1'b0;
  else
    Mkwa17 <= P6q7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Kmwa17 <= 1'b0;
  else
    Kmwa17 <= Rbl8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Iowa17 <= 1'b0;
  else
    Iowa17 <= Mcl8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fqwa17 <= 1'b0;
  else
    Fqwa17 <= B6q7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Wrwa17 <= 1'b0;
  else
    Wrwa17 <= Yfp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Utwa17 <= 1'b0;
  else
    Utwa17 <= Fgp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Svwa17 <= 1'b0;
  else
    Svwa17 <= Mgp7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qxwa17 <= 1'b0;
  else
    Qxwa17 <= Tgp7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ozwa17 <= 1'b1;
  else
    Ozwa17 <= K7q7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    K1xa17 <= 1'b0;
  else
    K1xa17 <= Ewq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    M4xa17 <= 1'b0;
  else
    M4xa17 <= R7q7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    O7xa17 <= 1'b0;
  else
    O7xa17 <= Kzq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vaxa17 <= 1'b0;
  else
    Vaxa17 <= Dzq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cexa17 <= 1'b0;
  else
    Cexa17 <= Rzq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Jhxa17 <= 1'b0;
  else
    Jhxa17 <= Pyq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Skxa17 <= 1'b0;
  else
    Skxa17 <= Ksq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Knxa17 <= 1'b0;
  else
    Knxa17 <= Dsq7v6;

always @(posedge FCLK) Cqxa17 <= Psp7v6;
always @(posedge FCLK) Nsxa17 <= Isp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yuxa17 <= 1'b0;
  else
    Yuxa17 <= Huq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Qxxa17 <= 1'b0;
  else
    Qxxa17 <= Auq7v6;

always @(posedge FCLK) I0ya17 <= Zqp7v6;
always @(posedge FCLK) T2ya17 <= Mmq7v6;
always @(posedge FCLK) E5ya17 <= Siq7v6;
always @(posedge FCLK) P7ya17 <= Ebq7v6;
always @(posedge FCLK) Aaya17 <= Sqp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lcya17 <= 1'b0;
  else
    Lcya17 <= Ttq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Dfya17 <= 1'b0;
  else
    Dfya17 <= Mtq7v6;

always @(posedge FCLK) Vhya17 <= Urp7v6;
always @(posedge FCLK) Gkya17 <= Nrp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rmya17 <= 1'b0;
  else
    Rmya17 <= Byq7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vpya17 <= 1'b0;
  else
    Vpya17 <= Zvr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Trya17 <= 1'b0;
  else
    Trya17 <= Atr7v6;

always @(posedge HCLK) Rtya17 <= Z1t7v6;
always @(posedge HCLK) Ovya17 <= G2t7v6;
always @(posedge HCLK) Lxya17 <= N2t7v6;
always @(posedge HCLK) Izya17 <= Vrt7v6;
always @(posedge HCLK) F1za17 <= Cst7v6;
always @(posedge HCLK) C3za17 <= Jst7v6;
always @(posedge HCLK) Z4za17 <= Xet7v6;
always @(posedge HCLK) W6za17 <= Eft7v6;
always @(posedge HCLK) T8za17 <= Lft7v6;
always @(posedge HCLK) Qaza17 <= T4u7v6;
always @(posedge HCLK) Ncza17 <= A5u7v6;
always @(posedge HCLK) Keza17 <= H5u7v6;
always @(posedge HCLK) Hgza17 <= L8t7v6;
always @(posedge HCLK) Eiza17 <= S8t7v6;
always @(posedge HCLK) Bkza17 <= Z8t7v6;
always @(posedge HCLK) Ylza17 <= Hyt7v6;
always @(posedge HCLK) Vnza17 <= Oyt7v6;
always @(posedge HCLK) Spza17 <= Vyt7v6;
always @(posedge HCLK) Prza17 <= Jlt7v6;
always @(posedge HCLK) Mtza17 <= Qlt7v6;
always @(posedge HCLK) Jvza17 <= Xlt7v6;
always @(posedge HCLK) Gxza17 <= Fbu7v6;
always @(posedge HCLK) Dzza17 <= Mbu7v6;
always @(posedge HCLK) A10b17 <= Tbu7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    X20b17 <= 1'b0;
  else
    X20b17 <= Z2s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    S40b17 <= 1'b0;
  else
    S40b17 <= O0s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Q60b17 <= 1'b0;
  else
    Q60b17 <= Kyr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    O80b17 <= 1'b0;
  else
    O80b17 <= Gwr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ma0b17 <= 1'b0;
  else
    Ma0b17 <= Htr7v6;

always @(posedge HCLK) Kc0b17 <= J0t7v6;
always @(posedge HCLK) He0b17 <= Q0t7v6;
always @(posedge HCLK) Eg0b17 <= X0t7v6;
always @(posedge HCLK) Bi0b17 <= Fqt7v6;
always @(posedge HCLK) Yj0b17 <= Mqt7v6;
always @(posedge HCLK) Vl0b17 <= Tqt7v6;
always @(posedge HCLK) Sn0b17 <= V6t7v6;
always @(posedge HCLK) Pp0b17 <= C7t7v6;
always @(posedge HCLK) Mr0b17 <= J7t7v6;
always @(posedge HCLK) Jt0b17 <= Rwt7v6;
always @(posedge HCLK) Gv0b17 <= Ywt7v6;
always @(posedge HCLK) Dx0b17 <= Fxt7v6;
always @(posedge HCLK) Az0b17 <= Hdt7v6;
always @(posedge HCLK) X01b17 <= Odt7v6;
always @(posedge HCLK) U21b17 <= Vdt7v6;
always @(posedge HCLK) R41b17 <= D3u7v6;
always @(posedge HCLK) O61b17 <= K3u7v6;
always @(posedge HCLK) L81b17 <= R3u7v6;
always @(posedge HCLK) Ia1b17 <= Tjt7v6;
always @(posedge HCLK) Fc1b17 <= Akt7v6;
always @(posedge HCLK) Ce1b17 <= Hkt7v6;
always @(posedge HCLK) Zf1b17 <= Ozs7v6;
always @(posedge HCLK) Wh1b17 <= Vzs7v6;
always @(posedge HCLK) Tj1b17 <= C0t7v6;
always @(posedge HCLK) Ql1b17 <= Kpt7v6;
always @(posedge HCLK) Nn1b17 <= Rpt7v6;
always @(posedge HCLK) Kp1b17 <= Ypt7v6;
always @(posedge HCLK) Hr1b17 <= A6t7v6;
always @(posedge HCLK) Et1b17 <= H6t7v6;
always @(posedge HCLK) Bv1b17 <= Wvt7v6;
always @(posedge HCLK) Yw1b17 <= Dwt7v6;
always @(posedge HCLK) Vy1b17 <= Kwt7v6;
always @(posedge HCLK) S02b17 <= Mct7v6;
always @(posedge HCLK) P22b17 <= Tct7v6;
always @(posedge HCLK) M42b17 <= Adt7v6;
always @(posedge HCLK) J62b17 <= I2u7v6;
always @(posedge HCLK) G82b17 <= P2u7v6;
always @(posedge HCLK) Da2b17 <= W2u7v6;
always @(posedge HCLK) Ac2b17 <= Yit7v6;
always @(posedge HCLK) Xd2b17 <= Fjt7v6;
always @(posedge HCLK) Uf2b17 <= Mjt7v6;
always @(posedge HCLK) Rh2b17 <= U8u7v6;
always @(posedge HCLK) Oj2b17 <= B9u7v6;
always @(posedge HCLK) Ll2b17 <= I9u7v6;
always @(posedge HCLK) In2b17 <= F5t7v6;
always @(posedge HCLK) Fp2b17 <= M5t7v6;
always @(posedge HCLK) Cr2b17 <= T5t7v6;
always @(posedge HCLK) Zs2b17 <= Bvt7v6;
always @(posedge HCLK) Wu2b17 <= Ivt7v6;
always @(posedge HCLK) Tw2b17 <= Pvt7v6;
always @(posedge HCLK) Qy2b17 <= Dit7v6;
always @(posedge HCLK) N03b17 <= Kit7v6;
always @(posedge HCLK) K23b17 <= Rit7v6;
always @(posedge HCLK) H43b17 <= Z7u7v6;
always @(posedge HCLK) E63b17 <= G8u7v6;
always @(posedge HCLK) B83b17 <= N8u7v6;
always @(posedge HCLK) Y93b17 <= E1t7v6;
always @(posedge HCLK) Vb3b17 <= L1t7v6;
always @(posedge HCLK) Sd3b17 <= S1t7v6;
always @(posedge HCLK) Pf3b17 <= Art7v6;
always @(posedge HCLK) Mh3b17 <= Hrt7v6;
always @(posedge HCLK) Jj3b17 <= Ort7v6;
always @(posedge HCLK) Gl3b17 <= Cet7v6;
always @(posedge HCLK) Dn3b17 <= Jet7v6;
always @(posedge HCLK) Ap3b17 <= Qet7v6;
always @(posedge HCLK) Xq3b17 <= Y3u7v6;
always @(posedge HCLK) Us3b17 <= F4u7v6;
always @(posedge HCLK) Ru3b17 <= M4u7v6;
always @(posedge HCLK) Ow3b17 <= Q7t7v6;
always @(posedge HCLK) Ly3b17 <= X7t7v6;
always @(posedge HCLK) I04b17 <= E8t7v6;
always @(posedge HCLK) F24b17 <= Mxt7v6;
always @(posedge HCLK) C44b17 <= Txt7v6;
always @(posedge HCLK) Z54b17 <= Ayt7v6;
always @(posedge HCLK) W74b17 <= Okt7v6;
always @(posedge HCLK) T94b17 <= Vkt7v6;
always @(posedge HCLK) Qb4b17 <= Clt7v6;
always @(posedge HCLK) Nd4b17 <= Kau7v6;
always @(posedge HCLK) Kf4b17 <= Rau7v6;
always @(posedge HCLK) Hh4b17 <= Yau7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ej4b17 <= 1'b0;
  else
    Ej4b17 <= G3s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zk4b17 <= 1'b0;
  else
    Zk4b17 <= V0s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xm4b17 <= 1'b0;
  else
    Xm4b17 <= Ryr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vo4b17 <= 1'b0;
  else
    Vo4b17 <= Nwr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Tq4b17 <= 1'b0;
  else
    Tq4b17 <= Otr7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Rs4b17 <= 1'b0;
  else
    Rs4b17 <= Tgw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pu4b17 <= 1'b0;
  else
    Pu4b17 <= Bpk8v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Nw4b17 <= 1'b0;
  else
    Nw4b17 <= S088v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uy4b17 <= 1'b0;
  else
    Uy4b17 <= Bp68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    X05b17 <= 1'b0;
  else
    X05b17 <= Mvo7v6;

always @(posedge HCLK) D45b17 <= Lg68v6;
always @(posedge HCLK) U55b17 <= E968v6;
always @(posedge HCLK) K75b17 <= C168v6;
always @(posedge HCLK) A95b17 <= At58v6;
always @(posedge HCLK) Qa5b17 <= Yk58v6;
always @(posedge HCLK) Gc5b17 <= Wc58v6;
always @(posedge HCLK) Wd5b17 <= U458v6;
always @(posedge HCLK) Mf5b17 <= Sw48v6;
always @(posedge HCLK) Ch5b17 <= Ep48v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Si5b17 <= 1'b0;
  else
    Si5b17 <= Zay7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sk5b17 <= 1'b0;
  else
    Sk5b17 <= A1y7v6;

always @(posedge FCLK) Um5b17 <= X2r7v6;
always @(posedge FCLK) Ro5b17 <= F8q7v6;
always @(posedge FCLK) Cr5b17 <= M8q7v6;
always @(posedge FCLK) Nt5b17 <= H9q7v6;
always @(posedge FCLK) Yv5b17 <= V9q7v6;
always @(posedge FCLK) Jy5b17 <= Caq7v6;
always @(posedge FCLK) U06b17 <= Qaq7v6;
always @(posedge FCLK) F36b17 <= Xaq7v6;
always @(posedge HCLK) Q56b17 <= Li48v6;
always @(posedge HCLK) T86b17 <= Si48v6;
always @(posedge HCLK) Wb6b17 <= Nsh7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qe6b17 <= 1'b0;
  else
    Qe6b17 <= Rq68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tg6b17 <= 1'b0;
  else
    Tg6b17 <= Cxo7v6;

always @(posedge HCLK) Zj6b17 <= Bi68v6;
always @(posedge HCLK) Ql6b17 <= Ua68v6;
always @(posedge HCLK) Gn6b17 <= S268v6;
always @(posedge HCLK) Wo6b17 <= Qu58v6;
always @(posedge HCLK) Mq6b17 <= Om58v6;
always @(posedge HCLK) Cs6b17 <= Me58v6;
always @(posedge HCLK) St6b17 <= K658v6;
always @(posedge HCLK) Iv6b17 <= Iy48v6;
always @(posedge HCLK) Yw6b17 <= Uq48v6;
always @(posedge FCLK) Oy6b17 <= N4r7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L07b17 <= 1'b0;
  else
    L07b17 <= Xll8v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    M37b17 <= 1'b0;
  else
    M37b17 <= Hlk8v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Q57b17 <= 1'b0;
  else
    Q57b17 <= V3w7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    R67b17 <= 1'b0;
  else
    R67b17 <= Pmv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    T77b17 <= 1'b0;
  else
    T77b17 <= Wmv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    V87b17 <= 1'b0;
  else
    V87b17 <= H3w7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    W97b17 <= 1'b0;
  else
    W97b17 <= A3w7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Xa7b17 <= 1'b0;
  else
    Xa7b17 <= T2w7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Yb7b17 <= 1'b0;
  else
    Yb7b17 <= M2w7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Zc7b17 <= 1'b0;
  else
    Zc7b17 <= Y1w7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Yg5m17 <= 1'b0;
  else
    Yg5m17 <= R1w7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Ai5m17 <= 1'b0;
  else
    Ai5m17 <= K1w7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Cj5m17 <= 1'b0;
  else
    Cj5m17 <= D1w7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Ek5m17 <= 1'b0;
  else
    Ek5m17 <= W0w7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Gl5m17 <= 1'b0;
  else
    Gl5m17 <= P0w7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Im5m17 <= 1'b0;
  else
    Im5m17 <= I0w7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Kn5m17 <= 1'b0;
  else
    Kn5m17 <= B0w7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Mo5m17 <= 1'b0;
  else
    Mo5m17 <= Uzv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Op5m17 <= 1'b0;
  else
    Op5m17 <= Gzv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Qq5m17 <= 1'b0;
  else
    Qq5m17 <= Zyv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Sr5m17 <= 1'b0;
  else
    Sr5m17 <= Syv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Us5m17 <= 1'b0;
  else
    Us5m17 <= Lyv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Wt5m17 <= 1'b0;
  else
    Wt5m17 <= Eyv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Yu5m17 <= 1'b0;
  else
    Yu5m17 <= Xxv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Aw5m17 <= 1'b0;
  else
    Aw5m17 <= Qxv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Cx5m17 <= 1'b0;
  else
    Cx5m17 <= Jxv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Ey5m17 <= 1'b0;
  else
    Ey5m17 <= Cxv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Gz5m17 <= 1'b0;
  else
    Gz5m17 <= Vwv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    I06m17 <= 1'b0;
  else
    I06m17 <= Owv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    K16m17 <= 1'b0;
  else
    K16m17 <= Hwv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    M26m17 <= 1'b0;
  else
    M26m17 <= Awv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    O36m17 <= 1'b0;
  else
    O36m17 <= Tvv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Q46m17 <= 1'b0;
  else
    Q46m17 <= Mvv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    S56m17 <= 1'b0;
  else
    S56m17 <= Fvv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    U66m17 <= 1'b0;
  else
    U66m17 <= Yuv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    W76m17 <= 1'b0;
  else
    W76m17 <= Ruv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Y86m17 <= 1'b0;
  else
    Y86m17 <= Kuv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Aa6m17 <= 1'b0;
  else
    Aa6m17 <= Duv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Cb6m17 <= 1'b0;
  else
    Cb6m17 <= Wtv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Ec6m17 <= 1'b0;
  else
    Ec6m17 <= Ptv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Gd6m17 <= 1'b0;
  else
    Gd6m17 <= Itv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Ie6m17 <= 1'b0;
  else
    Ie6m17 <= Btv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Kf6m17 <= 1'b0;
  else
    Kf6m17 <= Usv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Mg6m17 <= 1'b0;
  else
    Mg6m17 <= Nsv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Oh6m17 <= 1'b0;
  else
    Oh6m17 <= Gsv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Qi6m17 <= 1'b0;
  else
    Qi6m17 <= Zrv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Sj6m17 <= 1'b0;
  else
    Sj6m17 <= Srv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Uk6m17 <= 1'b0;
  else
    Uk6m17 <= Lrv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Wl6m17 <= 1'b0;
  else
    Wl6m17 <= Erv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Ym6m17 <= 1'b0;
  else
    Ym6m17 <= Xqv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Ao6m17 <= 1'b0;
  else
    Ao6m17 <= Qqv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Cp6m17 <= 1'b0;
  else
    Cp6m17 <= Jqv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Eq6m17 <= 1'b0;
  else
    Eq6m17 <= Cqv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Gr6m17 <= 1'b0;
  else
    Gr6m17 <= Vpv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Is6m17 <= 1'b0;
  else
    Is6m17 <= Opv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Kt6m17 <= 1'b0;
  else
    Kt6m17 <= Hpv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Mu6m17 <= 1'b0;
  else
    Mu6m17 <= Apv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Ov6m17 <= 1'b0;
  else
    Ov6m17 <= Mov7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Qw6m17 <= 1'b0;
  else
    Qw6m17 <= Fov7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Sx6m17 <= 1'b0;
  else
    Sx6m17 <= Ynv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Uy6m17 <= 1'b0;
  else
    Uy6m17 <= Rnv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Wz6m17 <= 1'b0;
  else
    Wz6m17 <= Knv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Y07m17 <= 1'b0;
  else
    Y07m17 <= Dnv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    A27m17 <= 1'b0;
  else
    A27m17 <= O3w7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    B37m17 <= 1'b0;
  else
    B37m17 <= Bxr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Z47m17 <= 1'b0;
  else
    Z47m17 <= Cur7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    X67m17 <= 1'b0;
  else
    X67m17 <= Gsh7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y87m17 <= 1'b0;
  else
    Y87m17 <= W4k8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fb7m17 <= 1'b0;
  else
    Fb7m17 <= S9s7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Je7m17 <= 1'b0;
  else
    Je7m17 <= O7s7v6;

always @(posedge FCLK) Nh7m17 <= Qa48v6;
always @(posedge FCLK) Tj7m17 <= Xa48v6;
always @(posedge FCLK) Zl7m17 <= Eb48v6;
always @(posedge FCLK) Fo7m17 <= Lb48v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Lq7m17 <= 1'b0;
  else
    Lq7m17 <= Uwr7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Js7m17 <= 1'b0;
  else
    Js7m17 <= Vtr7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hu7m17 <= 1'b0;
  else
    Hu7m17 <= Nrw7v6;

always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fw7m17 <= 1'b0;
  else
    Fw7m17 <= Ozfet6;

always @(posedge FCLK) Jy7m17 <= M7r7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    G08m17 <= 1'b1;
  else
    G08m17 <= Ftq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    N28m17 <= 1'b0;
  else
    N28m17 <= Ysq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    E58m17 <= 1'b0;
  else
    E58m17 <= Rsq7v6;

always @(posedge FCLK) V78m17 <= Jaq7v6;
always @(posedge FCLK) Ka8m17 <= Grp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zc8m17 <= 1'b0;
  else
    Zc8m17 <= Rkr7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ye8m17 <= 1'b0;
  else
    Ye8m17 <= Kkr7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ph8m17 <= 1'b0;
  else
    Ph8m17 <= Dkr7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Gk8m17 <= 1'b1;
  else
    Gk8m17 <= Wjr7v6;

always @(posedge FCLK) Nm8m17 <= Xpp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Cp8m17 <= 1'b1;
  else
    Cp8m17 <= Tlr7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Br8m17 <= 1'b0;
  else
    Br8m17 <= Mlr7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    At8m17 <= 1'b0;
  else
    At8m17 <= Flr7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zu8m17 <= 1'b0;
  else
    Zu8m17 <= Ykr7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yw8m17 <= 1'b1;
  else
    Yw8m17 <= Wrq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fz8m17 <= 1'b0;
  else
    Fz8m17 <= Prq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    W19m17 <= 1'b0;
  else
    W19m17 <= Irq7v6;

always @(posedge FCLK) N49m17 <= O9q7v6;
always @(posedge FCLK) C79m17 <= Bsp7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    R99m17 <= 1'b1;
  else
    R99m17 <= Cvq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Yb9m17 <= 1'b0;
  else
    Yb9m17 <= Vuq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Pe9m17 <= 1'b0;
  else
    Pe9m17 <= Ouq7v6;

always @(posedge FCLK) Gh9m17 <= Y7q7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Vj9m17 <= 1'b0;
  else
    Vj9m17 <= Gqq7v6;

always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Mm9m17 <= 1'b0;
  else
    Mm9m17 <= Zpq7v6;

always @(posedge FCLK) Dp9m17 <= A9q7v6;
always @(posedge FCLK) Or9m17 <= T8q7v6;
always @(posedge FCLK) Du9m17 <= Dtp7v6;
always @(posedge FCLK) Ow9m17 <= Wsp7v6;
always @(posedge HCLK) Dz9m17 <= Cf68v6;
always @(posedge HCLK) T0am17 <= He68v6;
always @(posedge HCLK) I2am17 <= F668v6;
always @(posedge HCLK) X3am17 <= Dy58v6;
always @(posedge HCLK) M5am17 <= Bq58v6;
always @(posedge HCLK) B7am17 <= Zh58v6;
always @(posedge HCLK) Q8am17 <= X958v6;
always @(posedge HCLK) Faam17 <= V158v6;
always @(posedge HCLK) Ubam17 <= Hu48v6;
always @(posedge FCLK) Jdam17 <= Cjv7v6;
always @(posedge FCLK) Pfam17 <= Ygv7v6;
always @(posedge FCLK) Vham17 <= A8r7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sjam17 <= 1'b0;
  else
    Sjam17 <= H7s7v6;

always @(posedge FCLK) Wmam17 <= O1r7v6;
always @(posedge FCLK) Toam17 <= O948v6;
always @(posedge FCLK) Zqam17 <= Nxq7v6;
always @(posedge FCLK) Ntam17 <= Rgv7v6;
always @(posedge FCLK) Tvam17 <= T7r7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Qxam17 <= 1'b0;
  else
    Qxam17 <= A7s7v6;

always @(posedge FCLK) U0bm17 <= Oiv7v6;
always @(posedge FCLK) A3bm17 <= Zwq7v6;
always @(posedge FCLK) O5bm17 <= Z3r7v6;
always @(posedge FCLK) L7bm17 <= D6r7v6;
always @(posedge FCLK) I9bm17 <= H2q7v6;
always @(posedge FCLK) Tbbm17 <= O2q7v6;
always @(posedge FCLK) Eebm17 <= Hop7v6;
always @(posedge FCLK) Tgbm17 <= C3q7v6;
always @(posedge FCLK) Ejbm17 <= J3q7v6;
always @(posedge FCLK) Plbm17 <= V2q7v6;
always @(posedge FCLK) Eobm17 <= X3q7v6;
always @(posedge FCLK) Pqbm17 <= E4q7v6;
always @(posedge FCLK) Atbm17 <= Q3q7v6;
always @(posedge FCLK) Pvbm17 <= S4q7v6;
always @(posedge FCLK) Aybm17 <= Z4q7v6;
always @(posedge FCLK) L0cm17 <= L4q7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    A3cm17 <= 1'b0;
  else
    A3cm17 <= Pol8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    B6cm17 <= 1'b0;
  else
    B6cm17 <= Owo7v6;

always @(posedge HCLK) H9cm17 <= G3z7v6;
always @(posedge HCLK) Rbcm17 <= Ofy7v6;
always @(posedge FCLK) Pecm17 <= C2r7v6;
always @(posedge HCLK) Mgcm17 <= Suz7v6;
always @(posedge HCLK) Djcm17 <= I308v6;
always @(posedge HCLK) Ulcm17 <= Yb08v6;
always @(posedge HCLK) Locm17 <= Ok08v6;
always @(posedge HCLK) Crcm17 <= Et08v6;
always @(posedge HCLK) Ttcm17 <= U118v6;
always @(posedge HCLK) Kwcm17 <= Ka18v6;
always @(posedge HCLK) Bzcm17 <= Aj18v6;
always @(posedge HCLK) S1dm17 <= Qr18v6;
always @(posedge HCLK) J4dm17 <= G028v6;
always @(posedge HCLK) B7dm17 <= W828v6;
always @(posedge HCLK) T9dm17 <= Mh28v6;
always @(posedge HCLK) Lcdm17 <= Op28v6;
always @(posedge HCLK) Dfdm17 <= Ey28v6;
always @(posedge HCLK) Vhdm17 <= G638v6;
always @(posedge HCLK) Nkdm17 <= Ozk8v6;
always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Endm17 <= 1'b0;
  else
    Endm17 <= Zqw7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fodm17 <= 1'b0;
  else
    Fodm17 <= Nas7v6;

always @(posedge FCLK) Irdm17 <= Q2r7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ftdm17 <= 1'b0;
  else
    Ftdm17 <= J8s7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jwdm17 <= 1'b0;
  else
    Jwdm17 <= Pp68v6;

always @(posedge HCLK) Mydm17 <= Zg68v6;
always @(posedge HCLK) D0em17 <= S968v6;
always @(posedge HCLK) T1em17 <= Q168v6;
always @(posedge HCLK) J3em17 <= Ot58v6;
always @(posedge HCLK) Z4em17 <= Ml58v6;
always @(posedge HCLK) P6em17 <= Kd58v6;
always @(posedge HCLK) F8em17 <= I558v6;
always @(posedge HCLK) V9em17 <= Gx48v6;
always @(posedge HCLK) Lbem17 <= Sp48v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bdem17 <= 1'b0;
  else
    Bdem17 <= O1y7v6;

always @(posedge FCLK) Dfem17 <= L3r7v6;
always @(posedge FCLK) Ahem17 <= Tup7v6;
always @(posedge FCLK) Ljem17 <= Avp7v6;
always @(posedge FCLK) Wlem17 <= Jpp7v6;
always @(posedge FCLK) Loem17 <= Ovp7v6;
always @(posedge FCLK) Wqem17 <= Vvp7v6;
always @(posedge FCLK) Htem17 <= Hvp7v6;
always @(posedge FCLK) Wvem17 <= Jwp7v6;
always @(posedge FCLK) Hyem17 <= Qwp7v6;
always @(posedge FCLK) S0fm17 <= Cwp7v6;
always @(posedge FCLK) H3fm17 <= Exp7v6;
always @(posedge FCLK) S5fm17 <= Lxp7v6;
always @(posedge FCLK) D8fm17 <= Xwp7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Safm17 <= 1'b0;
  else
    Safm17 <= Dpl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tdfm17 <= 1'b0;
  else
    Tdfm17 <= Awo7v6;

always @(posedge HCLK) Zgfm17 <= V3p7v6;
always @(posedge FCLK) Dkfm17 <= D8w7v6;
always @(posedge FCLK) Rmfm17 <= Haw7v6;
always @(posedge FCLK) Fpfm17 <= Lcw7v6;
always @(posedge FCLK) Srfm17 <= Anq7v6;
always @(posedge FCLK) Dufm17 <= Hnq7v6;
always @(posedge FCLK) Owfm17 <= Qpp7v6;
always @(posedge FCLK) Dzfm17 <= Vnq7v6;
always @(posedge FCLK) O1gm17 <= Coq7v6;
always @(posedge FCLK) Z3gm17 <= Onq7v6;
always @(posedge FCLK) O6gm17 <= Qoq7v6;
always @(posedge FCLK) Z8gm17 <= Xoq7v6;
always @(posedge FCLK) Kbgm17 <= Joq7v6;
always @(posedge FCLK) Zdgm17 <= Lpq7v6;
always @(posedge FCLK) Kggm17 <= Spq7v6;
always @(posedge FCLK) Vigm17 <= Epq7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Klgm17 <= 1'b0;
  else
    Klgm17 <= P4s7v6;

always @(posedge FCLK) Oogm17 <= C9r7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kqgm17 <= 1'b0;
  else
    Kqgm17 <= F6s7v6;

always @(posedge FCLK) Otgm17 <= Y6r7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lvgm17 <= 1'b0;
  else
    Lvgm17 <= Orl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lygm17 <= 1'b0;
  else
    Lygm17 <= Xsl8v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    M1hm17 <= 1'b0;
  else
    M1hm17 <= Tov7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    O2hm17 <= 1'b0;
  else
    O2hm17 <= Nzv7v6;

always @(posedge FCLK or negedge Py9dt6)
  if(~Py9dt6)
    Q3hm17 <= 1'b0;
  else
    Q3hm17 <= F2w7v6;

always @(posedge FCLK) R4hm17 <= R6r7v6;
always @(posedge FCLK) O6hm17 <= Tfq7v6;
always @(posedge FCLK) Z8hm17 <= Agq7v6;
always @(posedge FCLK) Kbhm17 <= Mfq7v6;
always @(posedge FCLK) Zdhm17 <= Ogq7v6;
always @(posedge FCLK) Kghm17 <= Vgq7v6;
always @(posedge FCLK) Vihm17 <= Hgq7v6;
always @(posedge FCLK) Klhm17 <= Jhq7v6;
always @(posedge FCLK) Vnhm17 <= Qhq7v6;
always @(posedge FCLK) Gqhm17 <= Chq7v6;
always @(posedge FCLK) Vshm17 <= Eiq7v6;
always @(posedge FCLK) Gvhm17 <= Liq7v6;
always @(posedge FCLK) Rxhm17 <= Xhq7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    G0im17 <= 1'b0;
  else
    G0im17 <= Uxi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    J3im17 <= 1'b0;
  else
    J3im17 <= Y5s7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    N6im17 <= 1'b0;
  else
    N6im17 <= Dmp7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    L8im17 <= 1'b0;
  else
    L8im17 <= Zrh7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Maim17 <= 1'b0;
  else
    Maim17 <= Kq68v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pcim17 <= 1'b0;
  else
    Pcim17 <= Vwo7v6;

always @(posedge HCLK) Vfim17 <= Uh68v6;
always @(posedge HCLK) Mhim17 <= Na68v6;
always @(posedge HCLK) Cjim17 <= L268v6;
always @(posedge HCLK) Skim17 <= Ju58v6;
always @(posedge HCLK) Imim17 <= Hm58v6;
always @(posedge HCLK) Ynim17 <= Fe58v6;
always @(posedge HCLK) Opim17 <= D658v6;
always @(posedge HCLK) Erim17 <= By48v6;
always @(posedge HCLK) Usim17 <= Nq48v6;
always @(posedge FCLK) Kuim17 <= G4r7v6;
always @(posedge FCLK) Hwim17 <= Njq7v6;
always @(posedge FCLK) Syim17 <= Ujq7v6;
always @(posedge FCLK) D1jm17 <= Gjq7v6;
always @(posedge FCLK) S3jm17 <= Ikq7v6;
always @(posedge FCLK) D6jm17 <= Pkq7v6;
always @(posedge FCLK) O8jm17 <= Bkq7v6;
always @(posedge FCLK) Dbjm17 <= Dlq7v6;
always @(posedge FCLK) Odjm17 <= Klq7v6;
always @(posedge FCLK) Zfjm17 <= Wkq7v6;
always @(posedge FCLK) Oijm17 <= Ylq7v6;
always @(posedge FCLK) Zkjm17 <= Fmq7v6;
always @(posedge FCLK) Knjm17 <= Rlq7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Zpjm17 <= 1'b0;
  else
    Zpjm17 <= Blp7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Xrjm17 <= 1'b0;
  else
    Xrjm17 <= Srh7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ytjm17 <= 1'b0;
  else
    Ytjm17 <= Akl8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ywjm17 <= 1'b0;
  else
    Ywjm17 <= D1p7v6;

always @(posedge HCLK) D0km17 <= E5p7v6;
always @(posedge HCLK) H3km17 <= S2k8v6;
always @(posedge HCLK) A5km17 <= L2k8v6;
always @(posedge HCLK) T6km17 <= Ddj8v6;
always @(posedge HCLK) M8km17 <= Pcj8v6;
always @(posedge HCLK) Fakm17 <= Sxh8v6;
always @(posedge HCLK) Wbkm17 <= Iu88v6;
always @(posedge HCLK) Pdkm17 <= Vj88v6;
always @(posedge HCLK) Ifkm17 <= Hj88v6;
always @(posedge HCLK) Fhkm17 <= Ikx7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yikm17 <= 1'b0;
  else
    Yikm17 <= V1y7v6;

always @(posedge FCLK) Alkm17 <= S3r7v6;
always @(posedge FCLK) Xmkm17 <= W5r7v6;
always @(posedge FCLK) Uokm17 <= Nyp7v6;
always @(posedge FCLK) Frkm17 <= Uyp7v6;
always @(posedge FCLK) Qtkm17 <= Vop7v6;
always @(posedge FCLK) Fwkm17 <= Izp7v6;
always @(posedge FCLK) Qykm17 <= Pzp7v6;
always @(posedge FCLK) B1lm17 <= Bzp7v6;
always @(posedge FCLK) Q3lm17 <= D0q7v6;
always @(posedge FCLK) B6lm17 <= K0q7v6;
always @(posedge FCLK) M8lm17 <= Wzp7v6;
always @(posedge FCLK) Bblm17 <= Y0q7v6;
always @(posedge FCLK) Mdlm17 <= F1q7v6;
always @(posedge FCLK) Xflm17 <= R0q7v6;
always @(posedge FCLK) Milm17 <= T1q7v6;
always @(posedge FCLK) Xklm17 <= A2q7v6;
always @(posedge FCLK) Inlm17 <= M1q7v6;
always @(posedge FCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xplm17 <= 1'b0;
  else
    Xplm17 <= Oop7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Xrlm17 <= 1'b0;
  else
    Xrlm17 <= Xip7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Vtlm17 <= 1'b0;
  else
    Vtlm17 <= Lrh7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Wvlm17 <= 1'b0;
  else
    Wvlm17 <= A3p7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xylm17 <= 1'b0;
  else
    Xylm17 <= M2p7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Y1mm17 <= 1'b0;
  else
    Y1mm17 <= T2p7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z4mm17 <= 1'b0;
  else
    Z4mm17 <= W0p7v6;

always @(posedge HCLK) E8mm17 <= Nqi8v6;
always @(posedge HCLK) Abmm17 <= Spi8v6;
always @(posedge HCLK) Wdmm17 <= Chx7v6;
always @(posedge HCLK) Sgmm17 <= Sro7v6;
always @(posedge HCLK) Mjmm17 <= Uso7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Cmmm17 <= 1'b0;
  else
    Cmmm17 <= Ox88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xomm17 <= 1'b0;
  else
    Xomm17 <= Byi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Asmm17 <= 1'b0;
  else
    Asmm17 <= Vx88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Vumm17 <= 1'b0;
  else
    Vumm17 <= Iyi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Yxmm17 <= 1'b0;
  else
    Yxmm17 <= Cy88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    T0nm17 <= 1'b0;
  else
    T0nm17 <= Pyi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    W3nm17 <= 1'b0;
  else
    W3nm17 <= Jy88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    R6nm17 <= 1'b0;
  else
    R6nm17 <= Qy88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M9nm17 <= 1'b0;
  else
    M9nm17 <= Dzi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pcnm17 <= 1'b0;
  else
    Pcnm17 <= Xy88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Kfnm17 <= 1'b0;
  else
    Kfnm17 <= Kzi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ninm17 <= 1'b0;
  else
    Ninm17 <= Ez88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ilnm17 <= 1'b0;
  else
    Ilnm17 <= Rzi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lonm17 <= 1'b0;
  else
    Lonm17 <= Lz88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Grnm17 <= 1'b0;
  else
    Grnm17 <= Yzi8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Junm17 <= 1'b0;
  else
    Junm17 <= Sz88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Exnm17 <= 1'b0;
  else
    Exnm17 <= F0j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    I0om17 <= 1'b0;
  else
    I0om17 <= Zz88v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D3om17 <= 1'b0;
  else
    D3om17 <= M0j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    H6om17 <= 1'b0;
  else
    H6om17 <= T0j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    L9om17 <= 1'b0;
  else
    L9om17 <= A1j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Pcom17 <= 1'b0;
  else
    Pcom17 <= H1j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tfom17 <= 1'b0;
  else
    Tfom17 <= O1j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xiom17 <= 1'b0;
  else
    Xiom17 <= V1j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Bmom17 <= 1'b0;
  else
    Bmom17 <= C2j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fpom17 <= 1'b0;
  else
    Fpom17 <= J2j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jsom17 <= 1'b0;
  else
    Jsom17 <= Q2j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Nvom17 <= 1'b0;
  else
    Nvom17 <= X2j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ryom17 <= 1'b0;
  else
    Ryom17 <= E3j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V1pm17 <= 1'b0;
  else
    V1pm17 <= L3j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Z4pm17 <= 1'b0;
  else
    Z4pm17 <= S3j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    D8pm17 <= 1'b0;
  else
    D8pm17 <= Z3j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Hbpm17 <= 1'b0;
  else
    Hbpm17 <= G4j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Lepm17 <= 1'b0;
  else
    Lepm17 <= N4j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Phpm17 <= 1'b0;
  else
    Phpm17 <= U4j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Tkpm17 <= 1'b0;
  else
    Tkpm17 <= B5j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Xnpm17 <= 1'b0;
  else
    Xnpm17 <= I5j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Brpm17 <= 1'b0;
  else
    Brpm17 <= P5j8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Fupm17 <= 1'b0;
  else
    Fupm17 <= Qel8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Jxpm17 <= 1'b0;
  else
    Jxpm17 <= Nxi8v6;

always @(posedge HCLK) M0qm17 <= Qbp7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    P3qm17 <= 1'b0;
  else
    P3qm17 <= An48v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    A5qm17 <= 1'b0;
  else
    A5qm17 <= Wal8v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Y6qm17 <= 1'b0;
  else
    Y6qm17 <= Erh7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Z8qm17 <= 1'b0;
  else
    Z8qm17 <= Rfp7v6;

always @(posedge TRACECLKIN) Xaqm17 <= Xqh7v6;
always @(posedge TRACECLKIN) Wcqm17 <= Qqh7v6;
always @(posedge TRACECLKIN) Veqm17 <= Jqh7v6;
always @(posedge TRACECLKIN) Ugqm17 <= Cqh7v6;
always @(posedge TRACECLKIN) Tiqm17 <= Vph7v6;
always @(posedge TRACECLKIN) Skqm17 <= Oph7v6;
always @(posedge TRACECLKIN) Rmqm17 <= Hph7v6;
always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Qoqm17 <= 1'b0;
  else
    Qoqm17 <= Wep7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Rqqm17 <= 1'b0;
  else
    Rqqm17 <= Pep7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Ssqm17 <= 1'b0;
  else
    Ssqm17 <= Bep7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Tuqm17 <= 1'b0;
  else
    Tuqm17 <= Ndp7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Uwqm17 <= 1'b0;
  else
    Uwqm17 <= Zcp7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Syqm17 <= 1'b0;
  else
    Syqm17 <= Kfp7v6;

always @(posedge FCLK) T0rm17 <= U4r7v6;
always @(posedge FCLK) Q2rm17 <= Zbq7v6;
always @(posedge FCLK) B5rm17 <= Gcq7v6;
always @(posedge FCLK) M7rm17 <= Sbq7v6;
always @(posedge FCLK) Barm17 <= Ucq7v6;
always @(posedge FCLK) Mcrm17 <= Bdq7v6;
always @(posedge FCLK) Xerm17 <= Ncq7v6;
always @(posedge FCLK) Mhrm17 <= Pdq7v6;
always @(posedge FCLK) Xjrm17 <= Wdq7v6;
always @(posedge FCLK) Imrm17 <= Idq7v6;
always @(posedge FCLK) Xorm17 <= Keq7v6;
always @(posedge FCLK) Irrm17 <= Req7v6;
always @(posedge FCLK) Ttrm17 <= Deq7v6;
always @(posedge FCLK) Iwrm17 <= Yeq7v6;
always @(posedge FCLK) Tyrm17 <= Ffq7v6;
always @(posedge FCLK) E1sm17 <= Rmp7v6;
always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    T3sm17 <= 1'b0;
  else
    T3sm17 <= Yvu7v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    V5sm17 <= 1'b0;
  else
    V5sm17 <= Ive8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    N7sm17 <= 1'b0;
  else
    N7sm17 <= Lme8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    A9sm17 <= 1'b0;
  else
    A9sm17 <= Eme8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Oasm17 <= 1'b0;
  else
    Oasm17 <= Wyi8v6;

always @(posedge HCLK) Rdsm17 <= T9p7v6;
always @(posedge FCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ugsm17 <= 1'b0;
  else
    Ugsm17 <= Idi8v6;

always @(posedge HCLK) Ajsm17 <= Oj88v6;
always @(posedge HCLK) Tksm17 <= Gso7v6;
always @(posedge HCLK) Jnsm17 <= Aph7v6;
always @(posedge HCLK) Dqsm17 <= Aj88v6;
always @(posedge HCLK) Assm17 <= Ero7v6;
always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Uusm17 <= 1'b0;
  else
    Uusm17 <= Mg38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Sxsm17 <= 1'b0;
  else
    Sxsm17 <= Hh38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Q0tm17 <= 1'b0;
  else
    Q0tm17 <= Q0l8v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    O3tm17 <= 1'b0;
  else
    O3tm17 <= Oh38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    M6tm17 <= 1'b0;
  else
    M6tm17 <= Ah38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    K9tm17 <= 1'b0;
  else
    K9tm17 <= Tg38v6;

always @(posedge HCLK or negedge H8bdt6)
  if(~H8bdt6)
    Ictm17 <= 1'b0;
  else
    Ictm17 <= Tly7v6;

always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Fftm17 <= 1'b0;
  else
    Fftm17 <= Zjp7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Dhtm17 <= 1'b0;
  else
    Dhtm17 <= Toh7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Ejtm17 <= 1'b0;
  else
    Ejtm17 <= Iep7v6;

always @(posedge HCLK) Fltm17 <= Cr88v6;
always @(posedge HCLK) Vntm17 <= Vq88v6;
always @(posedge HCLK) Lqtm17 <= Oq88v6;
always @(posedge HCLK) Bttm17 <= Hq88v6;
always @(posedge HCLK) Svtm17 <= Aq88v6;
always @(posedge HCLK) Jytm17 <= Tp88v6;
always @(posedge HCLK) A1um17 <= Mp88v6;
always @(posedge HCLK) R3um17 <= Fp88v6;
always @(posedge HCLK) I6um17 <= Yo88v6;
always @(posedge HCLK) Z8um17 <= Ro88v6;
always @(posedge HCLK) Qbum17 <= Ko88v6;
always @(posedge HCLK) Heum17 <= Do88v6;
always @(posedge HCLK) Ygum17 <= Wn88v6;
always @(posedge HCLK) Pjum17 <= Pn88v6;
always @(posedge HCLK) Gmum17 <= In88v6;
always @(posedge HCLK) Xoum17 <= Bn88v6;
always @(posedge HCLK) Orum17 <= Um88v6;
always @(posedge HCLK) Fuum17 <= Nm88v6;
always @(posedge HCLK) Wwum17 <= Gm88v6;
always @(posedge HCLK) Nzum17 <= Zl88v6;
always @(posedge HCLK) E2vm17 <= Sl88v6;
always @(posedge HCLK) V4vm17 <= Ll88v6;
always @(posedge HCLK) M7vm17 <= El88v6;
always @(posedge HCLK) Davm17 <= Xk88v6;
always @(posedge HCLK) Ucvm17 <= Qk88v6;
always @(posedge FCLK) Lfvm17 <= A1r7v6;
always @(posedge HCLK or negedge Ox9dt6)
  if(~Ox9dt6)
    Ihvm17 <= 1'b0;
  else
    Ihvm17 <= Vhp7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Gjvm17 <= 1'b0;
  else
    Gjvm17 <= Moh7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Hlvm17 <= 1'b0;
  else
    Hlvm17 <= Udp7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Invm17 <= 1'b0;
  else
    Invm17 <= Lcp7v6;

always @(posedge HCLK) Gpvm17 <= H3p7v6;
always @(posedge HCLK) Ksvm17 <= Foh7v6;
always @(posedge HCLK) Duvm17 <= Zns7v6;
always @(posedge HCLK) Wvvm17 <= Sns7v6;
always @(posedge HCLK) Pxvm17 <= Lns7v6;
always @(posedge HCLK) Izvm17 <= Ynh7v6;
always @(posedge HCLK) B1wm17 <= Pto7v6;
always @(posedge HCLK) U2wm17 <= Bto7v6;
always @(posedge HCLK) N4wm17 <= Nso7v6;
always @(posedge HCLK) G6wm17 <= Zro7v6;
always @(posedge HCLK) Z7wm17 <= Lro7v6;
always @(posedge HCLK) W9wm17 <= Xqo7v6;
always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Tbwm17 <= 1'b0;
  else
    Tbwm17 <= Rnh7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Udwm17 <= 1'b0;
  else
    Udwm17 <= Dfp7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Vfwm17 <= 1'b0;
  else
    Vfwm17 <= Scp7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Thwm17 <= 1'b0;
  else
    Thwm17 <= Ecp7v6;

always @(posedge TRACECLKIN or negedge T0adt6)
  if(~T0adt6)
    Rjwm17 <= 1'b0;
  else
    Rjwm17 <= Gdp7v6;

endmodule

//------------------------------------------------------------------------------
// EOF
//------------------------------------------------------------------------------

