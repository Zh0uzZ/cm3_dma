module Decoder_7x128 (
  input wire [6:0] select,
  output wire [127:0] outputs
);

  reg [127:0] data;

  always @* begin
    case (select)
      7'b0000000: data = 128'h00000000000000000000000000000001;
      7'b0000001: data = 128'h00000000000000000000000000000002;
      7'b0000010: data = 128'h00000000000000000000000000000004;
      7'b0000011: data = 128'h00000000000000000000000000000008;
      7'b0000100: data = 128'h00000000000000000000000000000010;
      7'b0000101: data = 128'h00000000000000000000000000000020;
      7'b0000110: data = 128'h00000000000000000000000000000040;
      7'b0000111: data = 128'h00000000000000000000000000000080;
      7'b0001000: data = 128'h00000000000000000000000000000100;
      7'b0001001: data = 128'h00000000000000000000000000000200;
      7'b0001010: data = 128'h00000000000000000000000000000400;
      7'b0001011: data = 128'h00000000000000000000000000000800;
      7'b0001100: data = 128'h00000000000000000000000000001000;
      7'b0001101: data = 128'h00000000000000000000000000002000;
      7'b0001110: data = 128'h00000000000000000000000000004000;
      7'b0001111: data = 128'h00000000000000000000000000008000;
      7'b0010000: data = 128'h00000000000000000000000000010000;
      7'b0010001: data = 128'h00000000000000000000000000020000;
      7'b0010010: data = 128'h00000000000000000000000000040000;
      7'b0010011: data = 128'h00000000000000000000000000080000;
      7'b0010100: data = 128'h00000000000000000000000000100000;
      7'b0010101: data = 128'h00000000000000000000000000200000;
      7'b0010110: data = 128'h00000000000000000000000000400000;
      7'b0010111: data = 128'h00000000000000000000000000800000;
      7'b0011000: data = 128'h00000000000000000000000001000000;
      7'b0011001: data = 128'h00000000000000000000000002000000;
      7'b0011010: data = 128'h00000000000000000000000004000000;
      7'b0011011: data = 128'h00000000000000000000000008000000;
      7'b0011100: data = 128'h00000000000000000000000010000000;
      7'b0011101: data = 128'h00000000000000000000000020000000;
      7'b0011110: data = 128'h00000000000000000000000040000000;
      7'b0011111: data = 128'h00000000000000000000000080000000;
      7'b0100000: data = 128'h00000000000000000000000100000000;
      7'b0100001: data = 128'h00000000000000000000000200000000;
      7'b0100010: data = 128'h00000000000000000000000400000000;
      7'b0100011: data = 128'h00000000000000000000000800000000;
      7'b0100100: data = 128'h00000000000000000000001000000000;
      7'b0100101: data = 128'h00000000000000000000002000000000;
      7'b0100110: data = 128'h00000000000000000000004000000000;
      7'b0100111: data = 128'h00000000000000000000008000000000;
      7'b0101000: data = 128'h00000000000000000000010000000000;
      7'b0101001: data = 128'h00000000000000000000020000000000;
      7'b0101010: data = 128'h00000000000000000000040000000000;
      7'b0101011: data = 128'h00000000000000000000080000000000;
      7'b0101100: data = 128'h00000000000000000000100000000000;
      7'b0101101: data = 128'h00000000000000000000200000000000;
      7'b0101110: data = 128'h00000000000000000000400000000000;
      7'b0101111: data = 128'h00000000000000000000800000000000;
      7'b0110000: data = 128'h00000000000000000001000000000000;
      7'b0110001: data = 128'h00000000000000000002000000000000;
      7'b0110010: data = 128'h00000000000000000004000000000000;
      7'b0110011: data = 128'h00000000000000000008000000000000;
      7'b0110100: data = 128'h00000000000000000010000000000000;
      7'b0110101: data = 128'h00000000000000000020000000000000;
      7'b0110110: data = 128'h00000000000000000040000000000000;
      7'b0110111: data = 128'h00000000000000000080000000000000;
      7'b0111000: data = 128'h00000000000000000100000000000000;
      7'b0111001: data = 128'h00000000000000000200000000000000;
      7'b0111010: data = 128'h00000000000000000400000000000000;
      7'b0111011: data = 128'h00000000000000000800000000000000;
      7'b0111100: data = 128'h00000000000000001000000000000000;
      7'b0111101: data = 128'h00000000000000002000000000000000;
      7'b0111110: data = 128'h00000000000000004000000000000000;
      7'b0111111: data = 128'h00000000000000008000000000000000;
      7'b1000000: data = 128'h00000000000000010000000000000000;
      7'b1000001: data = 128'h00000000000000020000000000000000;
      7'b1000010: data = 128'h00000000000000040000000000000000;
      7'b1000011: data = 128'h00000000000000080000000000000000;
      7'b1000100: data = 128'h00000000000000100000000000000000;
      7'b1000101: data = 128'h00000000000000200000000000000000;
      7'b1000110: data = 128'h00000000000000400000000000000000;
      7'b1000111: data = 128'h00000000000000800000000000000000;
      7'b1001000: data = 128'h00000000000001000000000000000000;
      7'b1001001: data = 128'h00000000000002000000000000000000;
      7'b1001010: data = 128'h00000000000004000000000000000000;
      7'b1001011: data = 128'h00000000000008000000000000000000;
      7'b1001100: data = 128'h00000000000010000000000000000000;
      7'b1001101: data = 128'h00000000000020000000000000000000;
      7'b1001110: data = 128'h00000000000040000000000000000000;
      7'b1001111: data = 128'h00000000000080000000000000000000;
      7'b1010000: data = 128'h00000000000100000000000000000000;
      7'b1010001: data = 128'h00000000000200000000000000000000;
      7'b1010010: data = 128'h00000000000400000000000000000000;
      7'b1010011: data = 128'h00000000000800000000000000000000;
      7'b1010100: data = 128'h00000000001000000000000000000000;
      7'b1010101: data = 128'h00000000002000000000000000000000;
      7'b1010110: data = 128'h00000000004000000000000000000000;
      7'b1010111: data = 128'h00000000008000000000000000000000;
      7'b1011000: data = 128'h00000000010000000000000000000000;
      7'b1011001: data = 128'h00000000020000000000000000000000;
      7'b1011010: data = 128'h00000000040000000000000000000000;
      7'b1011011: data = 128'h00000000080000000000000000000000;
      7'b1011100: data = 128'h00000000100000000000000000000000;
      7'b1011101: data = 128'h00000000200000000000000000000000;
      7'b1011110: data = 128'h00000000400000000000000000000000;
      7'b1011111: data = 128'h00000000800000000000000000000000;
      7'b1100000: data = 128'h00000001000000000000000000000000;
      7'b1100001: data = 128'h00000002000000000000000000000000;
      7'b1100010: data = 128'h00000004000000000000000000000000;
      7'b1100011: data = 128'h00000008000000000000000000000000;
      7'b1100100: data = 128'h00000010000000000000000000000000;
      7'b1100101: data = 128'h00000020000000000000000000000000;
      7'b1100110: data = 128'h00000040000000000000000000000000;
      7'b1100111: data = 128'h00000080000000000000000000000000;
      7'b1101000: data = 128'h00000100000000000000000000000000;
      7'b1101001: data = 128'h00000200000000000000000000000000;
      7'b1101010: data = 128'h00000400000000000000000000000000;
      7'b1101011: data = 128'h00000800000000000000000000000000;
      7'b1101100: data = 128'h00001000000000000000000000000000;
      7'b1101101: data = 128'h00002000000000000000000000000000;
      7'b1101110: data = 128'h00004000000000000000000000000000;
      7'b1101111: data = 128'h00008000000000000000000000000000;
      7'b1110000: data = 128'h00010000000000000000000000000000;
      7'b1110001: data = 128'h00020000000000000000000000000000;
      7'b1110010: data = 128'h00040000000000000000000000000000;
      7'b1110011: data = 128'h00080000000000000000000000000000;
      7'b1110100: data = 128'h00100000000000000000000000000000;
      7'b1110101: data = 128'h00200000000000000000000000000000;
      7'b1110110: data = 128'h00400000000000000000000000000000;
      7'b1110111: data = 128'h00800000000000000000000000000000;
      7'b1111000: data = 128'h01000000000000000000000000000000;
      7'b1111001: data = 128'h02000000000000000000000000000000;
      7'b1111010: data = 128'h04000000000000000000000000000000;
      7'b1111011: data = 128'h08000000000000000000000000000000;
      7'b1111100: data = 128'h10000000000000000000000000000000;
      7'b1111101: data = 128'h20000000000000000000000000000000;
      7'b1111110: data = 128'h40000000000000000000000000000000;
      7'b1111111: data = 128'h80000000000000000000000000000000;
      default: data = 128'h00000000000000000000000000000000;
    endcase
  end

  assign outputs = data;

endmodule
